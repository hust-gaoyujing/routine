`include "ux607_defines.v"


















module ux607_gpio_top(
  input   clk,
  input   rst_n,

  input                      i_icb_cmd_valid,
  output                     i_icb_cmd_ready,
  input  [`UX607_PA_SIZE-1:0]            i_icb_cmd_addr, 
  input                      i_icb_cmd_read, 
  input  [32-1:0]            i_icb_cmd_wdata,
  
  output                     i_icb_rsp_valid,
  input                      i_icb_rsp_ready,
  output [32-1:0]            i_icb_rsp_rdata,

  output  gpio_irq_0,
  output  gpio_irq_1,
  output  gpio_irq_2,
  output  gpio_irq_3,
  output  gpio_irq_4,
  output  gpio_irq_5,
  output  gpio_irq_6,
  output  gpio_irq_7,
  output  gpio_irq_8,
  output  gpio_irq_9,
  output  gpio_irq_10,
  output  gpio_irq_11,
  output  gpio_irq_12,
  output  gpio_irq_13,
  output  gpio_irq_14,
  output  gpio_irq_15,
  output  gpio_irq_16,
  output  gpio_irq_17,
  output  gpio_irq_18,
  output  gpio_irq_19,
  output  gpio_irq_20,
  output  gpio_irq_21,
  output  gpio_irq_22,
  output  gpio_irq_23,
  output  gpio_irq_24,
  output  gpio_irq_25,
  output  gpio_irq_26,
  output  gpio_irq_27,
  output  gpio_irq_28,
  output  gpio_irq_29,
  output  gpio_irq_30,
  output  gpio_irq_31,

  input   io_port_pins_0_i_ival,
  output  io_port_pins_0_o_oval,
  output  io_port_pins_0_o_oe,
  output  io_port_pins_0_o_ie,
  output  io_port_pins_0_o_pue,
  output  io_port_pins_0_o_ds,
  input   io_port_pins_1_i_ival,
  output  io_port_pins_1_o_oval,
  output  io_port_pins_1_o_oe,
  output  io_port_pins_1_o_ie,
  output  io_port_pins_1_o_pue,
  output  io_port_pins_1_o_ds,
  input   io_port_pins_2_i_ival,
  output  io_port_pins_2_o_oval,
  output  io_port_pins_2_o_oe,
  output  io_port_pins_2_o_ie,
  output  io_port_pins_2_o_pue,
  output  io_port_pins_2_o_ds,
  input   io_port_pins_3_i_ival,
  output  io_port_pins_3_o_oval,
  output  io_port_pins_3_o_oe,
  output  io_port_pins_3_o_ie,
  output  io_port_pins_3_o_pue,
  output  io_port_pins_3_o_ds,
  input   io_port_pins_4_i_ival,
  output  io_port_pins_4_o_oval,
  output  io_port_pins_4_o_oe,
  output  io_port_pins_4_o_ie,
  output  io_port_pins_4_o_pue,
  output  io_port_pins_4_o_ds,
  input   io_port_pins_5_i_ival,
  output  io_port_pins_5_o_oval,
  output  io_port_pins_5_o_oe,
  output  io_port_pins_5_o_ie,
  output  io_port_pins_5_o_pue,
  output  io_port_pins_5_o_ds,
  input   io_port_pins_6_i_ival,
  output  io_port_pins_6_o_oval,
  output  io_port_pins_6_o_oe,
  output  io_port_pins_6_o_ie,
  output  io_port_pins_6_o_pue,
  output  io_port_pins_6_o_ds,
  input   io_port_pins_7_i_ival,
  output  io_port_pins_7_o_oval,
  output  io_port_pins_7_o_oe,
  output  io_port_pins_7_o_ie,
  output  io_port_pins_7_o_pue,
  output  io_port_pins_7_o_ds,
  input   io_port_pins_8_i_ival,
  output  io_port_pins_8_o_oval,
  output  io_port_pins_8_o_oe,
  output  io_port_pins_8_o_ie,
  output  io_port_pins_8_o_pue,
  output  io_port_pins_8_o_ds,
  input   io_port_pins_9_i_ival,
  output  io_port_pins_9_o_oval,
  output  io_port_pins_9_o_oe,
  output  io_port_pins_9_o_ie,
  output  io_port_pins_9_o_pue,
  output  io_port_pins_9_o_ds,
  input   io_port_pins_10_i_ival,
  output  io_port_pins_10_o_oval,
  output  io_port_pins_10_o_oe,
  output  io_port_pins_10_o_ie,
  output  io_port_pins_10_o_pue,
  output  io_port_pins_10_o_ds,
  input   io_port_pins_11_i_ival,
  output  io_port_pins_11_o_oval,
  output  io_port_pins_11_o_oe,
  output  io_port_pins_11_o_ie,
  output  io_port_pins_11_o_pue,
  output  io_port_pins_11_o_ds,
  input   io_port_pins_12_i_ival,
  output  io_port_pins_12_o_oval,
  output  io_port_pins_12_o_oe,
  output  io_port_pins_12_o_ie,
  output  io_port_pins_12_o_pue,
  output  io_port_pins_12_o_ds,
  input   io_port_pins_13_i_ival,
  output  io_port_pins_13_o_oval,
  output  io_port_pins_13_o_oe,
  output  io_port_pins_13_o_ie,
  output  io_port_pins_13_o_pue,
  output  io_port_pins_13_o_ds,
  input   io_port_pins_14_i_ival,
  output  io_port_pins_14_o_oval,
  output  io_port_pins_14_o_oe,
  output  io_port_pins_14_o_ie,
  output  io_port_pins_14_o_pue,
  output  io_port_pins_14_o_ds,
  input   io_port_pins_15_i_ival,
  output  io_port_pins_15_o_oval,
  output  io_port_pins_15_o_oe,
  output  io_port_pins_15_o_ie,
  output  io_port_pins_15_o_pue,
  output  io_port_pins_15_o_ds,
  input   io_port_pins_16_i_ival,
  output  io_port_pins_16_o_oval,
  output  io_port_pins_16_o_oe,
  output  io_port_pins_16_o_ie,
  output  io_port_pins_16_o_pue,
  output  io_port_pins_16_o_ds,
  input   io_port_pins_17_i_ival,
  output  io_port_pins_17_o_oval,
  output  io_port_pins_17_o_oe,
  output  io_port_pins_17_o_ie,
  output  io_port_pins_17_o_pue,
  output  io_port_pins_17_o_ds,
  input   io_port_pins_18_i_ival,
  output  io_port_pins_18_o_oval,
  output  io_port_pins_18_o_oe,
  output  io_port_pins_18_o_ie,
  output  io_port_pins_18_o_pue,
  output  io_port_pins_18_o_ds,
  input   io_port_pins_19_i_ival,
  output  io_port_pins_19_o_oval,
  output  io_port_pins_19_o_oe,
  output  io_port_pins_19_o_ie,
  output  io_port_pins_19_o_pue,
  output  io_port_pins_19_o_ds,
  input   io_port_pins_20_i_ival,
  output  io_port_pins_20_o_oval,
  output  io_port_pins_20_o_oe,
  output  io_port_pins_20_o_ie,
  output  io_port_pins_20_o_pue,
  output  io_port_pins_20_o_ds,
  input   io_port_pins_21_i_ival,
  output  io_port_pins_21_o_oval,
  output  io_port_pins_21_o_oe,
  output  io_port_pins_21_o_ie,
  output  io_port_pins_21_o_pue,
  output  io_port_pins_21_o_ds,
  input   io_port_pins_22_i_ival,
  output  io_port_pins_22_o_oval,
  output  io_port_pins_22_o_oe,
  output  io_port_pins_22_o_ie,
  output  io_port_pins_22_o_pue,
  output  io_port_pins_22_o_ds,
  input   io_port_pins_23_i_ival,
  output  io_port_pins_23_o_oval,
  output  io_port_pins_23_o_oe,
  output  io_port_pins_23_o_ie,
  output  io_port_pins_23_o_pue,
  output  io_port_pins_23_o_ds,
  input   io_port_pins_24_i_ival,
  output  io_port_pins_24_o_oval,
  output  io_port_pins_24_o_oe,
  output  io_port_pins_24_o_ie,
  output  io_port_pins_24_o_pue,
  output  io_port_pins_24_o_ds,
  input   io_port_pins_25_i_ival,
  output  io_port_pins_25_o_oval,
  output  io_port_pins_25_o_oe,
  output  io_port_pins_25_o_ie,
  output  io_port_pins_25_o_pue,
  output  io_port_pins_25_o_ds,
  input   io_port_pins_26_i_ival,
  output  io_port_pins_26_o_oval,
  output  io_port_pins_26_o_oe,
  output  io_port_pins_26_o_ie,
  output  io_port_pins_26_o_pue,
  output  io_port_pins_26_o_ds,
  input   io_port_pins_27_i_ival,
  output  io_port_pins_27_o_oval,
  output  io_port_pins_27_o_oe,
  output  io_port_pins_27_o_ie,
  output  io_port_pins_27_o_pue,
  output  io_port_pins_27_o_ds,
  input   io_port_pins_28_i_ival,
  output  io_port_pins_28_o_oval,
  output  io_port_pins_28_o_oe,
  output  io_port_pins_28_o_ie,
  output  io_port_pins_28_o_pue,
  output  io_port_pins_28_o_ds,
  input   io_port_pins_29_i_ival,
  output  io_port_pins_29_o_oval,
  output  io_port_pins_29_o_oe,
  output  io_port_pins_29_o_ie,
  output  io_port_pins_29_o_pue,
  output  io_port_pins_29_o_ds,
  input   io_port_pins_30_i_ival,
  output  io_port_pins_30_o_oval,
  output  io_port_pins_30_o_oe,
  output  io_port_pins_30_o_ie,
  output  io_port_pins_30_o_pue,
  output  io_port_pins_30_o_ds,
  input   io_port_pins_31_i_ival,
  output  io_port_pins_31_o_oval,
  output  io_port_pins_31_o_oe,
  output  io_port_pins_31_o_ie,
  output  io_port_pins_31_o_pue,
  output  io_port_pins_31_o_ds,

  output  io_port_iof_0_0_i_ival,
  input   io_port_iof_0_0_o_oval,
  input   io_port_iof_0_0_o_oe,
  input   io_port_iof_0_0_o_ie,
  input   io_port_iof_0_0_o_valid,
  output  io_port_iof_0_1_i_ival,
  input   io_port_iof_0_1_o_oval,
  input   io_port_iof_0_1_o_oe,
  input   io_port_iof_0_1_o_ie,
  input   io_port_iof_0_1_o_valid,
  output  io_port_iof_0_2_i_ival,
  input   io_port_iof_0_2_o_oval,
  input   io_port_iof_0_2_o_oe,
  input   io_port_iof_0_2_o_ie,
  input   io_port_iof_0_2_o_valid,
  output  io_port_iof_0_3_i_ival,
  input   io_port_iof_0_3_o_oval,
  input   io_port_iof_0_3_o_oe,
  input   io_port_iof_0_3_o_ie,
  input   io_port_iof_0_3_o_valid,
  output  io_port_iof_0_4_i_ival,
  input   io_port_iof_0_4_o_oval,
  input   io_port_iof_0_4_o_oe,
  input   io_port_iof_0_4_o_ie,
  input   io_port_iof_0_4_o_valid,
  output  io_port_iof_0_5_i_ival,
  input   io_port_iof_0_5_o_oval,
  input   io_port_iof_0_5_o_oe,
  input   io_port_iof_0_5_o_ie,
  input   io_port_iof_0_5_o_valid,
  output  io_port_iof_0_6_i_ival,
  input   io_port_iof_0_6_o_oval,
  input   io_port_iof_0_6_o_oe,
  input   io_port_iof_0_6_o_ie,
  input   io_port_iof_0_6_o_valid,
  output  io_port_iof_0_7_i_ival,
  input   io_port_iof_0_7_o_oval,
  input   io_port_iof_0_7_o_oe,
  input   io_port_iof_0_7_o_ie,
  input   io_port_iof_0_7_o_valid,
  output  io_port_iof_0_8_i_ival,
  input   io_port_iof_0_8_o_oval,
  input   io_port_iof_0_8_o_oe,
  input   io_port_iof_0_8_o_ie,
  input   io_port_iof_0_8_o_valid,
  output  io_port_iof_0_9_i_ival,
  input   io_port_iof_0_9_o_oval,
  input   io_port_iof_0_9_o_oe,
  input   io_port_iof_0_9_o_ie,
  input   io_port_iof_0_9_o_valid,
  output  io_port_iof_0_10_i_ival,
  input   io_port_iof_0_10_o_oval,
  input   io_port_iof_0_10_o_oe,
  input   io_port_iof_0_10_o_ie,
  input   io_port_iof_0_10_o_valid,
  output  io_port_iof_0_11_i_ival,
  input   io_port_iof_0_11_o_oval,
  input   io_port_iof_0_11_o_oe,
  input   io_port_iof_0_11_o_ie,
  input   io_port_iof_0_11_o_valid,
  output  io_port_iof_0_12_i_ival,
  input   io_port_iof_0_12_o_oval,
  input   io_port_iof_0_12_o_oe,
  input   io_port_iof_0_12_o_ie,
  input   io_port_iof_0_12_o_valid,
  output  io_port_iof_0_13_i_ival,
  input   io_port_iof_0_13_o_oval,
  input   io_port_iof_0_13_o_oe,
  input   io_port_iof_0_13_o_ie,
  input   io_port_iof_0_13_o_valid,
  output  io_port_iof_0_14_i_ival,
  input   io_port_iof_0_14_o_oval,
  input   io_port_iof_0_14_o_oe,
  input   io_port_iof_0_14_o_ie,
  input   io_port_iof_0_14_o_valid,
  output  io_port_iof_0_15_i_ival,
  input   io_port_iof_0_15_o_oval,
  input   io_port_iof_0_15_o_oe,
  input   io_port_iof_0_15_o_ie,
  input   io_port_iof_0_15_o_valid,
  output  io_port_iof_0_16_i_ival,
  input   io_port_iof_0_16_o_oval,
  input   io_port_iof_0_16_o_oe,
  input   io_port_iof_0_16_o_ie,
  input   io_port_iof_0_16_o_valid,
  output  io_port_iof_0_17_i_ival,
  input   io_port_iof_0_17_o_oval,
  input   io_port_iof_0_17_o_oe,
  input   io_port_iof_0_17_o_ie,
  input   io_port_iof_0_17_o_valid,
  output  io_port_iof_0_18_i_ival,
  input   io_port_iof_0_18_o_oval,
  input   io_port_iof_0_18_o_oe,
  input   io_port_iof_0_18_o_ie,
  input   io_port_iof_0_18_o_valid,
  output  io_port_iof_0_19_i_ival,
  input   io_port_iof_0_19_o_oval,
  input   io_port_iof_0_19_o_oe,
  input   io_port_iof_0_19_o_ie,
  input   io_port_iof_0_19_o_valid,
  output  io_port_iof_0_20_i_ival,
  input   io_port_iof_0_20_o_oval,
  input   io_port_iof_0_20_o_oe,
  input   io_port_iof_0_20_o_ie,
  input   io_port_iof_0_20_o_valid,
  output  io_port_iof_0_21_i_ival,
  input   io_port_iof_0_21_o_oval,
  input   io_port_iof_0_21_o_oe,
  input   io_port_iof_0_21_o_ie,
  input   io_port_iof_0_21_o_valid,
  output  io_port_iof_0_22_i_ival,
  input   io_port_iof_0_22_o_oval,
  input   io_port_iof_0_22_o_oe,
  input   io_port_iof_0_22_o_ie,
  input   io_port_iof_0_22_o_valid,
  output  io_port_iof_0_23_i_ival,
  input   io_port_iof_0_23_o_oval,
  input   io_port_iof_0_23_o_oe,
  input   io_port_iof_0_23_o_ie,
  input   io_port_iof_0_23_o_valid,
  output  io_port_iof_0_24_i_ival,
  input   io_port_iof_0_24_o_oval,
  input   io_port_iof_0_24_o_oe,
  input   io_port_iof_0_24_o_ie,
  input   io_port_iof_0_24_o_valid,
  output  io_port_iof_0_25_i_ival,
  input   io_port_iof_0_25_o_oval,
  input   io_port_iof_0_25_o_oe,
  input   io_port_iof_0_25_o_ie,
  input   io_port_iof_0_25_o_valid,
  output  io_port_iof_0_26_i_ival,
  input   io_port_iof_0_26_o_oval,
  input   io_port_iof_0_26_o_oe,
  input   io_port_iof_0_26_o_ie,
  input   io_port_iof_0_26_o_valid,
  output  io_port_iof_0_27_i_ival,
  input   io_port_iof_0_27_o_oval,
  input   io_port_iof_0_27_o_oe,
  input   io_port_iof_0_27_o_ie,
  input   io_port_iof_0_27_o_valid,
  output  io_port_iof_0_28_i_ival,
  input   io_port_iof_0_28_o_oval,
  input   io_port_iof_0_28_o_oe,
  input   io_port_iof_0_28_o_ie,
  input   io_port_iof_0_28_o_valid,
  output  io_port_iof_0_29_i_ival,
  input   io_port_iof_0_29_o_oval,
  input   io_port_iof_0_29_o_oe,
  input   io_port_iof_0_29_o_ie,
  input   io_port_iof_0_29_o_valid,
  output  io_port_iof_0_30_i_ival,
  input   io_port_iof_0_30_o_oval,
  input   io_port_iof_0_30_o_oe,
  input   io_port_iof_0_30_o_ie,
  input   io_port_iof_0_30_o_valid,
  output  io_port_iof_0_31_i_ival,
  input   io_port_iof_0_31_o_oval,
  input   io_port_iof_0_31_o_oe,
  input   io_port_iof_0_31_o_ie,
  input   io_port_iof_0_31_o_valid,

  output  io_port_iof_1_0_i_ival,
  input   io_port_iof_1_0_o_oval,
  input   io_port_iof_1_0_o_oe,
  input   io_port_iof_1_0_o_ie,
  input   io_port_iof_1_0_o_valid,
  output  io_port_iof_1_1_i_ival,
  input   io_port_iof_1_1_o_oval,
  input   io_port_iof_1_1_o_oe,
  input   io_port_iof_1_1_o_ie,
  input   io_port_iof_1_1_o_valid,
  output  io_port_iof_1_2_i_ival,
  input   io_port_iof_1_2_o_oval,
  input   io_port_iof_1_2_o_oe,
  input   io_port_iof_1_2_o_ie,
  input   io_port_iof_1_2_o_valid,
  output  io_port_iof_1_3_i_ival,
  input   io_port_iof_1_3_o_oval,
  input   io_port_iof_1_3_o_oe,
  input   io_port_iof_1_3_o_ie,
  input   io_port_iof_1_3_o_valid,
  output  io_port_iof_1_4_i_ival,
  input   io_port_iof_1_4_o_oval,
  input   io_port_iof_1_4_o_oe,
  input   io_port_iof_1_4_o_ie,
  input   io_port_iof_1_4_o_valid,
  output  io_port_iof_1_5_i_ival,
  input   io_port_iof_1_5_o_oval,
  input   io_port_iof_1_5_o_oe,
  input   io_port_iof_1_5_o_ie,
  input   io_port_iof_1_5_o_valid,
  output  io_port_iof_1_6_i_ival,
  input   io_port_iof_1_6_o_oval,
  input   io_port_iof_1_6_o_oe,
  input   io_port_iof_1_6_o_ie,
  input   io_port_iof_1_6_o_valid,
  output  io_port_iof_1_7_i_ival,
  input   io_port_iof_1_7_o_oval,
  input   io_port_iof_1_7_o_oe,
  input   io_port_iof_1_7_o_ie,
  input   io_port_iof_1_7_o_valid,
  output  io_port_iof_1_8_i_ival,
  input   io_port_iof_1_8_o_oval,
  input   io_port_iof_1_8_o_oe,
  input   io_port_iof_1_8_o_ie,
  input   io_port_iof_1_8_o_valid,
  output  io_port_iof_1_9_i_ival,
  input   io_port_iof_1_9_o_oval,
  input   io_port_iof_1_9_o_oe,
  input   io_port_iof_1_9_o_ie,
  input   io_port_iof_1_9_o_valid,
  output  io_port_iof_1_10_i_ival,
  input   io_port_iof_1_10_o_oval,
  input   io_port_iof_1_10_o_oe,
  input   io_port_iof_1_10_o_ie,
  input   io_port_iof_1_10_o_valid,
  output  io_port_iof_1_11_i_ival,
  input   io_port_iof_1_11_o_oval,
  input   io_port_iof_1_11_o_oe,
  input   io_port_iof_1_11_o_ie,
  input   io_port_iof_1_11_o_valid,
  output  io_port_iof_1_12_i_ival,
  input   io_port_iof_1_12_o_oval,
  input   io_port_iof_1_12_o_oe,
  input   io_port_iof_1_12_o_ie,
  input   io_port_iof_1_12_o_valid,
  output  io_port_iof_1_13_i_ival,
  input   io_port_iof_1_13_o_oval,
  input   io_port_iof_1_13_o_oe,
  input   io_port_iof_1_13_o_ie,
  input   io_port_iof_1_13_o_valid,
  output  io_port_iof_1_14_i_ival,
  input   io_port_iof_1_14_o_oval,
  input   io_port_iof_1_14_o_oe,
  input   io_port_iof_1_14_o_ie,
  input   io_port_iof_1_14_o_valid,
  output  io_port_iof_1_15_i_ival,
  input   io_port_iof_1_15_o_oval,
  input   io_port_iof_1_15_o_oe,
  input   io_port_iof_1_15_o_ie,
  input   io_port_iof_1_15_o_valid,
  output  io_port_iof_1_16_i_ival,
  input   io_port_iof_1_16_o_oval,
  input   io_port_iof_1_16_o_oe,
  input   io_port_iof_1_16_o_ie,
  input   io_port_iof_1_16_o_valid,
  output  io_port_iof_1_17_i_ival,
  input   io_port_iof_1_17_o_oval,
  input   io_port_iof_1_17_o_oe,
  input   io_port_iof_1_17_o_ie,
  input   io_port_iof_1_17_o_valid,
  output  io_port_iof_1_18_i_ival,
  input   io_port_iof_1_18_o_oval,
  input   io_port_iof_1_18_o_oe,
  input   io_port_iof_1_18_o_ie,
  input   io_port_iof_1_18_o_valid,
  output  io_port_iof_1_19_i_ival,
  input   io_port_iof_1_19_o_oval,
  input   io_port_iof_1_19_o_oe,
  input   io_port_iof_1_19_o_ie,
  input   io_port_iof_1_19_o_valid,
  output  io_port_iof_1_20_i_ival,
  input   io_port_iof_1_20_o_oval,
  input   io_port_iof_1_20_o_oe,
  input   io_port_iof_1_20_o_ie,
  input   io_port_iof_1_20_o_valid,
  output  io_port_iof_1_21_i_ival,
  input   io_port_iof_1_21_o_oval,
  input   io_port_iof_1_21_o_oe,
  input   io_port_iof_1_21_o_ie,
  input   io_port_iof_1_21_o_valid,
  output  io_port_iof_1_22_i_ival,
  input   io_port_iof_1_22_o_oval,
  input   io_port_iof_1_22_o_oe,
  input   io_port_iof_1_22_o_ie,
  input   io_port_iof_1_22_o_valid,
  output  io_port_iof_1_23_i_ival,
  input   io_port_iof_1_23_o_oval,
  input   io_port_iof_1_23_o_oe,
  input   io_port_iof_1_23_o_ie,
  input   io_port_iof_1_23_o_valid,
  output  io_port_iof_1_24_i_ival,
  input   io_port_iof_1_24_o_oval,
  input   io_port_iof_1_24_o_oe,
  input   io_port_iof_1_24_o_ie,
  input   io_port_iof_1_24_o_valid,
  output  io_port_iof_1_25_i_ival,
  input   io_port_iof_1_25_o_oval,
  input   io_port_iof_1_25_o_oe,
  input   io_port_iof_1_25_o_ie,
  input   io_port_iof_1_25_o_valid,
  output  io_port_iof_1_26_i_ival,
  input   io_port_iof_1_26_o_oval,
  input   io_port_iof_1_26_o_oe,
  input   io_port_iof_1_26_o_ie,
  input   io_port_iof_1_26_o_valid,
  output  io_port_iof_1_27_i_ival,
  input   io_port_iof_1_27_o_oval,
  input   io_port_iof_1_27_o_oe,
  input   io_port_iof_1_27_o_ie,
  input   io_port_iof_1_27_o_valid,
  output  io_port_iof_1_28_i_ival,
  input   io_port_iof_1_28_o_oval,
  input   io_port_iof_1_28_o_oe,
  input   io_port_iof_1_28_o_ie,
  input   io_port_iof_1_28_o_valid,
  output  io_port_iof_1_29_i_ival,
  input   io_port_iof_1_29_o_oval,
  input   io_port_iof_1_29_o_oe,
  input   io_port_iof_1_29_o_ie,
  input   io_port_iof_1_29_o_valid,
  output  io_port_iof_1_30_i_ival,
  input   io_port_iof_1_30_o_oval,
  input   io_port_iof_1_30_o_oe,
  input   io_port_iof_1_30_o_ie,
  input   io_port_iof_1_30_o_valid,
  output  io_port_iof_1_31_i_ival,
  input   io_port_iof_1_31_o_oval,
  input   io_port_iof_1_31_o_oe,
  input   io_port_iof_1_31_o_ie,
  input   io_port_iof_1_31_o_valid
);

 
 
 

 
 
 
 
 
 
 
 
 
 
 
 
 
 
 


  wire  io_in_0_a_ready;
  assign  i_icb_cmd_ready  = io_in_0_a_ready;
  wire  io_in_0_a_valid  = i_icb_cmd_valid;
  wire  [2:0] io_in_0_a_bits_opcode  = i_icb_cmd_read ? 3'h4 : 3'h0;
  wire  [2:0] io_in_0_a_bits_param  = 3'b0;
  wire  [2:0] io_in_0_a_bits_size = 3'd2;
  wire  [4:0] io_in_0_a_bits_source  = 5'b0;
  wire  [28:0] io_in_0_a_bits_address  = {5'b0,i_icb_cmd_addr[23:0]};
  wire  [3:0] io_in_0_a_bits_mask  = 4'b1111;
  wire  [31:0] io_in_0_a_bits_data  = i_icb_cmd_wdata;

  
  wire  io_in_0_d_ready = i_icb_rsp_ready;

  wire  [2:0] io_in_0_d_bits_opcode;
  wire  [1:0] io_in_0_d_bits_param;
  wire  [2:0] io_in_0_d_bits_size;
  wire  [4:0] io_in_0_d_bits_source;
  wire  io_in_0_d_bits_sink;
  wire  [1:0] io_in_0_d_bits_addr_lo;
  wire  [31:0] io_in_0_d_bits_data;
  wire  io_in_0_d_bits_error;
  wire  io_in_0_d_valid;

  assign  i_icb_rsp_valid = io_in_0_d_valid;
  assign  i_icb_rsp_rdata = io_in_0_d_bits_data;

  
  wire  io_in_0_b_ready = 1'b0;
  wire  io_in_0_b_valid;
  wire  [2:0] io_in_0_b_bits_opcode;
  wire  [1:0] io_in_0_b_bits_param;
  wire  [2:0] io_in_0_b_bits_size;
  wire  [4:0] io_in_0_b_bits_source;
  wire  [28:0] io_in_0_b_bits_address;
  wire  [3:0] io_in_0_b_bits_mask;
  wire  [31:0] io_in_0_b_bits_data;

  
  wire  io_in_0_c_ready;
  wire  io_in_0_c_valid = 1'b0;
  wire  [2:0] io_in_0_c_bits_opcode = 3'b0;
  wire  [2:0] io_in_0_c_bits_param = 3'b0;
  wire  [2:0] io_in_0_c_bits_size = 3'd2;
  wire  [4:0] io_in_0_c_bits_source = 5'b0;
  wire  [28:0] io_in_0_c_bits_address = 29'b0;
  wire  [31:0] io_in_0_c_bits_data = 32'b0;
  wire  io_in_0_c_bits_error = 1'b0;

  
  wire  io_in_0_e_ready;
  wire  io_in_0_e_valid = 1'b0;
  wire  io_in_0_e_bits_sink = 1'b0;

ux607_gpio u_ux607_gpio(
  .clock                            (clk                              ),
  .reset                            (~rst_n                           ),

  .io_in_0_a_ready                  (io_in_0_a_ready                  ),
  .io_in_0_a_valid                  (io_in_0_a_valid                  ),
  .io_in_0_a_bits_opcode            (io_in_0_a_bits_opcode            ),
  .io_in_0_a_bits_param             (io_in_0_a_bits_param             ),
  .io_in_0_a_bits_size              (io_in_0_a_bits_size              ),
  .io_in_0_a_bits_source            (io_in_0_a_bits_source            ),
  .io_in_0_a_bits_address           (io_in_0_a_bits_address           ),
  .io_in_0_a_bits_mask              (io_in_0_a_bits_mask              ),
  .io_in_0_a_bits_data              (io_in_0_a_bits_data              ),
  .io_in_0_b_ready                  (io_in_0_b_ready                  ),
  .io_in_0_b_valid                  (io_in_0_b_valid                  ),
  .io_in_0_b_bits_opcode            (io_in_0_b_bits_opcode            ),
  .io_in_0_b_bits_param             (io_in_0_b_bits_param             ),
  .io_in_0_b_bits_size              (io_in_0_b_bits_size              ),
  .io_in_0_b_bits_source            (io_in_0_b_bits_source            ),
  .io_in_0_b_bits_address           (io_in_0_b_bits_address           ),
  .io_in_0_b_bits_mask              (io_in_0_b_bits_mask              ),
  .io_in_0_b_bits_data              (io_in_0_b_bits_data              ),
  .io_in_0_c_ready                  (io_in_0_c_ready                  ),
  .io_in_0_c_valid                  (io_in_0_c_valid                  ),
  .io_in_0_c_bits_opcode            (io_in_0_c_bits_opcode            ),
  .io_in_0_c_bits_param             (io_in_0_c_bits_param             ),
  .io_in_0_c_bits_size              (io_in_0_c_bits_size              ),
  .io_in_0_c_bits_source            (io_in_0_c_bits_source            ),
  .io_in_0_c_bits_address           (io_in_0_c_bits_address           ),
  .io_in_0_c_bits_data              (io_in_0_c_bits_data              ),
  .io_in_0_c_bits_error             (io_in_0_c_bits_error             ),
  .io_in_0_d_ready                  (io_in_0_d_ready                  ),
  .io_in_0_d_valid                  (io_in_0_d_valid                  ),
  .io_in_0_d_bits_opcode            (io_in_0_d_bits_opcode            ),
  .io_in_0_d_bits_param             (io_in_0_d_bits_param             ),
  .io_in_0_d_bits_size              (io_in_0_d_bits_size              ),
  .io_in_0_d_bits_source            (io_in_0_d_bits_source            ),
  .io_in_0_d_bits_sink              (io_in_0_d_bits_sink              ),
  .io_in_0_d_bits_addr_lo           (io_in_0_d_bits_addr_lo           ),
  .io_in_0_d_bits_data              (io_in_0_d_bits_data              ),
  .io_in_0_d_bits_error             (io_in_0_d_bits_error             ),
  .io_in_0_e_ready                  (io_in_0_e_ready                  ),
  .io_in_0_e_valid                  (io_in_0_e_valid                  ),
  .io_in_0_e_bits_sink              (io_in_0_e_bits_sink              ),

  .io_interrupts_0_0               (gpio_irq_0),
  .io_interrupts_0_1               (gpio_irq_1),
  .io_interrupts_0_2               (gpio_irq_2),
  .io_interrupts_0_3               (gpio_irq_3),
  .io_interrupts_0_4               (gpio_irq_4),
  .io_interrupts_0_5               (gpio_irq_5),
  .io_interrupts_0_6               (gpio_irq_6),
  .io_interrupts_0_7               (gpio_irq_7),
  .io_interrupts_0_8               (gpio_irq_8),
  .io_interrupts_0_9               (gpio_irq_9),
  .io_interrupts_0_10              (gpio_irq_10),
  .io_interrupts_0_11              (gpio_irq_11),
  .io_interrupts_0_12              (gpio_irq_12),
  .io_interrupts_0_13              (gpio_irq_13),
  .io_interrupts_0_14              (gpio_irq_14),
  .io_interrupts_0_15              (gpio_irq_15),
  .io_interrupts_0_16              (gpio_irq_16),
  .io_interrupts_0_17              (gpio_irq_17),
  .io_interrupts_0_18              (gpio_irq_18),
  .io_interrupts_0_19              (gpio_irq_19),
  .io_interrupts_0_20              (gpio_irq_20),
  .io_interrupts_0_21              (gpio_irq_21),
  .io_interrupts_0_22              (gpio_irq_22),
  .io_interrupts_0_23              (gpio_irq_23),
  .io_interrupts_0_24              (gpio_irq_24),
  .io_interrupts_0_25              (gpio_irq_25),
  .io_interrupts_0_26              (gpio_irq_26),
  .io_interrupts_0_27              (gpio_irq_27),
  .io_interrupts_0_28              (gpio_irq_28),
  .io_interrupts_0_29              (gpio_irq_29),
  .io_interrupts_0_30              (gpio_irq_30),
  .io_interrupts_0_31              (gpio_irq_31),
 
  .io_port_pins_0_i_ival           (io_port_pins_0_i_ival),
  .io_port_pins_0_o_oval           (io_port_pins_0_o_oval),
  .io_port_pins_0_o_oe             (io_port_pins_0_o_oe),
  .io_port_pins_0_o_ie             (io_port_pins_0_o_ie),
  .io_port_pins_0_o_pue            (io_port_pins_0_o_pue),
  .io_port_pins_0_o_ds             (io_port_pins_0_o_ds),
  .io_port_pins_1_i_ival           (io_port_pins_1_i_ival),
  .io_port_pins_1_o_oval           (io_port_pins_1_o_oval),
  .io_port_pins_1_o_oe             (io_port_pins_1_o_oe),
  .io_port_pins_1_o_ie             (io_port_pins_1_o_ie),
  .io_port_pins_1_o_pue            (io_port_pins_1_o_pue),
  .io_port_pins_1_o_ds             (io_port_pins_1_o_ds),
  .io_port_pins_2_i_ival           (io_port_pins_2_i_ival),
  .io_port_pins_2_o_oval           (io_port_pins_2_o_oval),
  .io_port_pins_2_o_oe             (io_port_pins_2_o_oe),
  .io_port_pins_2_o_ie             (io_port_pins_2_o_ie),
  .io_port_pins_2_o_pue            (io_port_pins_2_o_pue),
  .io_port_pins_2_o_ds             (io_port_pins_2_o_ds),
  .io_port_pins_3_i_ival           (io_port_pins_3_i_ival),
  .io_port_pins_3_o_oval           (io_port_pins_3_o_oval),
  .io_port_pins_3_o_oe             (io_port_pins_3_o_oe),
  .io_port_pins_3_o_ie             (io_port_pins_3_o_ie),
  .io_port_pins_3_o_pue            (io_port_pins_3_o_pue),
  .io_port_pins_3_o_ds             (io_port_pins_3_o_ds),
  .io_port_pins_4_i_ival           (io_port_pins_4_i_ival),
  .io_port_pins_4_o_oval           (io_port_pins_4_o_oval),
  .io_port_pins_4_o_oe             (io_port_pins_4_o_oe),
  .io_port_pins_4_o_ie             (io_port_pins_4_o_ie),
  .io_port_pins_4_o_pue            (io_port_pins_4_o_pue),
  .io_port_pins_4_o_ds             (io_port_pins_4_o_ds),
  .io_port_pins_5_i_ival           (io_port_pins_5_i_ival),
  .io_port_pins_5_o_oval           (io_port_pins_5_o_oval),
  .io_port_pins_5_o_oe             (io_port_pins_5_o_oe),
  .io_port_pins_5_o_ie             (io_port_pins_5_o_ie),
  .io_port_pins_5_o_pue            (io_port_pins_5_o_pue),
  .io_port_pins_5_o_ds             (io_port_pins_5_o_ds),
  .io_port_pins_6_i_ival           (io_port_pins_6_i_ival),
  .io_port_pins_6_o_oval           (io_port_pins_6_o_oval),
  .io_port_pins_6_o_oe             (io_port_pins_6_o_oe),
  .io_port_pins_6_o_ie             (io_port_pins_6_o_ie),
  .io_port_pins_6_o_pue            (io_port_pins_6_o_pue),
  .io_port_pins_6_o_ds             (io_port_pins_6_o_ds),
  .io_port_pins_7_i_ival           (io_port_pins_7_i_ival),
  .io_port_pins_7_o_oval           (io_port_pins_7_o_oval),
  .io_port_pins_7_o_oe             (io_port_pins_7_o_oe),
  .io_port_pins_7_o_ie             (io_port_pins_7_o_ie),
  .io_port_pins_7_o_pue            (io_port_pins_7_o_pue),
  .io_port_pins_7_o_ds             (io_port_pins_7_o_ds),
  .io_port_pins_8_i_ival           (io_port_pins_8_i_ival),
  .io_port_pins_8_o_oval           (io_port_pins_8_o_oval),
  .io_port_pins_8_o_oe             (io_port_pins_8_o_oe),
  .io_port_pins_8_o_ie             (io_port_pins_8_o_ie),
  .io_port_pins_8_o_pue            (io_port_pins_8_o_pue),
  .io_port_pins_8_o_ds             (io_port_pins_8_o_ds),
  .io_port_pins_9_i_ival           (io_port_pins_9_i_ival),
  .io_port_pins_9_o_oval           (io_port_pins_9_o_oval),
  .io_port_pins_9_o_oe             (io_port_pins_9_o_oe),
  .io_port_pins_9_o_ie             (io_port_pins_9_o_ie),
  .io_port_pins_9_o_pue            (io_port_pins_9_o_pue),
  .io_port_pins_9_o_ds             (io_port_pins_9_o_ds),
  .io_port_pins_10_i_ival          (io_port_pins_10_i_ival),
  .io_port_pins_10_o_oval          (io_port_pins_10_o_oval),
  .io_port_pins_10_o_oe            (io_port_pins_10_o_oe),
  .io_port_pins_10_o_ie            (io_port_pins_10_o_ie),
  .io_port_pins_10_o_pue           (io_port_pins_10_o_pue),
  .io_port_pins_10_o_ds            (io_port_pins_10_o_ds),
  .io_port_pins_11_i_ival          (io_port_pins_11_i_ival),
  .io_port_pins_11_o_oval          (io_port_pins_11_o_oval),
  .io_port_pins_11_o_oe            (io_port_pins_11_o_oe),
  .io_port_pins_11_o_ie            (io_port_pins_11_o_ie),
  .io_port_pins_11_o_pue           (io_port_pins_11_o_pue),
  .io_port_pins_11_o_ds            (io_port_pins_11_o_ds),
  .io_port_pins_12_i_ival          (io_port_pins_12_i_ival),
  .io_port_pins_12_o_oval          (io_port_pins_12_o_oval),
  .io_port_pins_12_o_oe            (io_port_pins_12_o_oe),
  .io_port_pins_12_o_ie            (io_port_pins_12_o_ie),
  .io_port_pins_12_o_pue           (io_port_pins_12_o_pue),
  .io_port_pins_12_o_ds            (io_port_pins_12_o_ds),
  .io_port_pins_13_i_ival          (io_port_pins_13_i_ival),
  .io_port_pins_13_o_oval          (io_port_pins_13_o_oval),
  .io_port_pins_13_o_oe            (io_port_pins_13_o_oe),
  .io_port_pins_13_o_ie            (io_port_pins_13_o_ie),
  .io_port_pins_13_o_pue           (io_port_pins_13_o_pue),
  .io_port_pins_13_o_ds            (io_port_pins_13_o_ds),
  .io_port_pins_14_i_ival          (io_port_pins_14_i_ival),
  .io_port_pins_14_o_oval          (io_port_pins_14_o_oval),
  .io_port_pins_14_o_oe            (io_port_pins_14_o_oe),
  .io_port_pins_14_o_ie            (io_port_pins_14_o_ie),
  .io_port_pins_14_o_pue           (io_port_pins_14_o_pue),
  .io_port_pins_14_o_ds            (io_port_pins_14_o_ds),
  .io_port_pins_15_i_ival          (io_port_pins_15_i_ival),
  .io_port_pins_15_o_oval          (io_port_pins_15_o_oval),
  .io_port_pins_15_o_oe            (io_port_pins_15_o_oe),
  .io_port_pins_15_o_ie            (io_port_pins_15_o_ie),
  .io_port_pins_15_o_pue           (io_port_pins_15_o_pue),
  .io_port_pins_15_o_ds            (io_port_pins_15_o_ds),
  .io_port_pins_16_i_ival          (io_port_pins_16_i_ival),
  .io_port_pins_16_o_oval          (io_port_pins_16_o_oval),
  .io_port_pins_16_o_oe            (io_port_pins_16_o_oe),
  .io_port_pins_16_o_ie            (io_port_pins_16_o_ie),
  .io_port_pins_16_o_pue           (io_port_pins_16_o_pue),
  .io_port_pins_16_o_ds            (io_port_pins_16_o_ds),
  .io_port_pins_17_i_ival          (io_port_pins_17_i_ival),
  .io_port_pins_17_o_oval          (io_port_pins_17_o_oval),
  .io_port_pins_17_o_oe            (io_port_pins_17_o_oe),
  .io_port_pins_17_o_ie            (io_port_pins_17_o_ie),
  .io_port_pins_17_o_pue           (io_port_pins_17_o_pue),
  .io_port_pins_17_o_ds            (io_port_pins_17_o_ds),
  .io_port_pins_18_i_ival          (io_port_pins_18_i_ival),
  .io_port_pins_18_o_oval          (io_port_pins_18_o_oval),
  .io_port_pins_18_o_oe            (io_port_pins_18_o_oe),
  .io_port_pins_18_o_ie            (io_port_pins_18_o_ie),
  .io_port_pins_18_o_pue           (io_port_pins_18_o_pue),
  .io_port_pins_18_o_ds            (io_port_pins_18_o_ds),
  .io_port_pins_19_i_ival          (io_port_pins_19_i_ival),
  .io_port_pins_19_o_oval          (io_port_pins_19_o_oval),
  .io_port_pins_19_o_oe            (io_port_pins_19_o_oe),
  .io_port_pins_19_o_ie            (io_port_pins_19_o_ie),
  .io_port_pins_19_o_pue           (io_port_pins_19_o_pue),
  .io_port_pins_19_o_ds            (io_port_pins_19_o_ds),
  .io_port_pins_20_i_ival          (io_port_pins_20_i_ival),
  .io_port_pins_20_o_oval          (io_port_pins_20_o_oval),
  .io_port_pins_20_o_oe            (io_port_pins_20_o_oe),
  .io_port_pins_20_o_ie            (io_port_pins_20_o_ie),
  .io_port_pins_20_o_pue           (io_port_pins_20_o_pue),
  .io_port_pins_20_o_ds            (io_port_pins_20_o_ds),
  .io_port_pins_21_i_ival          (io_port_pins_21_i_ival),
  .io_port_pins_21_o_oval          (io_port_pins_21_o_oval),
  .io_port_pins_21_o_oe            (io_port_pins_21_o_oe),
  .io_port_pins_21_o_ie            (io_port_pins_21_o_ie),
  .io_port_pins_21_o_pue           (io_port_pins_21_o_pue),
  .io_port_pins_21_o_ds            (io_port_pins_21_o_ds),
  .io_port_pins_22_i_ival          (io_port_pins_22_i_ival),
  .io_port_pins_22_o_oval          (io_port_pins_22_o_oval),
  .io_port_pins_22_o_oe            (io_port_pins_22_o_oe),
  .io_port_pins_22_o_ie            (io_port_pins_22_o_ie),
  .io_port_pins_22_o_pue           (io_port_pins_22_o_pue),
  .io_port_pins_22_o_ds            (io_port_pins_22_o_ds),
  .io_port_pins_23_i_ival          (io_port_pins_23_i_ival),
  .io_port_pins_23_o_oval          (io_port_pins_23_o_oval),
  .io_port_pins_23_o_oe            (io_port_pins_23_o_oe),
  .io_port_pins_23_o_ie            (io_port_pins_23_o_ie),
  .io_port_pins_23_o_pue           (io_port_pins_23_o_pue),
  .io_port_pins_23_o_ds            (io_port_pins_23_o_ds),
  .io_port_pins_24_i_ival          (io_port_pins_24_i_ival),
  .io_port_pins_24_o_oval          (io_port_pins_24_o_oval),
  .io_port_pins_24_o_oe            (io_port_pins_24_o_oe),
  .io_port_pins_24_o_ie            (io_port_pins_24_o_ie),
  .io_port_pins_24_o_pue           (io_port_pins_24_o_pue),
  .io_port_pins_24_o_ds            (io_port_pins_24_o_ds),
  .io_port_pins_25_i_ival          (io_port_pins_25_i_ival),
  .io_port_pins_25_o_oval          (io_port_pins_25_o_oval),
  .io_port_pins_25_o_oe            (io_port_pins_25_o_oe),
  .io_port_pins_25_o_ie            (io_port_pins_25_o_ie),
  .io_port_pins_25_o_pue           (io_port_pins_25_o_pue),
  .io_port_pins_25_o_ds            (io_port_pins_25_o_ds),
  .io_port_pins_26_i_ival          (io_port_pins_26_i_ival),
  .io_port_pins_26_o_oval          (io_port_pins_26_o_oval),
  .io_port_pins_26_o_oe            (io_port_pins_26_o_oe),
  .io_port_pins_26_o_ie            (io_port_pins_26_o_ie),
  .io_port_pins_26_o_pue           (io_port_pins_26_o_pue),
  .io_port_pins_26_o_ds            (io_port_pins_26_o_ds),
  .io_port_pins_27_i_ival          (io_port_pins_27_i_ival),
  .io_port_pins_27_o_oval          (io_port_pins_27_o_oval),
  .io_port_pins_27_o_oe            (io_port_pins_27_o_oe),
  .io_port_pins_27_o_ie            (io_port_pins_27_o_ie),
  .io_port_pins_27_o_pue           (io_port_pins_27_o_pue),
  .io_port_pins_27_o_ds            (io_port_pins_27_o_ds),
  .io_port_pins_28_i_ival          (io_port_pins_28_i_ival),
  .io_port_pins_28_o_oval          (io_port_pins_28_o_oval),
  .io_port_pins_28_o_oe            (io_port_pins_28_o_oe),
  .io_port_pins_28_o_ie            (io_port_pins_28_o_ie),
  .io_port_pins_28_o_pue           (io_port_pins_28_o_pue),
  .io_port_pins_28_o_ds            (io_port_pins_28_o_ds),
  .io_port_pins_29_i_ival          (io_port_pins_29_i_ival),
  .io_port_pins_29_o_oval          (io_port_pins_29_o_oval),
  .io_port_pins_29_o_oe            (io_port_pins_29_o_oe),
  .io_port_pins_29_o_ie            (io_port_pins_29_o_ie),
  .io_port_pins_29_o_pue           (io_port_pins_29_o_pue),
  .io_port_pins_29_o_ds            (io_port_pins_29_o_ds),
  .io_port_pins_30_i_ival          (io_port_pins_30_i_ival),
  .io_port_pins_30_o_oval          (io_port_pins_30_o_oval),
  .io_port_pins_30_o_oe            (io_port_pins_30_o_oe),
  .io_port_pins_30_o_ie            (io_port_pins_30_o_ie),
  .io_port_pins_30_o_pue           (io_port_pins_30_o_pue),
  .io_port_pins_30_o_ds            (io_port_pins_30_o_ds),
  .io_port_pins_31_i_ival          (io_port_pins_31_i_ival),
  .io_port_pins_31_o_oval          (io_port_pins_31_o_oval),
  .io_port_pins_31_o_oe            (io_port_pins_31_o_oe),
  .io_port_pins_31_o_ie            (io_port_pins_31_o_ie),
  .io_port_pins_31_o_pue           (io_port_pins_31_o_pue),
  .io_port_pins_31_o_ds            (io_port_pins_31_o_ds),
  .io_port_iof_0_0_i_ival          (io_port_iof_0_0_i_ival),
  .io_port_iof_0_0_o_oval          (io_port_iof_0_0_o_oval),
  .io_port_iof_0_0_o_oe            (io_port_iof_0_0_o_oe),
  .io_port_iof_0_0_o_ie            (io_port_iof_0_0_o_ie),
  .io_port_iof_0_0_o_valid         (io_port_iof_0_0_o_valid),
  .io_port_iof_0_1_i_ival          (io_port_iof_0_1_i_ival),
  .io_port_iof_0_1_o_oval          (io_port_iof_0_1_o_oval),
  .io_port_iof_0_1_o_oe            (io_port_iof_0_1_o_oe),
  .io_port_iof_0_1_o_ie            (io_port_iof_0_1_o_ie),
  .io_port_iof_0_1_o_valid         (io_port_iof_0_1_o_valid),
  .io_port_iof_0_2_i_ival          (io_port_iof_0_2_i_ival),
  .io_port_iof_0_2_o_oval          (io_port_iof_0_2_o_oval),
  .io_port_iof_0_2_o_oe            (io_port_iof_0_2_o_oe),
  .io_port_iof_0_2_o_ie            (io_port_iof_0_2_o_ie),
  .io_port_iof_0_2_o_valid         (io_port_iof_0_2_o_valid),
  .io_port_iof_0_3_i_ival          (io_port_iof_0_3_i_ival),
  .io_port_iof_0_3_o_oval          (io_port_iof_0_3_o_oval),
  .io_port_iof_0_3_o_oe            (io_port_iof_0_3_o_oe),
  .io_port_iof_0_3_o_ie            (io_port_iof_0_3_o_ie),
  .io_port_iof_0_3_o_valid         (io_port_iof_0_3_o_valid),
  .io_port_iof_0_4_i_ival          (io_port_iof_0_4_i_ival),
  .io_port_iof_0_4_o_oval          (io_port_iof_0_4_o_oval),
  .io_port_iof_0_4_o_oe            (io_port_iof_0_4_o_oe),
  .io_port_iof_0_4_o_ie            (io_port_iof_0_4_o_ie),
  .io_port_iof_0_4_o_valid         (io_port_iof_0_4_o_valid),
  .io_port_iof_0_5_i_ival          (io_port_iof_0_5_i_ival),
  .io_port_iof_0_5_o_oval          (io_port_iof_0_5_o_oval),
  .io_port_iof_0_5_o_oe            (io_port_iof_0_5_o_oe),
  .io_port_iof_0_5_o_ie            (io_port_iof_0_5_o_ie),
  .io_port_iof_0_5_o_valid         (io_port_iof_0_5_o_valid),
  .io_port_iof_0_6_i_ival          (io_port_iof_0_6_i_ival),
  .io_port_iof_0_6_o_oval          (io_port_iof_0_6_o_oval),
  .io_port_iof_0_6_o_oe            (io_port_iof_0_6_o_oe),
  .io_port_iof_0_6_o_ie            (io_port_iof_0_6_o_ie),
  .io_port_iof_0_6_o_valid         (io_port_iof_0_6_o_valid),
  .io_port_iof_0_7_i_ival          (io_port_iof_0_7_i_ival),
  .io_port_iof_0_7_o_oval          (io_port_iof_0_7_o_oval),
  .io_port_iof_0_7_o_oe            (io_port_iof_0_7_o_oe),
  .io_port_iof_0_7_o_ie            (io_port_iof_0_7_o_ie),
  .io_port_iof_0_7_o_valid         (io_port_iof_0_7_o_valid),
  .io_port_iof_0_8_i_ival          (io_port_iof_0_8_i_ival),
  .io_port_iof_0_8_o_oval          (io_port_iof_0_8_o_oval),
  .io_port_iof_0_8_o_oe            (io_port_iof_0_8_o_oe),
  .io_port_iof_0_8_o_ie            (io_port_iof_0_8_o_ie),
  .io_port_iof_0_8_o_valid         (io_port_iof_0_8_o_valid),
  .io_port_iof_0_9_i_ival          (io_port_iof_0_9_i_ival),
  .io_port_iof_0_9_o_oval          (io_port_iof_0_9_o_oval),
  .io_port_iof_0_9_o_oe            (io_port_iof_0_9_o_oe),
  .io_port_iof_0_9_o_ie            (io_port_iof_0_9_o_ie),
  .io_port_iof_0_9_o_valid         (io_port_iof_0_9_o_valid),
  .io_port_iof_0_10_i_ival         (io_port_iof_0_10_i_ival),
  .io_port_iof_0_10_o_oval         (io_port_iof_0_10_o_oval),
  .io_port_iof_0_10_o_oe           (io_port_iof_0_10_o_oe),
  .io_port_iof_0_10_o_ie           (io_port_iof_0_10_o_ie),
  .io_port_iof_0_10_o_valid        (io_port_iof_0_10_o_valid),
  .io_port_iof_0_11_i_ival         (io_port_iof_0_11_i_ival),
  .io_port_iof_0_11_o_oval         (io_port_iof_0_11_o_oval),
  .io_port_iof_0_11_o_oe           (io_port_iof_0_11_o_oe),
  .io_port_iof_0_11_o_ie           (io_port_iof_0_11_o_ie),
  .io_port_iof_0_11_o_valid        (io_port_iof_0_11_o_valid),
  .io_port_iof_0_12_i_ival         (io_port_iof_0_12_i_ival),
  .io_port_iof_0_12_o_oval         (io_port_iof_0_12_o_oval),
  .io_port_iof_0_12_o_oe           (io_port_iof_0_12_o_oe),
  .io_port_iof_0_12_o_ie           (io_port_iof_0_12_o_ie),
  .io_port_iof_0_12_o_valid        (io_port_iof_0_12_o_valid),
  .io_port_iof_0_13_i_ival         (io_port_iof_0_13_i_ival),
  .io_port_iof_0_13_o_oval         (io_port_iof_0_13_o_oval),
  .io_port_iof_0_13_o_oe           (io_port_iof_0_13_o_oe),
  .io_port_iof_0_13_o_ie           (io_port_iof_0_13_o_ie),
  .io_port_iof_0_13_o_valid        (io_port_iof_0_13_o_valid),
  .io_port_iof_0_14_i_ival         (io_port_iof_0_14_i_ival),
  .io_port_iof_0_14_o_oval         (io_port_iof_0_14_o_oval),
  .io_port_iof_0_14_o_oe           (io_port_iof_0_14_o_oe),
  .io_port_iof_0_14_o_ie           (io_port_iof_0_14_o_ie),
  .io_port_iof_0_14_o_valid        (io_port_iof_0_14_o_valid),
  .io_port_iof_0_15_i_ival         (io_port_iof_0_15_i_ival),
  .io_port_iof_0_15_o_oval         (io_port_iof_0_15_o_oval),
  .io_port_iof_0_15_o_oe           (io_port_iof_0_15_o_oe),
  .io_port_iof_0_15_o_ie           (io_port_iof_0_15_o_ie),
  .io_port_iof_0_15_o_valid        (io_port_iof_0_15_o_valid),
  .io_port_iof_0_16_i_ival         (io_port_iof_0_16_i_ival),
  .io_port_iof_0_16_o_oval         (io_port_iof_0_16_o_oval),
  .io_port_iof_0_16_o_oe           (io_port_iof_0_16_o_oe),
  .io_port_iof_0_16_o_ie           (io_port_iof_0_16_o_ie),
  .io_port_iof_0_16_o_valid        (io_port_iof_0_16_o_valid),
  .io_port_iof_0_17_i_ival         (io_port_iof_0_17_i_ival),
  .io_port_iof_0_17_o_oval         (io_port_iof_0_17_o_oval),
  .io_port_iof_0_17_o_oe           (io_port_iof_0_17_o_oe),
  .io_port_iof_0_17_o_ie           (io_port_iof_0_17_o_ie),
  .io_port_iof_0_17_o_valid        (io_port_iof_0_17_o_valid),
  .io_port_iof_0_18_i_ival         (io_port_iof_0_18_i_ival),
  .io_port_iof_0_18_o_oval         (io_port_iof_0_18_o_oval),
  .io_port_iof_0_18_o_oe           (io_port_iof_0_18_o_oe),
  .io_port_iof_0_18_o_ie           (io_port_iof_0_18_o_ie),
  .io_port_iof_0_18_o_valid        (io_port_iof_0_18_o_valid),
  .io_port_iof_0_19_i_ival         (io_port_iof_0_19_i_ival),
  .io_port_iof_0_19_o_oval         (io_port_iof_0_19_o_oval),
  .io_port_iof_0_19_o_oe           (io_port_iof_0_19_o_oe),
  .io_port_iof_0_19_o_ie           (io_port_iof_0_19_o_ie),
  .io_port_iof_0_19_o_valid        (io_port_iof_0_19_o_valid),
  .io_port_iof_0_20_i_ival         (io_port_iof_0_20_i_ival),
  .io_port_iof_0_20_o_oval         (io_port_iof_0_20_o_oval),
  .io_port_iof_0_20_o_oe           (io_port_iof_0_20_o_oe),
  .io_port_iof_0_20_o_ie           (io_port_iof_0_20_o_ie),
  .io_port_iof_0_20_o_valid        (io_port_iof_0_20_o_valid),
  .io_port_iof_0_21_i_ival         (io_port_iof_0_21_i_ival),
  .io_port_iof_0_21_o_oval         (io_port_iof_0_21_o_oval),
  .io_port_iof_0_21_o_oe           (io_port_iof_0_21_o_oe),
  .io_port_iof_0_21_o_ie           (io_port_iof_0_21_o_ie),
  .io_port_iof_0_21_o_valid        (io_port_iof_0_21_o_valid),
  .io_port_iof_0_22_i_ival         (io_port_iof_0_22_i_ival),
  .io_port_iof_0_22_o_oval         (io_port_iof_0_22_o_oval),
  .io_port_iof_0_22_o_oe           (io_port_iof_0_22_o_oe),
  .io_port_iof_0_22_o_ie           (io_port_iof_0_22_o_ie),
  .io_port_iof_0_22_o_valid        (io_port_iof_0_22_o_valid),
  .io_port_iof_0_23_i_ival         (io_port_iof_0_23_i_ival),
  .io_port_iof_0_23_o_oval         (io_port_iof_0_23_o_oval),
  .io_port_iof_0_23_o_oe           (io_port_iof_0_23_o_oe),
  .io_port_iof_0_23_o_ie           (io_port_iof_0_23_o_ie),
  .io_port_iof_0_23_o_valid        (io_port_iof_0_23_o_valid),
  .io_port_iof_0_24_i_ival         (io_port_iof_0_24_i_ival),
  .io_port_iof_0_24_o_oval         (io_port_iof_0_24_o_oval),
  .io_port_iof_0_24_o_oe           (io_port_iof_0_24_o_oe),
  .io_port_iof_0_24_o_ie           (io_port_iof_0_24_o_ie),
  .io_port_iof_0_24_o_valid        (io_port_iof_0_24_o_valid),
  .io_port_iof_0_25_i_ival         (io_port_iof_0_25_i_ival),
  .io_port_iof_0_25_o_oval         (io_port_iof_0_25_o_oval),
  .io_port_iof_0_25_o_oe           (io_port_iof_0_25_o_oe),
  .io_port_iof_0_25_o_ie           (io_port_iof_0_25_o_ie),
  .io_port_iof_0_25_o_valid        (io_port_iof_0_25_o_valid),
  .io_port_iof_0_26_i_ival         (io_port_iof_0_26_i_ival),
  .io_port_iof_0_26_o_oval         (io_port_iof_0_26_o_oval),
  .io_port_iof_0_26_o_oe           (io_port_iof_0_26_o_oe),
  .io_port_iof_0_26_o_ie           (io_port_iof_0_26_o_ie),
  .io_port_iof_0_26_o_valid        (io_port_iof_0_26_o_valid),
  .io_port_iof_0_27_i_ival         (io_port_iof_0_27_i_ival),
  .io_port_iof_0_27_o_oval         (io_port_iof_0_27_o_oval),
  .io_port_iof_0_27_o_oe           (io_port_iof_0_27_o_oe),
  .io_port_iof_0_27_o_ie           (io_port_iof_0_27_o_ie),
  .io_port_iof_0_27_o_valid        (io_port_iof_0_27_o_valid),
  .io_port_iof_0_28_i_ival         (io_port_iof_0_28_i_ival),
  .io_port_iof_0_28_o_oval         (io_port_iof_0_28_o_oval),
  .io_port_iof_0_28_o_oe           (io_port_iof_0_28_o_oe),
  .io_port_iof_0_28_o_ie           (io_port_iof_0_28_o_ie),
  .io_port_iof_0_28_o_valid        (io_port_iof_0_28_o_valid),
  .io_port_iof_0_29_i_ival         (io_port_iof_0_29_i_ival),
  .io_port_iof_0_29_o_oval         (io_port_iof_0_29_o_oval),
  .io_port_iof_0_29_o_oe           (io_port_iof_0_29_o_oe),
  .io_port_iof_0_29_o_ie           (io_port_iof_0_29_o_ie),
  .io_port_iof_0_29_o_valid        (io_port_iof_0_29_o_valid),
  .io_port_iof_0_30_i_ival         (io_port_iof_0_30_i_ival),
  .io_port_iof_0_30_o_oval         (io_port_iof_0_30_o_oval),
  .io_port_iof_0_30_o_oe           (io_port_iof_0_30_o_oe),
  .io_port_iof_0_30_o_ie           (io_port_iof_0_30_o_ie),
  .io_port_iof_0_30_o_valid        (io_port_iof_0_30_o_valid),
  .io_port_iof_0_31_i_ival         (io_port_iof_0_31_i_ival),
  .io_port_iof_0_31_o_oval         (io_port_iof_0_31_o_oval),
  .io_port_iof_0_31_o_oe           (io_port_iof_0_31_o_oe),
  .io_port_iof_0_31_o_ie           (io_port_iof_0_31_o_ie),
  .io_port_iof_0_31_o_valid        (io_port_iof_0_31_o_valid),
  .io_port_iof_1_0_i_ival          (io_port_iof_1_0_i_ival),
  .io_port_iof_1_0_o_oval          (io_port_iof_1_0_o_oval),
  .io_port_iof_1_0_o_oe            (io_port_iof_1_0_o_oe),
  .io_port_iof_1_0_o_ie            (io_port_iof_1_0_o_ie),
  .io_port_iof_1_0_o_valid         (io_port_iof_1_0_o_valid),
  .io_port_iof_1_1_i_ival          (io_port_iof_1_1_i_ival),
  .io_port_iof_1_1_o_oval          (io_port_iof_1_1_o_oval),
  .io_port_iof_1_1_o_oe            (io_port_iof_1_1_o_oe),
  .io_port_iof_1_1_o_ie            (io_port_iof_1_1_o_ie),
  .io_port_iof_1_1_o_valid         (io_port_iof_1_1_o_valid),
  .io_port_iof_1_2_i_ival          (io_port_iof_1_2_i_ival),
  .io_port_iof_1_2_o_oval          (io_port_iof_1_2_o_oval),
  .io_port_iof_1_2_o_oe            (io_port_iof_1_2_o_oe),
  .io_port_iof_1_2_o_ie            (io_port_iof_1_2_o_ie),
  .io_port_iof_1_2_o_valid         (io_port_iof_1_2_o_valid),
  .io_port_iof_1_3_i_ival          (io_port_iof_1_3_i_ival),
  .io_port_iof_1_3_o_oval          (io_port_iof_1_3_o_oval),
  .io_port_iof_1_3_o_oe            (io_port_iof_1_3_o_oe),
  .io_port_iof_1_3_o_ie            (io_port_iof_1_3_o_ie),
  .io_port_iof_1_3_o_valid         (io_port_iof_1_3_o_valid),
  .io_port_iof_1_4_i_ival          (io_port_iof_1_4_i_ival),
  .io_port_iof_1_4_o_oval          (io_port_iof_1_4_o_oval),
  .io_port_iof_1_4_o_oe            (io_port_iof_1_4_o_oe),
  .io_port_iof_1_4_o_ie            (io_port_iof_1_4_o_ie),
  .io_port_iof_1_4_o_valid         (io_port_iof_1_4_o_valid),
  .io_port_iof_1_5_i_ival          (io_port_iof_1_5_i_ival),
  .io_port_iof_1_5_o_oval          (io_port_iof_1_5_o_oval),
  .io_port_iof_1_5_o_oe            (io_port_iof_1_5_o_oe),
  .io_port_iof_1_5_o_ie            (io_port_iof_1_5_o_ie),
  .io_port_iof_1_5_o_valid         (io_port_iof_1_5_o_valid),
  .io_port_iof_1_6_i_ival          (io_port_iof_1_6_i_ival),
  .io_port_iof_1_6_o_oval          (io_port_iof_1_6_o_oval),
  .io_port_iof_1_6_o_oe            (io_port_iof_1_6_o_oe),
  .io_port_iof_1_6_o_ie            (io_port_iof_1_6_o_ie),
  .io_port_iof_1_6_o_valid         (io_port_iof_1_6_o_valid),
  .io_port_iof_1_7_i_ival          (io_port_iof_1_7_i_ival),
  .io_port_iof_1_7_o_oval          (io_port_iof_1_7_o_oval),
  .io_port_iof_1_7_o_oe            (io_port_iof_1_7_o_oe),
  .io_port_iof_1_7_o_ie            (io_port_iof_1_7_o_ie),
  .io_port_iof_1_7_o_valid         (io_port_iof_1_7_o_valid),
  .io_port_iof_1_8_i_ival          (io_port_iof_1_8_i_ival),
  .io_port_iof_1_8_o_oval          (io_port_iof_1_8_o_oval),
  .io_port_iof_1_8_o_oe            (io_port_iof_1_8_o_oe),
  .io_port_iof_1_8_o_ie            (io_port_iof_1_8_o_ie),
  .io_port_iof_1_8_o_valid         (io_port_iof_1_8_o_valid),
  .io_port_iof_1_9_i_ival          (io_port_iof_1_9_i_ival),
  .io_port_iof_1_9_o_oval          (io_port_iof_1_9_o_oval),
  .io_port_iof_1_9_o_oe            (io_port_iof_1_9_o_oe),
  .io_port_iof_1_9_o_ie            (io_port_iof_1_9_o_ie),
  .io_port_iof_1_9_o_valid         (io_port_iof_1_9_o_valid),
  .io_port_iof_1_10_i_ival         (io_port_iof_1_10_i_ival),
  .io_port_iof_1_10_o_oval         (io_port_iof_1_10_o_oval),
  .io_port_iof_1_10_o_oe           (io_port_iof_1_10_o_oe),
  .io_port_iof_1_10_o_ie           (io_port_iof_1_10_o_ie),
  .io_port_iof_1_10_o_valid        (io_port_iof_1_10_o_valid),
  .io_port_iof_1_11_i_ival         (io_port_iof_1_11_i_ival),
  .io_port_iof_1_11_o_oval         (io_port_iof_1_11_o_oval),
  .io_port_iof_1_11_o_oe           (io_port_iof_1_11_o_oe),
  .io_port_iof_1_11_o_ie           (io_port_iof_1_11_o_ie),
  .io_port_iof_1_11_o_valid        (io_port_iof_1_11_o_valid),
  .io_port_iof_1_12_i_ival         (io_port_iof_1_12_i_ival),
  .io_port_iof_1_12_o_oval         (io_port_iof_1_12_o_oval),
  .io_port_iof_1_12_o_oe           (io_port_iof_1_12_o_oe),
  .io_port_iof_1_12_o_ie           (io_port_iof_1_12_o_ie),
  .io_port_iof_1_12_o_valid        (io_port_iof_1_12_o_valid),
  .io_port_iof_1_13_i_ival         (io_port_iof_1_13_i_ival),
  .io_port_iof_1_13_o_oval         (io_port_iof_1_13_o_oval),
  .io_port_iof_1_13_o_oe           (io_port_iof_1_13_o_oe),
  .io_port_iof_1_13_o_ie           (io_port_iof_1_13_o_ie),
  .io_port_iof_1_13_o_valid        (io_port_iof_1_13_o_valid),
  .io_port_iof_1_14_i_ival         (io_port_iof_1_14_i_ival),
  .io_port_iof_1_14_o_oval         (io_port_iof_1_14_o_oval),
  .io_port_iof_1_14_o_oe           (io_port_iof_1_14_o_oe),
  .io_port_iof_1_14_o_ie           (io_port_iof_1_14_o_ie),
  .io_port_iof_1_14_o_valid        (io_port_iof_1_14_o_valid),
  .io_port_iof_1_15_i_ival         (io_port_iof_1_15_i_ival),
  .io_port_iof_1_15_o_oval         (io_port_iof_1_15_o_oval),
  .io_port_iof_1_15_o_oe           (io_port_iof_1_15_o_oe),
  .io_port_iof_1_15_o_ie           (io_port_iof_1_15_o_ie),
  .io_port_iof_1_15_o_valid        (io_port_iof_1_15_o_valid),
  .io_port_iof_1_16_i_ival         (io_port_iof_1_16_i_ival),
  .io_port_iof_1_16_o_oval         (io_port_iof_1_16_o_oval),
  .io_port_iof_1_16_o_oe           (io_port_iof_1_16_o_oe),
  .io_port_iof_1_16_o_ie           (io_port_iof_1_16_o_ie),
  .io_port_iof_1_16_o_valid        (io_port_iof_1_16_o_valid),
  .io_port_iof_1_17_i_ival         (io_port_iof_1_17_i_ival),
  .io_port_iof_1_17_o_oval         (io_port_iof_1_17_o_oval),
  .io_port_iof_1_17_o_oe           (io_port_iof_1_17_o_oe),
  .io_port_iof_1_17_o_ie           (io_port_iof_1_17_o_ie),
  .io_port_iof_1_17_o_valid        (io_port_iof_1_17_o_valid),
  .io_port_iof_1_18_i_ival         (io_port_iof_1_18_i_ival),
  .io_port_iof_1_18_o_oval         (io_port_iof_1_18_o_oval),
  .io_port_iof_1_18_o_oe           (io_port_iof_1_18_o_oe),
  .io_port_iof_1_18_o_ie           (io_port_iof_1_18_o_ie),
  .io_port_iof_1_18_o_valid        (io_port_iof_1_18_o_valid),
  .io_port_iof_1_19_i_ival         (io_port_iof_1_19_i_ival),
  .io_port_iof_1_19_o_oval         (io_port_iof_1_19_o_oval),
  .io_port_iof_1_19_o_oe           (io_port_iof_1_19_o_oe),
  .io_port_iof_1_19_o_ie           (io_port_iof_1_19_o_ie),
  .io_port_iof_1_19_o_valid        (io_port_iof_1_19_o_valid),
  .io_port_iof_1_20_i_ival         (io_port_iof_1_20_i_ival),
  .io_port_iof_1_20_o_oval         (io_port_iof_1_20_o_oval),
  .io_port_iof_1_20_o_oe           (io_port_iof_1_20_o_oe),
  .io_port_iof_1_20_o_ie           (io_port_iof_1_20_o_ie),
  .io_port_iof_1_20_o_valid        (io_port_iof_1_20_o_valid),
  .io_port_iof_1_21_i_ival         (io_port_iof_1_21_i_ival),
  .io_port_iof_1_21_o_oval         (io_port_iof_1_21_o_oval),
  .io_port_iof_1_21_o_oe           (io_port_iof_1_21_o_oe),
  .io_port_iof_1_21_o_ie           (io_port_iof_1_21_o_ie),
  .io_port_iof_1_21_o_valid        (io_port_iof_1_21_o_valid),
  .io_port_iof_1_22_i_ival         (io_port_iof_1_22_i_ival),
  .io_port_iof_1_22_o_oval         (io_port_iof_1_22_o_oval),
  .io_port_iof_1_22_o_oe           (io_port_iof_1_22_o_oe),
  .io_port_iof_1_22_o_ie           (io_port_iof_1_22_o_ie),
  .io_port_iof_1_22_o_valid        (io_port_iof_1_22_o_valid),
  .io_port_iof_1_23_i_ival         (io_port_iof_1_23_i_ival),
  .io_port_iof_1_23_o_oval         (io_port_iof_1_23_o_oval),
  .io_port_iof_1_23_o_oe           (io_port_iof_1_23_o_oe),
  .io_port_iof_1_23_o_ie           (io_port_iof_1_23_o_ie),
  .io_port_iof_1_23_o_valid        (io_port_iof_1_23_o_valid),
  .io_port_iof_1_24_i_ival         (io_port_iof_1_24_i_ival),
  .io_port_iof_1_24_o_oval         (io_port_iof_1_24_o_oval),
  .io_port_iof_1_24_o_oe           (io_port_iof_1_24_o_oe),
  .io_port_iof_1_24_o_ie           (io_port_iof_1_24_o_ie),
  .io_port_iof_1_24_o_valid        (io_port_iof_1_24_o_valid),
  .io_port_iof_1_25_i_ival         (io_port_iof_1_25_i_ival),
  .io_port_iof_1_25_o_oval         (io_port_iof_1_25_o_oval),
  .io_port_iof_1_25_o_oe           (io_port_iof_1_25_o_oe),
  .io_port_iof_1_25_o_ie           (io_port_iof_1_25_o_ie),
  .io_port_iof_1_25_o_valid        (io_port_iof_1_25_o_valid),
  .io_port_iof_1_26_i_ival         (io_port_iof_1_26_i_ival),
  .io_port_iof_1_26_o_oval         (io_port_iof_1_26_o_oval),
  .io_port_iof_1_26_o_oe           (io_port_iof_1_26_o_oe),
  .io_port_iof_1_26_o_ie           (io_port_iof_1_26_o_ie),
  .io_port_iof_1_26_o_valid        (io_port_iof_1_26_o_valid),
  .io_port_iof_1_27_i_ival         (io_port_iof_1_27_i_ival),
  .io_port_iof_1_27_o_oval         (io_port_iof_1_27_o_oval),
  .io_port_iof_1_27_o_oe           (io_port_iof_1_27_o_oe),
  .io_port_iof_1_27_o_ie           (io_port_iof_1_27_o_ie),
  .io_port_iof_1_27_o_valid        (io_port_iof_1_27_o_valid),
  .io_port_iof_1_28_i_ival         (io_port_iof_1_28_i_ival),
  .io_port_iof_1_28_o_oval         (io_port_iof_1_28_o_oval),
  .io_port_iof_1_28_o_oe           (io_port_iof_1_28_o_oe),
  .io_port_iof_1_28_o_ie           (io_port_iof_1_28_o_ie),
  .io_port_iof_1_28_o_valid        (io_port_iof_1_28_o_valid),
  .io_port_iof_1_29_i_ival         (io_port_iof_1_29_i_ival),
  .io_port_iof_1_29_o_oval         (io_port_iof_1_29_o_oval),
  .io_port_iof_1_29_o_oe           (io_port_iof_1_29_o_oe),
  .io_port_iof_1_29_o_ie           (io_port_iof_1_29_o_ie),
  .io_port_iof_1_29_o_valid        (io_port_iof_1_29_o_valid),
  .io_port_iof_1_30_i_ival         (io_port_iof_1_30_i_ival),
  .io_port_iof_1_30_o_oval         (io_port_iof_1_30_o_oval),
  .io_port_iof_1_30_o_oe           (io_port_iof_1_30_o_oe),
  .io_port_iof_1_30_o_ie           (io_port_iof_1_30_o_ie),
  .io_port_iof_1_30_o_valid        (io_port_iof_1_30_o_valid),
  .io_port_iof_1_31_i_ival         (io_port_iof_1_31_i_ival),
  .io_port_iof_1_31_o_oval         (io_port_iof_1_31_o_oval),
  .io_port_iof_1_31_o_oe           (io_port_iof_1_31_o_oe),
  .io_port_iof_1_31_o_ie           (io_port_iof_1_31_o_ie),
  .io_port_iof_1_31_o_valid        (io_port_iof_1_31_o_valid)
);

endmodule
