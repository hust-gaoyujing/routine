`default_nettype none

module gs_filter_5x5(




);





endmodule