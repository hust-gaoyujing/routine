 /*                                                                      
  *  Copyright (c) 2018-2020 Nuclei System Technology, Inc.              
  *  All rights reserved.                                                
  */                                                                     

























module ux607_core (


  
  
  input  jtag_TCK    ,
  input  jtag_TMS    ,
  input  jtag_TDI    ,
  output jtag_TDO    ,
  output jtag_DRV_TDO,

      
      
  output hart_halted,
  input  i_dbg_stop,    
  input  override_dm_sleep,    


  output sysrstreq,

  output trace_ivalid,
  output trace_iexception, 
  output trace_interrupt, 
  output [64-1:0] trace_cause, 
  output [64-1:0] trace_tval, 
  output [64-1:0] trace_iaddr, 
  output [32-1:0] trace_instr, 
  output [1:0] trace_priv, 
  output trace_bjp_taken,
  output trace_dmode,









  input  core_clk_aon,






  input  core_clk,



  input  core_reset_n,



  input  por_reset_n,


  input reset_bypass,

  input clkgate_bypass, 




  input  nmi,








  
      
  input  mtime_toggle_a,


      
      
  input  dbg_toggle_a,
     

  
      
      
  input [32-1:0] irq_i,






  output                        ilm_cs,  
  output [13-1:0] ilm_addr, 
  output [8-1:0] ilm_byte_we,
  output [64-1:0] ilm_wdata,          
  input  [64-1:0] ilm_rdata,
  output                        clk_ilm_ram,
  
 
 
 
 
 
 
 
 
 

 
 
 
 
 
 


  
  input                             mem_arready,
  output                            mem_arvalid,
  
  output [32-1:0]      mem_araddr,
  output [7:0]                      mem_arlen,
  output [2:0]                      mem_arsize,
  output [1:0]                      mem_arburst,
  output [1:0]                      mem_arlock,
  output [3:0]                      mem_arcache,
  output [2:0]                      mem_arprot,
  
  
  
  
  input                             mem_awready,
  output                            mem_awvalid,
  
  output [32-1:0]      mem_awaddr,
  output [7:0]                      mem_awlen,
  output [2:0]                      mem_awsize,
  output [1:0]                      mem_awburst,
  output [1:0]                      mem_awlock,
  output [3:0]                      mem_awcache,
  output [2:0]                      mem_awprot,
  
  
  

  input                             mem_wready,
  output                            mem_wvalid,
  
  output [64-1:0]           mem_wdata,
  output [8-1:0]        mem_wstrb,
  output                            mem_wlast,
  
  output                            mem_rready,
  input                             mem_rvalid,
  
  input [64-1:0]            mem_rdata,
  input [1:0]                       mem_rresp,
  input                             mem_rlast,
  
  output                            mem_bready,
  input                             mem_bvalid,
  
  input [1:0]                       mem_bresp,

  input                            mem_clk_en,




  
  
  
  
  
  
  
  
  output                        dlm0_cs,  
  output [13-1:0] dlm0_addr, 
  output [4-1:0] dlm0_byte_we,
  output [32-1:0] dlm0_wdata,          
  input  [32-1:0] dlm0_rdata,
  output                        clk_dlm0_ram,

  output                        dlm1_cs,  
  output [13-1:0] dlm1_addr, 
  output [4-1:0] dlm1_byte_we,
  output [32-1:0] dlm1_wdata,          
  input  [32-1:0] dlm1_rdata,
  output                        clk_dlm1_ram,
  

  
  
  
  
  
  
  
  
  
  
  
  
  

  
  
  
  
  
  

    
  input                            icache_disable_init,

  output                           icache_tag0_cs,  
  output                           icache_tag0_we,  
  output [7-1:0] icache_tag0_addr, 
  output [54-1:0] icache_tag0_wdata,          
  input  [54-1:0] icache_tag0_rdata,
  output                               clk_icache_tag0,

  output                           icache_data0_cs,  
  output                           icache_data0_we,  
  output [9-1:0] icache_data0_addr, 
  output [64-1:0] icache_data0_wdata,          
  input  [64-1:0] icache_data0_rdata,
  output                               clk_icache_data0,

  output                           icache_tag1_cs,  
  output                           icache_tag1_we,  
  output [7-1:0] icache_tag1_addr, 
  output [54-1:0] icache_tag1_wdata,          
  input  [54-1:0] icache_tag1_rdata,
  output                               clk_icache_tag1,

  
  output                           icache_data1_cs,  
  output                           icache_data1_we,  
  output [9-1:0] icache_data1_addr, 
  output [64-1:0] icache_data1_wdata,          
  input  [64-1:0] icache_data1_rdata,
  output                               clk_icache_data1,





  input  dcache_disable_init,
   
  output                          clk_dcache_w0_tram,  
  output                          dcache_w0_tram_cs,  
  output [6-1:0]  dcache_w0_tram_addr,
  output                          dcache_w0_tram_we ,
  output [24-1:0]  dcache_w0_tram_din,          
  input  [24-1:0]  dcache_w0_tram_dout,
   
  output                          clk_dcache_w1_tram,  
  output                          dcache_w1_tram_cs,  
  output [6-1:0]  dcache_w1_tram_addr, 
  output                          dcache_w1_tram_we ,
  output [24-1:0]  dcache_w1_tram_din,          
  input  [24-1:0]  dcache_w1_tram_dout,


  
  
  output                          clk_dcache_dram_b0,  
  output                          dcache_dram_b0_cs,  
  output [8-1:0] dcache_dram_b0_addr, 
  output [4-1:0] dcache_dram_b0_wem,
  output [32-1:0] dcache_dram_b0_din,          
  input  [32-1:0] dcache_dram_b0_dout,
                                                
  output                          clk_dcache_dram_b1,  
  output                          dcache_dram_b1_cs,  
  output [8-1:0] dcache_dram_b1_addr, 
  output [4-1:0] dcache_dram_b1_wem,
  output [32-1:0] dcache_dram_b1_din,          
  input  [32-1:0] dcache_dram_b1_dout,
                                                
  output                          clk_dcache_dram_b2,  
  output                          dcache_dram_b2_cs,  
  output [8-1:0] dcache_dram_b2_addr, 
  output [4-1:0] dcache_dram_b2_wem,
  output [32-1:0] dcache_dram_b2_din,          
  input  [32-1:0] dcache_dram_b2_dout,
                                                
  output                          clk_dcache_dram_b3,  
  output                          dcache_dram_b3_cs,  
  output [8-1:0] dcache_dram_b3_addr, 
  output [4-1:0] dcache_dram_b3_wem,
  output [32-1:0] dcache_dram_b3_din,          
  input  [32-1:0] dcache_dram_b3_dout,

  input                                           mmu_tlb_disable_init,
  
  output                                          clk_mmu_tlb_way0, 
  output                                          clk_mmu_tlb_way1, 
  output                                          mmu_tlb_way0_cs, 
  output                                          mmu_tlb_way1_cs, 
  output                                          mmu_tlb_way0_we, 
  output                                          mmu_tlb_way1_we, 
  output [66-1:0]               mmu_tlb_way0_wdata, 
  output [66-1:0]               mmu_tlb_way1_wdata,
  output [6-1:0]              mmu_tlb_way0_addr, 
  output [6-1:0]              mmu_tlb_way1_addr, 
  input  [66-1:0]               mmu_tlb_way0_dout, 
  input  [66-1:0]               mmu_tlb_way1_dout, 



  
  
  
  

























  
  
  
  
 
 
 
 
 
 
 
 
 
 
 
 
 
 
 
 
 
 
 

  output [1:0]                   ppi_ahbl_htrans  ,  
  output                         ppi_ahbl_hwrite  ,  
  output [32-1:0]   ppi_ahbl_haddr   ,  
  output [2:0]                   ppi_ahbl_hsize   ,  
  output [32-1:0]        ppi_ahbl_hwdata  ,  
  output [3:0]                   ppi_ahbl_hprot   ,

  input  [32-1:0]        ppi_ahbl_hrdata  ,  
  input  [1:0]                   ppi_ahbl_hresp   ,  
  input                          ppi_ahbl_hready  ,  

  input                          ppi_ahbl_clk_en, 










  output tx_evt,
  input  rx_evt,


  input  [64-1:0] hart_id,


  input  [64-1:0] reset_vector, 





  output core_wfi_mode, 


































































  output core_sleep_value

  );


  wire exu_i_valid;
  wire exu_i_ready;
  wire [64-1:0] x3;
  wire alu_cmt_i_valid;
  wire [64-1:0] alu_cmt_i_pc;
  wire mscratch_ena;
  wire [64-1:0] mscratch_nxt;
  wire sscratch_ena;
  wire [64-1:0] sscratch_nxt;

    localparam urjif1vu4pqgqxt4x8 = 51; 

  wire c4boo209;
  wire yukl2;

  wire zmxoq9ga;
  wire mtip;
  wire msip;

  assign zmxoq9ga = 1'b0 
                | msip
                ;

  wire x_cq40qmp6a;
  wire uc5qxb4d2b28ye5 ;
  wire o2qkf90r783 ;
  wire rn1o3sl83;
  wire z1l80uwh6vyyg34;
  wire zz5wo47gw146x4;
  wire fgr486jx5kevbua;
  wire pvfk1_6o89lmby;
  wire xx87vzbpchg;

  wire rst_aon;

  wire clic_int_mode;
  wire w00ret5k22yud = (~clic_int_mode) & c4boo209; 
  wire ff_heo9iuk1_06 = (~clic_int_mode) & yukl2; 
  wire nws29bnqq53 = (~clic_int_mode) & zmxoq9ga;
  wire le41_affnsq6 = (~clic_int_mode) & mtip;

  k6pp01__lz7owqwu u_ux607_irq_sync (
    .dk2xhkj77a  (core_clk_aon  ),
    .zh6e0v0mmz (core_clk),
    .ru_wi    (rst_aon    ),   
    .avs1_7j   (rx_evt   ),
    .wxmxi1zq5  (nmi  ),

    .g0sg4nb6l3f  (w00ret5k22yud),
    .aey60u5dsgv  (ff_heo9iuk1_06),
    .gf9zfb8tq9sv  (nws29bnqq53),
    .iqg2bp31t  (le41_affnsq6),

    .z1l80uwh6vyyg34(z1l80uwh6vyyg34),
    .rn1o3sl83(rn1o3sl83), 
    .zz5wo47gw146x4(zz5wo47gw146x4),
    .fgr486jx5kevbua(fgr486jx5kevbua),
    .pvfk1_6o89lmby(pvfk1_6o89lmby),
    .xx87vzbpchg(xx87vzbpchg),

    .uc5qxb4d2b28ye5 (uc5qxb4d2b28ye5 ),
    .o2qkf90r783 (o2qkf90r783 ) 
  );










  wire kxmsn0p4ualeps = 1'b0;
  wire ujj9wb8hyzso = 1'b0;





  wire j_r1zrxno8j;
  wire kjc1hiyz;


  wire rb077g2alw88;
  wire o5q5hev;
  wire c8fchlpwl;
  wire fid1178x5nxb;
  wire klwwlfrft;
  wire oi60pknul;


  wire h7fseh5_df0hbx;


  wire e5fbibk7anp8xhvl52n0ajx2; 
  assign core_sleep_value = core_wfi_mode & e5fbibk7anp8xhvl52n0ajx2; 

































































  wire h8xul8_er09on;
  wire emc_bywzarijbo;
  wire umnrzb6pv8dzc;
  wire nv5a7f_68p9ebw;
  wire bebngvg8sove;


  assign j_r1zrxno8j = c8fchlpwl;
  assign kjc1hiyz = rb077g2alw88;


  wire ip80u6bjne;
  wire qz0hhqemjh;
  wire imsbh3sgxkg4;
  wire vlb2az38tbnj4;

  wire u_ll4hq1b12s2i1;
  wire w41ourymsjpvm8q1e;



  u9lwna1kfmt_pjd_ u_ux607_rst_ctrl (
    .w41ourymsjpvm8q1e(w41ourymsjpvm8q1e),
    .dk2xhkj77a    (core_clk_aon  ),
    .kdnujwd70g0p(por_reset_n    ),
    .k9yxnxeuf0w1(core_reset_n    ),
    .yez0ldac23i95  (reset_bypass),

    .rb077g2alw88   (rb077g2alw88),






    .frilyw4z   (rst_aon) 
  );



   
  wire de1sbr3kjbswue;
  wire nm83rtc_qty;
assign sysrstreq = 1'b0
                 | de1sbr3kjbswue
                 | nm83rtc_qty
                 ;

  wire j4xe_w_yjq2;
  wire j2t29hqv0s6c7;
  wire aui65oshqn8b5_iz6;
  wire jmoafuo8zb_i1t;
  wire sa5of37yr6xn0s3e;
  wire o_dsdljul;
  wire juyzxopct4k03sl;
  wire qyqw_37_fxv8z;
  wire hyw0m71z3q3rpt1;
  wire fx_h7chccf02z;
  wire e592323mqvany;
  wire erv7j3wmd3gb_dp;
  wire wz_if_2q_23jhl2;
  wire n1wslu68m9v;

  wire dyl5g2vgrvy4mb3;
  wire viuu21jzrv;

  wire trtkzwpsx6l;
  wire h87jx93oz7;

  wire bf61lpqg8z;
  wire dnl01g_;



  wire b7ch4h6nrw1vm0;
  wire rcernpf1zf4   ;


  wire y12wg4mlovhn13;
  wire ais_l7yddpa00   ;

  wire b13zu8ysd3u;
  wire itcmps0ezqld   ;

  svx57a7v0ddpyua9ju u_ux607_clk_ctrl(
    .dk2xhkj77a      (core_clk_aon      ),
    .gf33atgy          (core_clk          ),
    .ru_wi        (rst_aon      ),
    .gc4b3kdcan6do88ta_(clkgate_bypass    ),

    .kxmsn0p4ualeps  (kxmsn0p4ualeps),

    .b7ch4h6nrw1vm0   (b7ch4h6nrw1vm0),
    .rcernpf1zf4      (rcernpf1zf4   ),

    .y12wg4mlovhn13   (y12wg4mlovhn13),
    .ais_l7yddpa00      (ais_l7yddpa00   ),

    .b13zu8ysd3u   (b13zu8ysd3u),
    .itcmps0ezqld      (itcmps0ezqld   ),


    .e592323mqvany (e592323mqvany),
    .erv7j3wmd3gb_dp    (erv7j3wmd3gb_dp   ),
    .j4xe_w_yjq2    (j4xe_w_yjq2),
    .j2t29hqv0s6c7 (j2t29hqv0s6c7),
    .aui65oshqn8b5_iz6(aui65oshqn8b5_iz6),
    .jmoafuo8zb_i1t(jmoafuo8zb_i1t),
    .sa5of37yr6xn0s3e(sa5of37yr6xn0s3e),
    .o_dsdljul       (o_dsdljul   ),
    .juyzxopct4k03sl   (juyzxopct4k03sl),
    .qyqw_37_fxv8z   (qyqw_37_fxv8z),
    .hyw0m71z3q3rpt1   (hyw0m71z3q3rpt1),
    .fx_h7chccf02z    (fx_h7chccf02z),

    .wz_if_2q_23jhl2 (wz_if_2q_23jhl2),
    .n1wslu68m9v    (n1wslu68m9v   ),
    .jxdeeywnwq          (),

    .dyl5g2vgrvy4mb3 (dyl5g2vgrvy4mb3),
    .viuu21jzrv    (viuu21jzrv   ),

    .trtkzwpsx6l   (trtkzwpsx6l),
    .h87jx93oz7      (h87jx93oz7   ),

    .bf61lpqg8z   (bf61lpqg8z),
    .dnl01g_      (dnl01g_   ),

    .o5q5hev (o5q5hev      ),
    .c8fchlpwl (c8fchlpwl      ),
    .fid1178x5nxb (fid1178x5nxb      ),
    .ip80u6bjne     (ip80u6bjne     ),
    .qz0hhqemjh  (qz0hhqemjh),
    .ub65ja5c      (),
    .imsbh3sgxkg4     (imsbh3sgxkg4     ),
    .vlb2az38tbnj4  (vlb2az38tbnj4),
    .s_lnrw      (),

    .h8xul8_er09on(h8xul8_er09on),
    .emc_bywzarijbo(emc_bywzarijbo),
    .umnrzb6pv8dzc(umnrzb6pv8dzc),

    .bebngvg8sove  (bebngvg8sove),
    .oi60pknul     (oi60pknul), 

    .nv5a7f_68p9ebw   (nv5a7f_68p9ebw),
    .klwwlfrft      (klwwlfrft   ) 
  );




    
  wire j0qaxhuqtdi;
  wire pbzpk52jinfscit4mm;
  wire gwj6ow6qvbhs0tc31;
  wire [12-1:0] mm0ssgy582fv_j;
  wire iwdkm52x_w4hpak_a2_w;
  wire [64-1:0] ir2913p9xpmq_1bvfd1;
  wire [64-1:0] bsjo0v5e0t556pph;
  wire mwegg_7inaca6povsw;
  wire wnkp7091zrsevkbl;

  wire  [64-1:0] qeb3z0x5;
  wire  ibhfuwrztbm8p4gg;
  wire  [3-1:0] i8_5wt0vppx;
  wire  osv2437qj_3nuf;
  wire b7g_vsn0zoewh6g1;
  wire [2-1:0] onnv64ydiajl;
  wire [2-1:0] r21i4by0bu3ks;
  wire [64-1:0] hn85hkp2yav;


  wire rn2mt6nngsc9w5cz;
  wire c5ewdqztjw9za;
  wire t5trf35s8vy;
  wire zbac123pv78sbz3;
  wire z4e_m564fxae0kpbjr;
  wire zmwq3e9oijvo7d7;

  wire hixy2y36a1pn0;
  wire ozwene1gdpatk6g;
  wire sxvvsxtbhyvt;

  wire [64*4-1:0] azll7rq5fab5ou;
  wire [64*4-1:0] n6a0r_0zddzrme8;
  wire ns0i7siujgkrghjpqv6;




  wire um8zsjyxn_4p; 





  
  
  
  
      
  wire              wex3zbl1x6s4be1en;
  wire [1:0]        pszbl2iobld50k;   
  wire              vfuu2l_7oof31qn0_a;   
  wire [32    -1:0] bvy9o58rgxtbjz_xph;    
  wire [2:0]        gcpthp2sfxb3cxo;
  wire [2:0]        xzjdk5deciqs4l3my_l;
  wire [3:0]        peug05ptx4vv93u4xc; 
  wire [64    -1:0] dlg9f36umgj9xdv0wa;   
  wire  [64    -1:0] yienty7ycnc25au;   
  wire  [1:0]        rxlx2eq69oye0ba3;    
  wire               j2amhrzbhku8dzd;  

  wire resethaltreq;

  
  
  
  wire                       fkm9up63o1aeauaqhjb;
  wire                       to_1lv9wnb3vmu6tvz5rc;
  wire [32-1:0] ju1kbeplcqy314lfj4; 
  wire                       r985fbe5k7hgzaq9i; 
  wire                       bb04gpwotp2s6c7_p1gqkq; 
  wire                       sqmey185cu3mtixhl; 
  wire                       rffcsd1o699ytclmx;
  wire  [64-1:0]     lbr88vbqtg8rht7320frde;
  wire  [8-1:0]  g7qq38mx3d58n1b15kcia;
  wire                       demg_fwfkmaeawq30t;
  wire                       grtb6ypa0px2gi1c;
  wire  [1:0]                f128d8ws0seoihu1;
  wire                       m2r7mfmq3afdd1ine;
  wire                       nhafiywg3hg_52kogwh;
  wire                       xrqayy6vigrw66z8a  ;
  wire                       jyy72ywt9nbo10f2jxupacld;
  wire [64-1:0]      drz92qecqx_qtxwro;
  wire                       st4f16aums5; 
  wire                       p05ld2ghmwh; 


  assign rn2mt6nngsc9w5cz = resethaltreq;

  wire q4gqhurcazjpsf4h;


  wire a02zzbowpjn06h;
  wire jzwasdy8fj0howe;


  pulwy5sk17o3m9m6x u_ux607_dbg_top(

    .idi3vfnshcpo    (core_clk_aon),
    .jzwasdy8fj0howe      (jzwasdy8fj0howe),
    .a02zzbowpjn06h  (a02zzbowpjn06h),
    .um8zsjyxn_4p       (um8zsjyxn_4p),
    .u_ll4hq1b12s2i1    (u_ll4hq1b12s2i1    ),
    .w41ourymsjpvm8q1e(w41ourymsjpvm8q1e),

    .t4bp4v54b9fmhin      (jtag_TDI), 
    .truuny5aeeb6afbba     (), 
    .dc8ehbd4k6bl2re764fz  (), 
    .i3cufk3oe15lxb_x      (1'b0), 
    .q9x26ou3eg17z     (jtag_TDO), 
    .mzb743s60gk6mhj37sy  (jtag_DRV_TDO), 
    .pom74hc61wlcgj8      (jtag_TMS), 
    .pik73_qshqijdw     (), 
    .h9xe65iyw9qxvfp6  (), 
    .ndlpsbtthtn7hv     (1'b0), 
    .v6pe_zs7a1rf5a    (), 
    .dz3fwvx3e10_j6bfrgbzu (), 
    .dlkg75fv         (jtag_TCK), 

    .v66uy2mvzfhls6     (dbg_toggle_a),

    .kdnujwd70g0p     (por_reset_n   ),   
    .yez0ldac23i95    (reset_bypass  ),
    .gc4b3kdcan6do88ta_  (clkgate_bypass),


    .agsknykmgwpc        (nm83rtc_qty   ),
    .u6j3yp5u249c9in70r6h(i_dbg_stop ),
    .pjy0x0i1ftpgz1lr_3dk(override_dm_sleep ),
                    
    .io5ukym11gp2utw    (resethaltreq   ),


    
    .rb050tnl        (j0qaxhuqtdi      ),
    .a94vd35etec4      (pbzpk52jinfscit4mm    ),
    .el7_p8jit09      (gwj6ow6qvbhs0tc31    ),
    .izhvh9xxvwe2   (iwdkm52x_w4hpak_a2_w ),
    .e1go3iu        (mm0ssgy582fv_j      ),
    .l9erxxpnphqd26vg9   (bsjo0v5e0t556pph ),
    .vf5xcr67bqhzlo43_   (ir2913p9xpmq_1bvfd1 ),
    .u2dvoyt5e7o_03z9z5 (mwegg_7inaca6povsw),
    .s904ol6a25v9zn8   (wnkp7091zrsevkbl),

      .qeb3z0x5         (qeb3z0x5        ),
      .ibhfuwrztbm8p4gg     (ibhfuwrztbm8p4gg    ),
      .i8_5wt0vppx      (i8_5wt0vppx     ),
      .osv2437qj_3nuf  (osv2437qj_3nuf ),


      .b7g_vsn0zoewh6g1    (b7g_vsn0zoewh6g1),
      .onnv64ydiajl        (onnv64ydiajl    ),
      .r21i4by0bu3ks       (r21i4by0bu3ks   ),
    .hn85hkp2yav       (hn85hkp2yav),
                             
    .azll7rq5fab5ou      (azll7rq5fab5ou      ),
    .n6a0r_0zddzrme8      (n6a0r_0zddzrme8      ),
    .ns0i7siujgkrghjpqv6(ns0i7siujgkrghjpqv6),

    .pydatzxqqi        (hart_halted),
    .t5trf35s8vy      (t5trf35s8vy),
    .zbac123pv78sbz3   (zbac123pv78sbz3),
    .z4e_m564fxae0kpbjr   (z4e_m564fxae0kpbjr),
    .zmwq3e9oijvo7d7   (zmwq3e9oijvo7d7),
    .q4gqhurcazjpsf4h    (q4gqhurcazjpsf4h),

    .c5ewdqztjw9za        (c5ewdqztjw9za),

    .hixy2y36a1pn0   (hixy2y36a1pn0),
    .ozwene1gdpatk6g      (ozwene1gdpatk6g   ),
    .sxvvsxtbhyvt      (sxvvsxtbhyvt   ),
    .rn1o3sl83       (rn1o3sl83    ),

	.wex3zbl1x6s4be1en    (wex3zbl1x6s4be1en    ),
	.pszbl2iobld50k    (pszbl2iobld50k    ),
	.vfuu2l_7oof31qn0_a    (vfuu2l_7oof31qn0_a    ),
	.bvy9o58rgxtbjz_xph     (bvy9o58rgxtbjz_xph     ),
	.gcpthp2sfxb3cxo     (gcpthp2sfxb3cxo     ),
	.xzjdk5deciqs4l3my_l    (xzjdk5deciqs4l3my_l    ),
	.dlg9f36umgj9xdv0wa    (dlg9f36umgj9xdv0wa    ),
	.peug05ptx4vv93u4xc     (peug05ptx4vv93u4xc     ),
	.yienty7ycnc25au    (yienty7ycnc25au    ),
	.j2amhrzbhku8dzd    (j2amhrzbhku8dzd    ),
	.rxlx2eq69oye0ba3     (rxlx2eq69oye0ba3     ),
	.fkm9up63o1aeauaqhjb (fkm9up63o1aeauaqhjb ),
	.to_1lv9wnb3vmu6tvz5rc (to_1lv9wnb3vmu6tvz5rc ),
	.ju1kbeplcqy314lfj4  (ju1kbeplcqy314lfj4  ), 
	.r985fbe5k7hgzaq9i  (r985fbe5k7hgzaq9i  ), 
	.bb04gpwotp2s6c7_p1gqkq (bb04gpwotp2s6c7_p1gqkq ), 
	.sqmey185cu3mtixhl (sqmey185cu3mtixhl ), 
	.rffcsd1o699ytclmx (rffcsd1o699ytclmx ),
	.lbr88vbqtg8rht7320frde (lbr88vbqtg8rht7320frde ),
	.g7qq38mx3d58n1b15kcia (g7qq38mx3d58n1b15kcia ),
	.demg_fwfkmaeawq30t  (demg_fwfkmaeawq30t  ),
	.grtb6ypa0px2gi1c  (grtb6ypa0px2gi1c  ),
	.f128d8ws0seoihu1  (f128d8ws0seoihu1  ),
	.m2r7mfmq3afdd1ine (m2r7mfmq3afdd1ine ),
	.nhafiywg3hg_52kogwh (nhafiywg3hg_52kogwh ),
	.xrqayy6vigrw66z8a   (xrqayy6vigrw66z8a   ),
	.jyy72ywt9nbo10f2jxupacld(jyy72ywt9nbo10f2jxupacld),
	.drz92qecqx_qtxwro (drz92qecqx_qtxwro ),
	.st4f16aums5         (st4f16aums5         ), 
	.p05ld2ghmwh         (p05ld2ghmwh         ), 

    .rb077g2alw88       (rb077g2alw88),

    .j_r1zrxno8j        (j_r1zrxno8j),
    .kjc1hiyz        (kjc1hiyz) 
  );













  wire                         l9z66pxhit_o_1iyjp;
  wire                         jdh22q4xq9e7wiznv;
  wire [32-1:0]   y_z_yc9_f4ppblmsch3z5; 
  wire                         nmp2x4e8pl59l6he_f9_; 
  wire                         yc7tq3wh6q569ueq7i07em; 
  wire                         yfy18a1ju6mptqd0_u; 
  wire                         gducqncehu9g7n4lydij_0; 
  wire [32-1:0]        dd_gpw58ph81_864rnspr;
  wire [4-1:0]      nhzg88_kzsk0fbtrtku;

  wire                         ixpwz6oo67i61vepd74;
  wire                         t7hb1k3tkjzooetwf;
  wire                         da2pgeraioxt6edc  ;
  wire [32-1:0]        u2fwd1l2_bdiuiftn;

  wire                         ooqxby68qkbvkc5xteznb_x;
  wire                         zhr6liff5rm5wfulyyq;
  wire [32-1:0]   xlsvmbo_v42zk9mypgihxz; 
  wire                         pzv82u11m6kxelyx220ilq5; 
  wire                         yhhbbaf9pqjys_bjgq6h4gj; 
  wire                         qbaqr2mf9nkictp7plgs; 
  wire                         ijehxhtls_byykogg4h; 
  wire [32-1:0]        ylsn7ect00nktb3n8gy6;
  wire [4-1:0]      etkmv0abc25lclz_o85;

  wire                         txrvwlqb8aeb5k6eo4p0tb2;
  wire                         q8mbpl9ben1u54xn_d;
  wire                         igk23ds0cu4_sziqf  ;
  wire [32-1:0]        rsvzuajc8qp4__n0807;
  wire                          dz0zrf512290tvcy4q;
  wire                          core_in_int;
  wire                          mnxti_valid_taken;

  wire                          mip_pmovi;
  wire                          mip_imecci;

  wire                          clic_irq_r;
  wire [9:0]                    clic_irq_id;
  wire                          clic_irq_shv;
  wire [7:0]                    mintstatus_mil_r;
  wire [7:0]                    clic_irq_lvl; 
  wire                          znzjygllppv1s0a8cqub3c;
  wire                          aw82i964do;
  wire                          y8_gkxsfle;
  wire                          fzdb65fcrotwcaccus_cwo;
  wire [7:0]                    tcy_87vt9vet39knuw;
  wire                          fc_4ns_w1nh4h02z_dgg;
  wire                          jqsukc5b5drcc1e78;
  wire                          gnn46rd7vvofruqij;

  wire                         sc9dq6vpj_vb3unfw0;
  wire                         ni7lsi0fuchbbgfizw0l;
  wire [32-1:0]   cvmgqobwfiy_kwo814x; 
  wire                         h_htd26ozpf1rjy0gsvy; 
  wire                         gbzyzsndu75k8rua21_v9c; 
  wire                         w2e5ixihsvl50pgq6b4; 
  wire [32-1:0]        tl_6em2dyajt9yrv4j794c;
  wire [4-1:0]     mf1rr9vurug23q2qsrv;

  wire                         m1vcvvn1ntgzmmwe1bse;
  wire                         f20ikomgiyzoonhphcz;
  wire                         q7emifz3jwxt_jv0_w  ;
  wire [32-1:0]        l1hbm4iglo7pz0pdg_ayjs;



  wire                         bm7mey1b6dibd5i6lfpukeue;

  wire                          a8h5u6ohzhowdrvqrnlllzd70h;
  wire                          pz92yc3xo60c49ayrztvq18a;
  wire  [16-1:0]   pwzrcrecvxehn8htjdn3kv2d0; 
  wire                         ksa323b46ngmxwazg70t76;
  wire                         bs4xe3ath5_4_iwylkfwppp;
  wire                         njyud2m27xz7r6j0g0ieq17m;
  wire                          m5itqssum7ljklhpn5nvzvd93; 
  wire  [64-1:0]        kkk0rwd1njowzq01nvxke;
  wire  [8-1:0]      a2kttuidwhopy02uoajaf;
  wire                          g4hx0dbyp7f7ou8x02a0;
  wire                          zce_icdtm3r9hzeanwhlu3fv;
  wire  [1:0]                   jkp1oke9n1q9ikytwx_7k;

  wire                          mu3ut_ezr05qz2bbi7_vc_aod;
  wire                          sk3bm3yc69h4ac84pc4killh;
  wire                          b7g_hkjxumf964flze01v6p  ;
  wire                          cmtnwdaxz9zk1858kalga2vt  ;
  wire  [64-1:0]        qjvmrd1013dapqkahq_f87b;

  wire                          x0i6aykuzxn1t7_hyw9s7r4to;
  wire                          pbyudse8quydhisrzo9pbl4;
  wire [16-1:0]    vapgj050raiah87lnzt_a; 
  wire                          cvksl3f95u8b10a3rmr6qvom;
  wire                          togorwkvhfveb6zwndvww;
  wire                          i036i6j05gm5ht39aak7k;
  wire                          xubhke6y45gk7d9bj7c1022icq;
  wire                          nao0kbyh1yex0kg7uycyc;

  wire                          c8u60qjfyfel53grl6lmf5_3; 
  wire                          vhl77l_vrkmhgbq9nx8p8ix;   
  wire [64-1:0]         sedkfhar7baq5_wmvydzjmit2; 
  wire                          sf4u33sbbh0akueinpc6j4ly8ue; 



  wire                          ndsqg7zrec89ncrv9yu3k;
  wire                          eth8quxx9hhjhxr4u9k2s77f;
  wire                          zw6mbnvv_8hcztypnytp87v_vy;
  wire  [16-1:0]   l_s_khzs83700pzjuq3_obo44; 
  wire                          kyvscpwy0vljnwysfxqxb;
  wire                          sl5cpfvi658e8pl6nh2cm4;
  wire                          tmqgi_fx924f3bq8ms4u8t0;
  wire                          tcrjx_8vlmtrlqjvk3tu; 
  wire  [64-1:0]      y0jaju01t8mqh2ycz05limpxfu;
  wire  [8-1:0]      x88dy7qz1z117o2jmbslutlpm;
  wire                          kykdx6vx9n3hm7k6oybv;
  wire                          b59iokn7e2645ocyqifdk6sp1;
  wire  [1:0]                   xs2l1_f3yynnrl_rw2zbe;

  wire                          hf8rqlrzsk0e9ho4orde_r;
  wire                          opns8_xijy8grr0gygeszh;
  wire                          hng3_y3ldjtyu4a9n45  ;
  wire                          y1ovf4ea_l0kgs84_pwk6czrs  ;
  wire  [64-1:0]        n6fa00b9i708mtqu7yc9wjvxip;


  wire  [31:0]                  nwk1l6uz4;
  wire  [31:0]                  ir_9aedxd8;

  wire [8*32-1:0] pcr4upio7_tx37; 
  wire [8*1-1:0] uzklqlncpqqm1rav;
  wire [8*1-1:0] ortueunvnkx_l5m_j;
  wire [8*1-1:0] hwuhtb7ucto_utk56;
  wire [8*2-1:0] i1env2kmns7qvvuuc;
  wire [8*1-1:0] g3s3vpafvy3i;

  wire [6-1:0] z6tf8fwcfv0tw03; 

  assign mmu_tlb_way0_addr = z6tf8fwcfv0tw03; 
  assign mmu_tlb_way1_addr = z6tf8fwcfv0tw03; 

  hdkje04yactero u_ux607_ucore(

    .sfyn3seo6gs      (exu_i_valid),
    .sgthjbo1oq1kw1e6      (exu_i_ready),
    .ollg7               (x3),
    .d3n7pwgwcgze9cr4  (alu_cmt_i_valid),
    .amc4c8vcbecv1i     (alu_cmt_i_pc   ),  
    .pby60vfdze02     (mscratch_ena),
    .vm3pyzc9nt95     (mscratch_nxt),
    .rbz4pv_atxqopdwt     (sscratch_ena),
    .qs1xgat7r8xow     (sscratch_nxt),

    .av1w8ld09cfofn     (trace_ivalid    ),
    .im2b5l0h98avl6t4sj (trace_iexception),
    .bw65wl7fvekfymd8vqx  (trace_interrupt ),
    .pecbpcoa04vq      (trace_cause     ),
    .tb_snaxyfs       (trace_tval      ),
    .zc4mldgm25r      (trace_iaddr     ),
    .d23wb5yh1iyvf      (trace_instr     ),
    .srim3bfnzhve       (trace_priv      ),
    .cy3nuhzm_v2p73mt  (trace_bjp_taken ), 
    .fvqwdz2hdbb      (trace_dmode     ),


    .w41ourymsjpvm8q1e(w41ourymsjpvm8q1e),
    .u_ll4hq1b12s2i1    (u_ll4hq1b12s2i1    ),
    .io5ukym11gp2utw    (resethaltreq   ),
     .a02zzbowpjn06h (a02zzbowpjn06h),


      .wd9dvepxj        (reset_vector),

      .tw5xnp59d8x        (core_wfi_mode),
      .um8zsjyxn_4p       (um8zsjyxn_4p),







      .h7fseh5_df0hbx    (h7fseh5_df0hbx),

      .i_x3a8jgmo8qd81tcr    (1'b0),


      .uc5qxb4d2b28ye5          (uc5qxb4d2b28ye5),
      .o2qkf90r783          (o2qkf90r783),

      .habgbg2jn3qi       (e5fbibk7anp8xhvl52n0ajx2),
      .dg4hzu_          (tx_evt     ),












      .j0qaxhuqtdi        (j0qaxhuqtdi      ),
      .pbzpk52jinfscit4mm      (pbzpk52jinfscit4mm    ),
      .gwj6ow6qvbhs0tc31      (gwj6ow6qvbhs0tc31    ),
      .iwdkm52x_w4hpak_a2_w   (iwdkm52x_w4hpak_a2_w ),
      .mm0ssgy582fv_j        (mm0ssgy582fv_j      ),
      .bsjo0v5e0t556pph   (bsjo0v5e0t556pph ),
      .ir2913p9xpmq_1bvfd1   (ir2913p9xpmq_1bvfd1 ),
      .mwegg_7inaca6povsw (mwegg_7inaca6povsw),
      .wnkp7091zrsevkbl   (wnkp7091zrsevkbl),


    
    
      .qeb3z0x5         (qeb3z0x5        ),
      .ibhfuwrztbm8p4gg     (ibhfuwrztbm8p4gg    ),
      .i8_5wt0vppx      (i8_5wt0vppx     ),
      .osv2437qj_3nuf  (osv2437qj_3nuf ),


      .b7g_vsn0zoewh6g1    (b7g_vsn0zoewh6g1),
      .onnv64ydiajl        (onnv64ydiajl    ),
      .r21i4by0bu3ks       (r21i4by0bu3ks   ),
      .hn85hkp2yav       (hn85hkp2yav),

      .azll7rq5fab5ou      (azll7rq5fab5ou      ),
      .n6a0r_0zddzrme8      (n6a0r_0zddzrme8      ),
      .ns0i7siujgkrghjpqv6(ns0i7siujgkrghjpqv6),

      .pydatzxqqi        (hart_halted),
      .t5trf35s8vy      (t5trf35s8vy),
      .zbac123pv78sbz3   (zbac123pv78sbz3),
      .z4e_m564fxae0kpbjr   (z4e_m564fxae0kpbjr),
      .zmwq3e9oijvo7d7   (zmwq3e9oijvo7d7),

      .c5ewdqztjw9za        (c5ewdqztjw9za  ),
      .rn2mt6nngsc9w5cz(rn2mt6nngsc9w5cz),

      .hixy2y36a1pn0   (hixy2y36a1pn0),
      .ozwene1gdpatk6g      (ozwene1gdpatk6g   ),
      .sxvvsxtbhyvt      (sxvvsxtbhyvt   ),

    

      .pcr4upio7_tx37     (pcr4upio7_tx37   ), 
      .uzklqlncpqqm1rav  (uzklqlncpqqm1rav),
      .ortueunvnkx_l5m_j  (ortueunvnkx_l5m_j),
      .hwuhtb7ucto_utk56  (hwuhtb7ucto_utk56),
      .i1env2kmns7qvvuuc  (i1env2kmns7qvvuuc),
      .g3s3vpafvy3i  (g3s3vpafvy3i),



      .v09gw6e6rfjf05qg    (hart_id),  




      .fcjh1nct4r             (clic_irq_r),
      .f_i1959b4xizzq9jea     (mintstatus_mil_r),
      .b4lwcgm6l21pi          (clic_irq_id),
      .hjrk_rwjkqj3zk_b         (clic_irq_lvl),
      .zwcbp7zqfei5xz         (clic_irq_shv),
      .znzjygllppv1s0a8cqub3c    (znzjygllppv1s0a8cqub3c), 
      .dxi_ue3gf5zqqqxwgq2a    (mnxti_valid_taken),
      .ix299qulxi5            (mip_pmovi    ),
      .jjj61w03m77lv           (mip_imecci    ),
      .gfy3zost37aq8qmr          (core_in_int),
      .dz0zrf512290tvcy4q        (dz0zrf512290tvcy4q),
      .dn8riluj40uunvq5        (clic_int_mode),
      .aw82i964do               (aw82i964do            ),
      .y8_gkxsfle               (y8_gkxsfle            ),
      .fzdb65fcrotwcaccus_cwo    (fzdb65fcrotwcaccus_cwo ),
      .tcy_87vt9vet39knuw     (tcy_87vt9vet39knuw  ),
      .fc_4ns_w1nh4h02z_dgg   (fc_4ns_w1nh4h02z_dgg),
      .jqsukc5b5drcc1e78       (jqsukc5b5drcc1e78    ),
      .gnn46rd7vvofruqij       (gnn46rd7vvofruqij    ),
      .x_cq40qmp6a          (x_cq40qmp6a       ),




      .z1l80uwh6vyyg34 (z1l80uwh6vyyg34),
      .rn1o3sl83     (rn1o3sl83),
      .zz5wo47gw146x4    (zz5wo47gw146x4),
      .fgr486jx5kevbua    (fgr486jx5kevbua),
      .pvfk1_6o89lmby     (pvfk1_6o89lmby),
      .xx87vzbpchg     (xx87vzbpchg),






    .ij_sgq3rtvw2          (nwk1l6uz4),
    .k9jntnqwqp         (ir_9aedxd8),


    .nv5a7f_68p9ebw   (nv5a7f_68p9ebw),
    .klwwlfrft      (klwwlfrft      ),

    .bebngvg8sove  (bebngvg8sove),
    .oi60pknul     (oi60pknul), 



    .bm7mey1b6dibd5i6lfpukeue      (bm7mey1b6dibd5i6lfpukeue    ),

    .a8h5u6ohzhowdrvqrnlllzd70h    (a8h5u6ohzhowdrvqrnlllzd70h  ),
    .pz92yc3xo60c49ayrztvq18a    (pz92yc3xo60c49ayrztvq18a  ),
    .pwzrcrecvxehn8htjdn3kv2d0     (pwzrcrecvxehn8htjdn3kv2d0   ),
    .ksa323b46ngmxwazg70t76    (ksa323b46ngmxwazg70t76  ),
    .bs4xe3ath5_4_iwylkfwppp    (bs4xe3ath5_4_iwylkfwppp  ),
    .njyud2m27xz7r6j0g0ieq17m    (njyud2m27xz7r6j0g0ieq17m  ),
    .m5itqssum7ljklhpn5nvzvd93     (m5itqssum7ljklhpn5nvzvd93   ),
    .kkk0rwd1njowzq01nvxke    (kkk0rwd1njowzq01nvxke  ),
    .a2kttuidwhopy02uoajaf    (a2kttuidwhopy02uoajaf  ),
    .g4hx0dbyp7f7ou8x02a0     (g4hx0dbyp7f7ou8x02a0   ),
    .zce_icdtm3r9hzeanwhlu3fv     (zce_icdtm3r9hzeanwhlu3fv   ),
    .jkp1oke9n1q9ikytwx_7k     (jkp1oke9n1q9ikytwx_7k   ),
                                                       
    .mu3ut_ezr05qz2bbi7_vc_aod    (mu3ut_ezr05qz2bbi7_vc_aod  ),
    .sk3bm3yc69h4ac84pc4killh    (sk3bm3yc69h4ac84pc4killh  ),
    .b7g_hkjxumf964flze01v6p      (b7g_hkjxumf964flze01v6p    ),
    .cmtnwdaxz9zk1858kalga2vt  (cmtnwdaxz9zk1858kalga2vt), 
    .qjvmrd1013dapqkahq_f87b    (qjvmrd1013dapqkahq_f87b  ),
                                                      
    .x0i6aykuzxn1t7_hyw9s7r4to    (x0i6aykuzxn1t7_hyw9s7r4to  ),
    .pbyudse8quydhisrzo9pbl4    (pbyudse8quydhisrzo9pbl4  ),
    .vapgj050raiah87lnzt_a     (vapgj050raiah87lnzt_a   ),
    .cvksl3f95u8b10a3rmr6qvom    (cvksl3f95u8b10a3rmr6qvom   ),
    .togorwkvhfveb6zwndvww    (togorwkvhfveb6zwndvww   ),
    .i036i6j05gm5ht39aak7k    (i036i6j05gm5ht39aak7k   ),
    .xubhke6y45gk7d9bj7c1022icq    (xubhke6y45gk7d9bj7c1022icq   ),
	.nao0kbyh1yex0kg7uycyc      (nao0kbyh1yex0kg7uycyc     ),
                                                     
    .c8u60qjfyfel53grl6lmf5_3    (c8u60qjfyfel53grl6lmf5_3  ),
    .vhl77l_vrkmhgbq9nx8p8ix      (vhl77l_vrkmhgbq9nx8p8ix    ),
    .sedkfhar7baq5_wmvydzjmit2    (sedkfhar7baq5_wmvydzjmit2  ),
    .sf4u33sbbh0akueinpc6j4ly8ue   (sf4u33sbbh0akueinpc6j4ly8ue ), 
                                                    

    .ndsqg7zrec89ncrv9yu3k      (ndsqg7zrec89ncrv9yu3k  ),

    .eth8quxx9hhjhxr4u9k2s77f    (eth8quxx9hhjhxr4u9k2s77f  ),
    .zw6mbnvv_8hcztypnytp87v_vy    (zw6mbnvv_8hcztypnytp87v_vy  ),
    .l_s_khzs83700pzjuq3_obo44     (l_s_khzs83700pzjuq3_obo44   ),
    .kyvscpwy0vljnwysfxqxb    (kyvscpwy0vljnwysfxqxb  ),
    .sl5cpfvi658e8pl6nh2cm4    (sl5cpfvi658e8pl6nh2cm4  ),
    .tmqgi_fx924f3bq8ms4u8t0    (tmqgi_fx924f3bq8ms4u8t0  ),
    .tcrjx_8vlmtrlqjvk3tu     (tcrjx_8vlmtrlqjvk3tu   ),
    .y0jaju01t8mqh2ycz05limpxfu    (y0jaju01t8mqh2ycz05limpxfu  ),
    .x88dy7qz1z117o2jmbslutlpm    (x88dy7qz1z117o2jmbslutlpm  ),
    .kykdx6vx9n3hm7k6oybv     (kykdx6vx9n3hm7k6oybv   ),
    .b59iokn7e2645ocyqifdk6sp1     (b59iokn7e2645ocyqifdk6sp1   ),
    .xs2l1_f3yynnrl_rw2zbe     (xs2l1_f3yynnrl_rw2zbe   ),
  
    .hf8rqlrzsk0e9ho4orde_r    (hf8rqlrzsk0e9ho4orde_r  ),
    .opns8_xijy8grr0gygeszh    (opns8_xijy8grr0gygeszh  ),
    .hng3_y3ldjtyu4a9n45      (hng3_y3ldjtyu4a9n45    ),
    .y1ovf4ea_l0kgs84_pwk6czrs  (y1ovf4ea_l0kgs84_pwk6czrs), 
    .n6fa00b9i708mtqu7yc9wjvxip    (n6fa00b9i708mtqu7yc9wjvxip  ),
    


    .ooqxby68qkbvkc5xteznb_x     (ooqxby68qkbvkc5xteznb_x),
    .zhr6liff5rm5wfulyyq     (zhr6liff5rm5wfulyyq),
    .xlsvmbo_v42zk9mypgihxz      (xlsvmbo_v42zk9mypgihxz ),
    .pzv82u11m6kxelyx220ilq5     (pzv82u11m6kxelyx220ilq5),
    .yhhbbaf9pqjys_bjgq6h4gj     (yhhbbaf9pqjys_bjgq6h4gj),
    .qbaqr2mf9nkictp7plgs     (qbaqr2mf9nkictp7plgs),
    .ijehxhtls_byykogg4h      (ijehxhtls_byykogg4h ),
    .ylsn7ect00nktb3n8gy6     (ylsn7ect00nktb3n8gy6),
    .etkmv0abc25lclz_o85     (etkmv0abc25lclz_o85),
    
    .txrvwlqb8aeb5k6eo4p0tb2     (txrvwlqb8aeb5k6eo4p0tb2),
    .q8mbpl9ben1u54xn_d     (q8mbpl9ben1u54xn_d),
    .igk23ds0cu4_sziqf       (igk23ds0cu4_sziqf  ),
    .rsvzuajc8qp4__n0807     (rsvzuajc8qp4__n0807),
    .sc9dq6vpj_vb3unfw0     (sc9dq6vpj_vb3unfw0),
    .ni7lsi0fuchbbgfizw0l     (ni7lsi0fuchbbgfizw0l),
    .cvmgqobwfiy_kwo814x      (cvmgqobwfiy_kwo814x ),
    .h_htd26ozpf1rjy0gsvy     (h_htd26ozpf1rjy0gsvy),
    .gbzyzsndu75k8rua21_v9c     (gbzyzsndu75k8rua21_v9c),
    .w2e5ixihsvl50pgq6b4      (w2e5ixihsvl50pgq6b4 ),
    .tl_6em2dyajt9yrv4j794c     (tl_6em2dyajt9yrv4j794c),
    .mf1rr9vurug23q2qsrv     (mf1rr9vurug23q2qsrv),
    
    .m1vcvvn1ntgzmmwe1bse     (m1vcvvn1ntgzmmwe1bse),
    .f20ikomgiyzoonhphcz     (f20ikomgiyzoonhphcz),
    .q7emifz3jwxt_jv0_w       (q7emifz3jwxt_jv0_w  ),
    .l1hbm4iglo7pz0pdg_ayjs     (l1hbm4iglo7pz0pdg_ayjs),

    .l9z66pxhit_o_1iyjp     (l9z66pxhit_o_1iyjp),
    .jdh22q4xq9e7wiznv     (jdh22q4xq9e7wiznv),
    .y_z_yc9_f4ppblmsch3z5      (y_z_yc9_f4ppblmsch3z5 ),
    .yc7tq3wh6q569ueq7i07em     (yc7tq3wh6q569ueq7i07em),
    .yfy18a1ju6mptqd0_u     (yfy18a1ju6mptqd0_u),
    .gducqncehu9g7n4lydij_0     (gducqncehu9g7n4lydij_0),
    .nmp2x4e8pl59l6he_f9_      (nmp2x4e8pl59l6he_f9_ ),
    .dd_gpw58ph81_864rnspr     (dd_gpw58ph81_864rnspr),
    .nhzg88_kzsk0fbtrtku     (nhzg88_kzsk0fbtrtku),
    
    .ixpwz6oo67i61vepd74     (ixpwz6oo67i61vepd74),
    .t7hb1k3tkjzooetwf     (t7hb1k3tkjzooetwf),
    .da2pgeraioxt6edc       (da2pgeraioxt6edc  ),
    .u2fwd1l2_bdiuiftn     (u2fwd1l2_bdiuiftn),



     .wh6iy6zpdqsnv2y (mem_arready),
     .bd6yatp5cqq (mem_arvalid),
     .fl1qsvyu    (        ),
     .b9889wezsu  (mem_araddr),
     .an__mxugc4   (mem_arlen),
     .poj6g8vw9e  (mem_arsize),
     .dafaivw3ze9g3hi (mem_arburst),
     .q2c0d6fxz_1bw  (mem_arlock),
     .wblesminvapwua (mem_arcache),
     .v3cim36gj8g  (mem_arprot),
     .ss22f8fuy2uhr   (         ),
     .hoaoalj5pcdnpnm0(            ),
     .rh8f1e3jgg3xi  (          ),
     .roral7fym4h3_ (mem_awready),
     .b_gwvq35iq0_yvk (mem_awvalid),
     .lqm2hm0cjm5zt    (        ),
     .f3n3tpjs44e0_  (mem_awaddr),
     .dmc59hxf352z   (mem_awlen),
     .a63l3og_8qak5jy  (mem_awsize),
     .m0wp58qmji79 (mem_awburst),
     .c8qmnfk1vqai  (mem_awlock),
     .pbov8g9yizcwr (mem_awcache),
     .t8qjehupeajtzjr  (mem_awprot),
     .hhp1rh0x0jn   (         ),
     .w9yptl69xj6p(            ),
     .yvcpy_gyehs4lji  (          ), 
     .kted7ph0krq  (mem_wready),
     .a93i3d2hji  (mem_wvalid),
     .of5p5cb8p4     (          ),
     .g1bi1xzuv64   (mem_wdata),
     .gj6p5b5ik3r9p   (mem_wstrb),
     .m1fmaas4oww6   (mem_wlast),
     .hjstsi51gm  (mem_rready),
     .onpqhy0s69  (mem_rvalid),
     .aw7xjbi     (4'h0),
     .z0cc2y_uzoh_   (mem_rdata),
     .y8tc_vywu82ugn   (mem_rresp),
     .o2h9d51o6m6   (mem_rlast),
     .nneek3ep5xykwl  (mem_bready),
     .g8khua4l0y77zjp  (mem_bvalid),
     .wmlp1a2b     (4'h0),
     .weop50xb_avne   (mem_bresp),
     .su81e8dxdzng9d (mem_clk_en),

 
    .lueem7uei21mn66 (ppi_ahbl_htrans) ,  
    .vgodhub5af4gihqv5eef (ppi_ahbl_hwrite) ,  
    .lueqjwqinfpts52  (ppi_ahbl_haddr ) ,  
    .lv9moee8_5_8dsy5  (ppi_ahbl_hsize ) ,  
    .ck0wbvgghs6n9j4 (ppi_ahbl_hwdata) ,  
    .uecfgtalcganlj42vmq  (ppi_ahbl_hprot ) ,
    .msxgfr_x73l96858p1s (ppi_ahbl_hrdata) ,  
    .tze074ath5y6h2m41  (ppi_ahbl_hresp ) ,  
    .o752t3g6xbcxc6if88wi (ppi_ahbl_hready) , 

    .nprvxoyk8ecm174bi8 (ppi_ahbl_clk_en) , 





	.wex3zbl1x6s4be1en    (wex3zbl1x6s4be1en    ),
	.pszbl2iobld50k    (pszbl2iobld50k    ),
	.vfuu2l_7oof31qn0_a    (vfuu2l_7oof31qn0_a    ),
	.bvy9o58rgxtbjz_xph     (bvy9o58rgxtbjz_xph     ),
	.gcpthp2sfxb3cxo     (gcpthp2sfxb3cxo     ),
	.xzjdk5deciqs4l3my_l    (xzjdk5deciqs4l3my_l    ),
	.dlg9f36umgj9xdv0wa    (dlg9f36umgj9xdv0wa    ),
	.peug05ptx4vv93u4xc     (peug05ptx4vv93u4xc     ),
	.yienty7ycnc25au    (yienty7ycnc25au    ),
	.j2amhrzbhku8dzd    (j2amhrzbhku8dzd    ),
	.rxlx2eq69oye0ba3     (rxlx2eq69oye0ba3     ),

	.fkm9up63o1aeauaqhjb (fkm9up63o1aeauaqhjb ),
	.to_1lv9wnb3vmu6tvz5rc (to_1lv9wnb3vmu6tvz5rc ),
	.ju1kbeplcqy314lfj4  (ju1kbeplcqy314lfj4  ), 
	.r985fbe5k7hgzaq9i  (r985fbe5k7hgzaq9i  ), 
	.bb04gpwotp2s6c7_p1gqkq (bb04gpwotp2s6c7_p1gqkq ), 
	.sqmey185cu3mtixhl (sqmey185cu3mtixhl ), 
	.rffcsd1o699ytclmx (rffcsd1o699ytclmx ),
	.lbr88vbqtg8rht7320frde (lbr88vbqtg8rht7320frde ),
	.g7qq38mx3d58n1b15kcia (g7qq38mx3d58n1b15kcia ),
	.demg_fwfkmaeawq30t  (demg_fwfkmaeawq30t  ),
	.grtb6ypa0px2gi1c  (grtb6ypa0px2gi1c  ),
	.f128d8ws0seoihu1  (f128d8ws0seoihu1  ),
	.m2r7mfmq3afdd1ine (m2r7mfmq3afdd1ine ),
	.nhafiywg3hg_52kogwh (nhafiywg3hg_52kogwh ),
	.xrqayy6vigrw66z8a   (xrqayy6vigrw66z8a   ),
	.jyy72ywt9nbo10f2jxupacld(jyy72ywt9nbo10f2jxupacld),
	.drz92qecqx_qtxwro (drz92qecqx_qtxwro ),
	.st4f16aums5         (st4f16aums5         ), 
	.p05ld2ghmwh         (p05ld2ghmwh         ), 



    .gc4b3kdcan6do88ta_   (clkgate_bypass), 

    .wz_if_2q_23jhl2  (wz_if_2q_23jhl2),
    .n1wslu68m9v     (n1wslu68m9v   ),

    .svlxg92fk8wh7_jgsa8x (icache_disable_init),

    .v0bybbiepfqv4kc_cdg         (icache_tag0_cs    ),
    .i28_g1tt8nk7e30         (icache_tag0_we    ),
    .m_aqi5ytp0maje5sj       (icache_tag0_addr  ),
    .e2iagwi42o6sun5_ykv9      (icache_tag0_wdata ),        
    .wa_f05baz0i8dkq7t_4y      (icache_tag0_rdata ),
                                                
    .hpf4dbs7lpgqzs89        (icache_data0_cs   ),
    .hlpyb4rsu9gt28ml_u        (icache_data0_we   ),
    .qh651fblp7os_lrh1rf5      (icache_data0_addr ),
    .yalqjjffhlwhb4fi3re     (icache_data0_wdata),        
    .s0j6brb1s7b0asp2o_4vmv0     (icache_data0_rdata),
                                               
    .a9pfw7vdfvtnr1l89         (icache_tag1_cs    ),
    .qmlhx0ddtv5q5m65mb2         (icache_tag1_we    ),
    .gg035mahjzmwm_850rpfm       (icache_tag1_addr  ),
    .faibzt_25z6u6lt9f      (icache_tag1_wdata ),        
    .n_6989smoxxpesripwzs5      (icache_tag1_rdata ),
                                               
    .pq_z6zyr2bjwut728ldr        (icache_data1_cs   ),
    .p4ls8ac9eyqc7uznlkv        (icache_data1_we   ),
    .utq6xdqs0m3irmvrgwe7      (icache_data1_addr ),
    .tw7hzxhmmtptsxpzz1x9d17     (icache_data1_wdata),        
    .tz_zq72t3w19dm7c3a0mu     (icache_data1_rdata),





    .dyl5g2vgrvy4mb3 (dyl5g2vgrvy4mb3),
    .viuu21jzrv    (viuu21jzrv   ),

    .f2qbwkn13kmm9hmrn159wahi (dcache_disable_init),
    
    .mum8f1rtatle7p_55y84     (dcache_w0_tram_cs  ),   
    .pn5bpwlp5ijfako9m5ao   (dcache_w0_tram_addr),
    .g3s0qe2adsxsx8e6z     (dcache_w0_tram_we  ),
    .a1rl4lmhqp8ydyk07kqkn    (dcache_w0_tram_din ),       
    .apnns9jlj7y3y5bg8ynz   (dcache_w0_tram_dout),
                                               
    .pmz7e4mgvbnmimqp0nghk     (dcache_w1_tram_cs  ),
    .j61algpxjoycxbswhgsuf   (dcache_w1_tram_addr),
    .omq1ehm8hp4q9jgp5n5vn     (dcache_w1_tram_we  ),
    .fbv1q6sraswzp91zcn    (dcache_w1_tram_din ),       
    .jv8kv41vzuir6an4iod   (dcache_w1_tram_dout),
                                               
                                               
    .qgl4363n31jx6xjyo05zkn     (dcache_dram_b0_cs  ),
    .zec78nyllxlfwmpsgncluudf   (dcache_dram_b0_addr),
    .dwvnjl0vxqkgd8t6dtvg5z    (dcache_dram_b0_wem ),
    .gngmcj5c1jd85csel9ntru    (dcache_dram_b0_din ),       
    .tkt93y5lfluzkia5plvksp   (dcache_dram_b0_dout),
                                               
    .km7co8hqm563od8ga_03_g     (dcache_dram_b1_cs  ),
    .j4mas6g26o63wvnsdquh8c4p   (dcache_dram_b1_addr),
    .nniah5mh0cunkhyln9    (dcache_dram_b1_wem ),
    .rcy_v3911lf33nza5j    (dcache_dram_b1_din ),       
    .g4nfgu53_rgc0632w8z97   (dcache_dram_b1_dout),
                                               
    .xzgkclcxsgfuseg87     (dcache_dram_b2_cs  ),
    .djwlah5bo0r6myit6cal0t   (dcache_dram_b2_addr),
    .qu_ju3lv6nvkdbo8h11uf    (dcache_dram_b2_wem ),
    .dydwz9i6k80alqfarffop    (dcache_dram_b2_din ),       
    .ql1c7hzoj9kf__7r97krm   (dcache_dram_b2_dout),
                                               
    .kp2j8kv1p1cjcg0lerwm     (dcache_dram_b3_cs  ),
    .v4a7g1wh3ivw0esp7dye0oiz   (dcache_dram_b3_addr),
    .x9zuk21gpaj58uszvm5    (dcache_dram_b3_wem ),
    .n_h5oz0c5bo5rpevwjcu8    (dcache_dram_b3_din ),       
    .ryid4_99ns1jc83at_88x   (dcache_dram_b3_dout),


    .trtkzwpsx6l                      (trtkzwpsx6l                        ),
    .h87jx93oz7                         (h87jx93oz7                           ),
    .moqs2k81l9fugde5v_581            (mmu_tlb_disable_init              ),
    .i0acx70llka5qu09r5jd                 (mmu_tlb_way0_cs                   ), 
    .e44u8ctdv_z5u19to                 (mmu_tlb_way1_cs                   ), 
    .h7k_k0xxi7vktla                 (mmu_tlb_way0_we                   ), 
    .v_vouzmjecsvtjxt                 (mmu_tlb_way1_we                   ), 
    .ef9y8yyld9onuy00de7o              (mmu_tlb_way0_wdata                ), 
    .ammhazyeeglt3ewt4p              (mmu_tlb_way1_wdata                ), 
    .xvwzwg7_3ek2tx                   (z6tf8fwcfv0tw03                      ), 
    .y8sg6kbsyavoh4usiqn               (mmu_tlb_way0_dout                 ), 
    .gnqkycbjc0k9k4_edoube               (mmu_tlb_way1_dout                 ), 


    .bf61lpqg8z  (bf61lpqg8z),
    .dnl01g_     (dnl01g_   ),

    .emc_bywzarijbo    (emc_bywzarijbo),
    .h8xul8_er09on    (h8xul8_er09on),
    .umnrzb6pv8dzc    (umnrzb6pv8dzc),
    .e592323mqvany (e592323mqvany), 
    .o5q5hev       (o5q5hev),
    .c8fchlpwl       (c8fchlpwl),
    .fid1178x5nxb       (fid1178x5nxb),


    .j4xe_w_yjq2     (j4xe_w_yjq2),
    .j2t29hqv0s6c7  (j2t29hqv0s6c7),
    .aui65oshqn8b5_iz6 (aui65oshqn8b5_iz6),
    .jmoafuo8zb_i1t (jmoafuo8zb_i1t),
    .sa5of37yr6xn0s3e (sa5of37yr6xn0s3e),
    .o_dsdljul        (o_dsdljul       ),
    .juyzxopct4k03sl    (juyzxopct4k03sl   ),
    .qyqw_37_fxv8z    (qyqw_37_fxv8z   ),
    .hyw0m71z3q3rpt1    (hyw0m71z3q3rpt1   ),
    .fx_h7chccf02z     (fx_h7chccf02z    ),
    .dk2xhkj77a        (core_clk_aon     ),
    .erv7j3wmd3gb_dp     (erv7j3wmd3gb_dp    ),

    .ru_wi        (rb077g2alw88    )
  );

  ux607_clkgate vrtyktpe3i8f8s7_ioyyl52(
    .clk_in   (core_clk),
    .clkgate_bypass(clkgate_bypass  ),
    .clock_en (icache_tag0_cs),
    .clk_out  (clk_icache_tag0)
  );

  ux607_clkgate bckv8giuqfvu16ft7fqxuml(
    .clk_in   (core_clk),
    .clkgate_bypass(clkgate_bypass  ),
    .clock_en (icache_data0_cs),
    .clk_out  (clk_icache_data0)
  );

  ux607_clkgate bpjz2p0buffvf46tmvn0f2d(
    .clk_in   (core_clk),
    .clkgate_bypass(clkgate_bypass  ),
    .clock_en (icache_tag1_cs),
    .clk_out  (clk_icache_tag1)
  );

  ux607_clkgate wqivggeo35kxu09r6twtw5rag(
    .clk_in   (core_clk),
    .clkgate_bypass(clkgate_bypass  ),
    .clock_en (icache_data1_cs),
    .clk_out  (clk_icache_data1)
  );


  ux607_clkgate eg0454_3y3y79nfyn2vsg9c_pvf(
    .clk_in   (core_clk),
    .clkgate_bypass(clkgate_bypass  ),
    .clock_en (dcache_w0_tram_cs),
    .clk_out  (clk_dcache_w0_tram)
  );

  ux607_clkgate bobvr5ao8ctobfc_vgjsxp_aymz(
    .clk_in   (core_clk),
    .clkgate_bypass(clkgate_bypass  ),
    .clock_en (dcache_w1_tram_cs),
    .clk_out  (clk_dcache_w1_tram)
  );
   
  
  
  ux607_clkgate tjyaxujqlt2nzvshbbaabywofr3(
    .clk_in   (core_clk),
    .clkgate_bypass(clkgate_bypass  ),
    .clock_en (dcache_dram_b0_cs),
    .clk_out  (clk_dcache_dram_b0)
  );

  ux607_clkgate m_3j06xnur7r8096qzrvdtni3z(
    .clk_in   (core_clk),
    .clkgate_bypass(clkgate_bypass  ),
    .clock_en (dcache_dram_b1_cs),
    .clk_out  (clk_dcache_dram_b1)
  );
   
  ux607_clkgate vud8p019crvir4n7juldjb7t(
    .clk_in   (core_clk),
    .clkgate_bypass(clkgate_bypass  ),
    .clock_en (dcache_dram_b2_cs),
    .clk_out  (clk_dcache_dram_b2)
  );
   
   
  ux607_clkgate dbyp7cacnepigvek3gu5lusb275b(
    .clk_in   (core_clk),
    .clkgate_bypass(clkgate_bypass  ),
    .clock_en (dcache_dram_b3_cs),
    .clk_out  (clk_dcache_dram_b3)
  );
   

  ux607_clkgate lkv9q4ni8kd4lq8hc54jmb(
    .clk_in   (core_clk),
    .clkgate_bypass(clkgate_bypass  ),
    .clock_en (mmu_tlb_way0_cs),
    .clk_out  (clk_mmu_tlb_way0)
  );

  ux607_clkgate ee0afbrgf0xodl6qvggbelu(
    .clk_in   (core_clk),
    .clkgate_bypass(clkgate_bypass  ),
    .clock_en (mmu_tlb_way1_cs),
    .clk_out  (clk_mmu_tlb_way1)
  );










  odg9yeykg220ymcco
   #(
      .nm_fj         (16),
      .onr7l         (64),
      .h1b         (8),
      .ktra3i     (3),
      .rm39njpb7w     (13),
      .wvmre88     (64),
      .bf0ngee0t   (1),
      .xbpsp4_i     (8),
      .k2qm7hpa_qinpd (0),
      .quofpn_rylwqbg9 (0) 
      ) r6ak_x8u809k624o_q (
    .qz0hhqemjh          (qz0hhqemjh),
    .ujj9wb8hyzso           (ujj9wb8hyzso),

    .ndsqg7zrec89ncrv9yu3k    (ndsqg7zrec89ncrv9yu3k  ),

    .bm7mey1b6dibd5i6lfpukeue    (bm7mey1b6dibd5i6lfpukeue    ),
                                                    
    .a8h5u6ohzhowdrvqrnlllzd70h  (a8h5u6ohzhowdrvqrnlllzd70h  ),
    .pz92yc3xo60c49ayrztvq18a  (pz92yc3xo60c49ayrztvq18a  ),
    .pwzrcrecvxehn8htjdn3kv2d0   (pwzrcrecvxehn8htjdn3kv2d0   ), 
    .m5itqssum7ljklhpn5nvzvd93   (m5itqssum7ljklhpn5nvzvd93   ), 
    .kkk0rwd1njowzq01nvxke  (kkk0rwd1njowzq01nvxke  ),
    .a2kttuidwhopy02uoajaf  (a2kttuidwhopy02uoajaf  ),
    .g4hx0dbyp7f7ou8x02a0   (g4hx0dbyp7f7ou8x02a0   ),
    .zce_icdtm3r9hzeanwhlu3fv   (zce_icdtm3r9hzeanwhlu3fv   ),
    .jkp1oke9n1q9ikytwx_7k   (jkp1oke9n1q9ikytwx_7k   ),
    .njyud2m27xz7r6j0g0ieq17m  (njyud2m27xz7r6j0g0ieq17m),
    .ksa323b46ngmxwazg70t76  (ksa323b46ngmxwazg70t76),
    .bs4xe3ath5_4_iwylkfwppp  (bs4xe3ath5_4_iwylkfwppp),
    
    .mu3ut_ezr05qz2bbi7_vc_aod  (mu3ut_ezr05qz2bbi7_vc_aod  ),
    .sk3bm3yc69h4ac84pc4killh  (sk3bm3yc69h4ac84pc4killh  ),
    .b7g_hkjxumf964flze01v6p    (b7g_hkjxumf964flze01v6p    ),
    .cmtnwdaxz9zk1858kalga2vt(cmtnwdaxz9zk1858kalga2vt),
    .qjvmrd1013dapqkahq_f87b  (qjvmrd1013dapqkahq_f87b  ),
    

    .c52ldkop361ts52m0    (x0i6aykuzxn1t7_hyw9s7r4to  ),
    .x88wat37r_vjsn57a    (pbyudse8quydhisrzo9pbl4  ),
    .z3k8ps_o7osj4uosf_6i5     (vapgj050raiah87lnzt_a [16-1:0]  ),
    .rzon56p292pybf35mi_    (cvksl3f95u8b10a3rmr6qvom),
    .jn_zyepkhmn_mdbqe1    (togorwkvhfveb6zwndvww),
    .w8k_3fawz__hfg4mk0mw7g    (i036i6j05gm5ht39aak7k),
    .i88maxesdvq1fkint66    (xubhke6y45gk7d9bj7c1022icq),
	.nao0kbyh1yex0kg7uycyc  (nao0kbyh1yex0kg7uycyc  ),
                                                
    .ult8a6a0b4agydwsws    (c8u60qjfyfel53grl6lmf5_3  ),
    .gkbxrtlrxlk7_fk4      (vhl77l_vrkmhgbq9nx8p8ix    ),
    .d27a6w261um4big8wy8    (sedkfhar7baq5_wmvydzjmit2  ),
    .bwdpzndejgg3liwep6q_   (sf4u33sbbh0akueinpc6j4ly8ue ), 
                                                    


    .d53gmmeaj           (ilm_cs   ),  
    .coouz2jyj2n         (ilm_addr ), 
    .dcmn368x8          (ilm_byte_we  ),
    .opsl7g4          (ilm_wdata  ),          
    .tn65z3ytg         (ilm_rdata ),
    .wzor2kya          (             ),

  

      .pcr4upio7_tx37     (pcr4upio7_tx37   ), 
      .uzklqlncpqqm1rav  (uzklqlncpqqm1rav),
      .ortueunvnkx_l5m_j  (ortueunvnkx_l5m_j),
      .hwuhtb7ucto_utk56  (hwuhtb7ucto_utk56),
      .i1env2kmns7qvvuuc  (i1env2kmns7qvvuuc),
      .g3s3vpafvy3i  (g3s3vpafvy3i),

    .gc4b3kdcan6do88ta_       (clkgate_bypass),
    .gf33atgy                  (ip80u6bjne),
    .ru_wi                (rst_aon) 
  );

  ux607_clkgate m7pjy2kppbajsk5ditlri01(
    .clk_in   (core_clk),
    .clkgate_bypass(clkgate_bypass  ),
    .clock_en (ilm_cs),
    .clk_out  (clk_ilm_ram)
  );

  
  
  wire [2-1:0] r6tkd_53z; 
  wire [13-1:0] cyop0l7lnv6j3; 
  wire [8-1:0] g9h1mnhtsaduuk;
  wire [64-1:0] pyxv3lgda85n;      
  wire [64-1:0] k90knfo82df2l;
  assign dlm0_addr = cyop0l7lnv6j3;
  assign dlm1_addr = cyop0l7lnv6j3;
  assign {dlm1_cs,dlm0_cs} = r6tkd_53z;
  assign {dlm1_byte_we, dlm0_byte_we} = g9h1mnhtsaduuk;
  assign {dlm1_wdata, dlm0_wdata}     = pyxv3lgda85n;
  assign k90knfo82df2l                    = {dlm1_rdata,dlm0_rdata};
  
  ad3c301j_tm48vb7x3
   #(
      .nm_fj         (16),
      .onr7l         (64),
      .h1b         (8),
      .ktra3i     (3),
      .rm39njpb7w     (13),
      .wvmre88     (64),
      .bf0ngee0t   (2),
      .xbpsp4_i     (8),
      .k2qm7hpa_qinpd (0),
      .quofpn_rylwqbg9 (0) 
      ) ne52xlcv8rmv6ffeim1 (
    .vlb2az38tbnj4           (vlb2az38tbnj4),
    .ujj9wb8hyzso           (ujj9wb8hyzso),

    .eth8quxx9hhjhxr4u9k2s77f    (eth8quxx9hhjhxr4u9k2s77f  ),
    .zw6mbnvv_8hcztypnytp87v_vy    (zw6mbnvv_8hcztypnytp87v_vy  ),
    .l_s_khzs83700pzjuq3_obo44     (l_s_khzs83700pzjuq3_obo44   ),
    .tcrjx_8vlmtrlqjvk3tu     (tcrjx_8vlmtrlqjvk3tu   ),
    .y0jaju01t8mqh2ycz05limpxfu    (y0jaju01t8mqh2ycz05limpxfu  ),
    .x88dy7qz1z117o2jmbslutlpm    (x88dy7qz1z117o2jmbslutlpm  ),
    .xs2l1_f3yynnrl_rw2zbe     (xs2l1_f3yynnrl_rw2zbe   ),
    .kyvscpwy0vljnwysfxqxb    (kyvscpwy0vljnwysfxqxb),
    .sl5cpfvi658e8pl6nh2cm4    (sl5cpfvi658e8pl6nh2cm4),
    .tmqgi_fx924f3bq8ms4u8t0    (tmqgi_fx924f3bq8ms4u8t0),
    .hf8rqlrzsk0e9ho4orde_r    (hf8rqlrzsk0e9ho4orde_r  ),
    .opns8_xijy8grr0gygeszh    (opns8_xijy8grr0gygeszh  ),
    .hng3_y3ldjtyu4a9n45      (hng3_y3ldjtyu4a9n45    ),
    .y1ovf4ea_l0kgs84_pwk6czrs  (y1ovf4ea_l0kgs84_pwk6czrs), 
    .n6fa00b9i708mtqu7yc9wjvxip    (n6fa00b9i708mtqu7yc9wjvxip  ),


                              
    .d53gmmeaj           (r6tkd_53z   ),  
    .coouz2jyj2n         (cyop0l7lnv6j3 ), 
    .dcmn368x8          (g9h1mnhtsaduuk  ),
    .opsl7g4          (pyxv3lgda85n  ),          
    .tn65z3ytg         (k90knfo82df2l ),
    .wzor2kya          (             ),

  

    .gc4b3kdcan6do88ta_       (clkgate_bypass),
    .gf33atgy                  (imsbh3sgxkg4),
    .ru_wi                (rst_aon) 
  );











  ux607_clkgate mhtsj557yyputg_bi_c9(
    .clk_in   (core_clk     ),
    .clkgate_bypass(clkgate_bypass  ),
    .clock_en (dlm0_cs),
    .clk_out  (clk_dlm0_ram)
  );

  ux607_clkgate vy5bv707gz0f4_lr5vo9i(
    .clk_in   (core_clk     ),
    .clkgate_bypass(clkgate_bypass  ),
    .clock_en (dlm1_cs),
    .clk_out  (clk_dlm1_ram)
  );


wire [32-1:0] fcjh1nct4r = clic_int_mode ? irq_i[32-1:0]: 32'b0;
 d2x3825_dhbv0h #(
     .vb1dh27fsxbyysw (urjif1vu4pqgqxt4x8),
     .t5twosugmt3qlv (3)
 ) u_ux607_clic_top(
    .dk2xhkj77a                     (core_clk_aon),
    .gf33atgy                         (ais_l7yddpa00),
    .zh6e0v0mmz                    (core_clk),
    .ru_wi                       (rst_aon),

    .a3v1iy5k0                        (zmxoq9ga),
    .cjwv                        (mtip),
    .fcjh1nct4r                    (fcjh1nct4r),
    .th06du2c8e2_b7k               (ooqxby68qkbvkc5xteznb_x),
    .irjoi8wvo25u209f_5               (zhr6liff5rm5wfulyyq),
    .zvk11dhgg2s67mkq                (xlsvmbo_v42zk9mypgihxz[15:0]),
    .lhibcc3xwm6cy               (etkmv0abc25lclz_o85),
    .zxe59xihintdqfy9d                (ijehxhtls_byykogg4h),
    .u4r4b_6kp09q767q               (ylsn7ect00nktb3n8gy6),

    .klkflmsyyf5w7ar               (txrvwlqb8aeb5k6eo4p0tb2),
    .wy36iirxspfw56864               (q8mbpl9ben1u54xn_d),
    .h7f6k_ims_9p3               (rsvzuajc8qp4__n0807),
    .lkjqs6kiuyj                 (igk23ds0cu4_sziqf),

    .aw82i964do                      (aw82i964do            ),
    .fbzs0o4ysyuzeg_qdj               (pzv82u11m6kxelyx220ilq5),
    .me1n4pvwxa7n3u8l05               (yhhbbaf9pqjys_bjgq6h4gj),
    .qaidts35dk5jcji0n               (qbaqr2mf9nkictp7plgs),
    .y8_gkxsfle                      (y8_gkxsfle            ),
    .fzdb65fcrotwcaccus_cwo           (fzdb65fcrotwcaccus_cwo ),
    .tcy_87vt9vet39knuw            (tcy_87vt9vet39knuw  ),
    .fc_4ns_w1nh4h02z_dgg          (fc_4ns_w1nh4h02z_dgg),
    .jqsukc5b5drcc1e78              (jqsukc5b5drcc1e78    ),
    .gnn46rd7vvofruqij              (gnn46rd7vvofruqij    ),

    .dz0zrf512290tvcy4q              (dz0zrf512290tvcy4q),
    .gfy3zost37aq8qmr                 (core_in_int ), 
    .dn8riluj40uunvq5               (clic_int_mode),
    .dxi_ue3gf5zqqqxwgq2a           (mnxti_valid_taken),
    .y12wg4mlovhn13                 (y12wg4mlovhn13),
    .kfrxhvr3mwznw                  (clic_irq_r),
    .b4lwcgm6l21pi                 (clic_irq_id),
    .zwcbp7zqfei5xz                (clic_irq_shv),
    .f_i1959b4xizzq9jea            (mintstatus_mil_r),
    .hjrk_rwjkqj3zk_b                (clic_irq_lvl),
    .znzjygllppv1s0a8cqub3c           (znzjygllppv1s0a8cqub3c)
  );

wire [32-1:0] t71as51n = irq_i;

 qc2dx_wo71_o92_z4 xkuia9tavvagp7ghtg(

    .v9ov1b3vn5k4ctkb     (sc9dq6vpj_vb3unfw0),
    .ub9pjiu4juf6nuqoq2w6     (ni7lsi0fuchbbgfizw0l),
    .aw0a19a967dn7n0x25w      (cvmgqobwfiy_kwo814x ),
    .ty6a2k41y0e9ir8_yzg     (h_htd26ozpf1rjy0gsvy),
    .cwkq4r6_upg_2884r     (gbzyzsndu75k8rua21_v9c),
    .ogvavqa7ta836s      (w2e5ixihsvl50pgq6b4 ),
    .sc169gxpr38lpe8     (tl_6em2dyajt9yrv4j794c),
    .hg1g2yh6yktfe_btdst7     (mf1rr9vurug23q2qsrv),
    
    .dy9ll1o6t6ytby71hf4     (m1vcvvn1ntgzmmwe1bse),
    .ow4hbh48f0mt6le4o     (f20ikomgiyzoonhphcz),
    .uzwj715coelxmfqs       (q7emifz3jwxt_jv0_w  ),
    .dek0xt7q6guk2vf6     (l1hbm4iglo7pz0pdg_ayjs),

    .da_yai4b0c6          (t71as51n),

    .qszs2_0t9_mzkmv3         (c4boo209),
    .x_cq40qmp6a         (x_cq40qmp6a),
    .ysjo7jpbga9zbsp         (yukl2),

    .b13zu8ysd3u         (b13zu8ysd3u),
    .dk2xhkj77a             (core_clk_aon),
    .gf33atgy                 (itcmps0ezqld),
    .ru_wi               (rst_aon) 
  );


ux607_tmr_top u_ux607_tmr_top(
    .i_icb_cmd_valid     (l9z66pxhit_o_1iyjp),
    .i_icb_cmd_ready     (jdh22q4xq9e7wiznv),
    .i_icb_cmd_addr      (y_z_yc9_f4ppblmsch3z5 ),
    .i_icb_cmd_read      (nmp2x4e8pl59l6he_f9_ ),
    .i_icb_cmd_wdata     (dd_gpw58ph81_864rnspr),
    .i_icb_cmd_wmask     (nhzg88_kzsk0fbtrtku),
    .i_icb_cmd_mmode     (yc7tq3wh6q569ueq7i07em),
    .i_icb_cmd_smode     (yfy18a1ju6mptqd0_u),
    .i_icb_cmd_dmode     (gducqncehu9g7n4lydij_0),
    
    .i_icb_rsp_valid     (ixpwz6oo67i61vepd74),
    .i_icb_rsp_ready     (t7hb1k3tkjzooetwf),
    .i_icb_rsp_err       (da2pgeraioxt6edc  ),
    .i_icb_rsp_rdata     (u2fwd1l2_bdiuiftn),

    .tmr_irq             (mtip),
    .sft_irq             (msip),

    .sft_rst_req         (de1sbr3kjbswue),

    .rtc_toggle_a        (mtime_toggle_a),
 
    .mtime               (nwk1l6uz4),
    .mtimeh              (ir_9aedxd8),

    .dbg_stoptime        (q4gqhurcazjpsf4h),

    .tmr_active          (b7ch4h6nrw1vm0),
    .clk                 (rcernpf1zf4   ),
    .clk_aon             (core_clk_aon   ),

    .rst_n               (rst_aon) 
  );







  
  
  
  
  
  

  
  
  
  
  
  




endmodule




















module hdkje04yactero (
    output sfyn3seo6gs,
    output sgthjbo1oq1kw1e6,
    output [64-1:0] ollg7,
    output d3n7pwgwcgze9cr4,
    output [64-1:0] amc4c8vcbecv1i,  
    output pby60vfdze02,
    output [64-1:0] vm3pyzc9nt95,
    output rbz4pv_atxqopdwt,
    output [64-1:0] qs1xgat7r8xow,

    output av1w8ld09cfofn,
    output im2b5l0h98avl6t4sj,
    output bw65wl7fvekfymd8vqx,
    output [64-1:0] pecbpcoa04vq,
    output [64-1:0] tb_snaxyfs,
    output [64-1:0] zc4mldgm25r,
    output [32-1:0] d23wb5yh1iyvf,
    output [1:0] srim3bfnzhve,
    output cy3nuhzm_v2p73mt,  
    output fvqwdz2hdbb,
    input  a02zzbowpjn06h,
    input  io5ukym11gp2utw,
    input  w41ourymsjpvm8q1e,
    output u_ll4hq1b12s2i1    ,









































































  input  svlxg92fk8wh7_jgsa8x,
  input  i_x3a8jgmo8qd81tcr,

  input   uc5qxb4d2b28ye5,
  output  o2qkf90r783,

  output habgbg2jn3qi,
  output dg4hzu_,
  output h7fseh5_df0hbx,










  output tw5xnp59d8x,
  output  um8zsjyxn_4p,  


  input  [64-1:0] wd9dvepxj,

  input  [64-1:0] v09gw6e6rfjf05qg,
  input fcjh1nct4r,
  output [7:0] f_i1959b4xizzq9jea,
  input [9:0] b4lwcgm6l21pi,
  input [7:0] hjrk_rwjkqj3zk_b,
  input zwcbp7zqfei5xz,
  input znzjygllppv1s0a8cqub3c, 
  output gfy3zost37aq8qmr,
  output dz0zrf512290tvcy4q,
  output dxi_ue3gf5zqqqxwgq2a,
  output ix299qulxi5, 
  output jjj61w03m77lv,
  output dn8riluj40uunvq5,
  output aw82i964do,
  output fzdb65fcrotwcaccus_cwo,
  output [7:0] tcy_87vt9vet39knuw,
  input  fc_4ns_w1nh4h02z_dgg,
  input  jqsukc5b5drcc1e78,
  input  gnn46rd7vvofruqij,
  output y8_gkxsfle,
  output x_cq40qmp6a,
  output z1l80uwh6vyyg34,
  input  rn1o3sl83,
  input  zz5wo47gw146x4,
  input  fgr486jx5kevbua,
  input  pvfk1_6o89lmby,
  input  xx87vzbpchg,

  
  
  input  c5ewdqztjw9za,
  input  rn2mt6nngsc9w5cz,

  output j0qaxhuqtdi,
  output pbzpk52jinfscit4mm,
  output gwj6ow6qvbhs0tc31,
  output iwdkm52x_w4hpak_a2_w,
  output [12-1:0] mm0ssgy582fv_j,
  output [64-1:0] ir2913p9xpmq_1bvfd1,
  input  [64-1:0] bsjo0v5e0t556pph,
  input  mwegg_7inaca6povsw,
  input  wnkp7091zrsevkbl,


  input  [64*4-1:0] azll7rq5fab5ou,
  input  [64*4-1:0] n6a0r_0zddzrme8,
  output ns0i7siujgkrghjpqv6,



  output  [64-1:0] qeb3z0x5,
  output  ibhfuwrztbm8p4gg,
  output  [3-1:0] i8_5wt0vppx,
  output  osv2437qj_3nuf,


  output  b7g_vsn0zoewh6g1,
  output  [2-1:0] onnv64ydiajl,
  input   [2-1:0] r21i4by0bu3ks,
  input  [64-1:0] hn85hkp2yav,

  input  pydatzxqqi,
  input  t5trf35s8vy,
  input  zbac123pv78sbz3,
  input  z4e_m564fxae0kpbjr,
  input  zmwq3e9oijvo7d7,
  input  hixy2y36a1pn0,
  input  ozwene1gdpatk6g,
  input  sxvvsxtbhyvt,

  output [8*32-1:0] pcr4upio7_tx37, 
  output [8*1-1:0] uzklqlncpqqm1rav,
  output [8*1-1:0] ortueunvnkx_l5m_j,
  output [8*1-1:0] hwuhtb7ucto_utk56,
  output [8*2-1:0] i1env2kmns7qvvuuc,
  output [8*1-1:0] g3s3vpafvy3i,






  output                         l9z66pxhit_o_1iyjp,
  input                          jdh22q4xq9e7wiznv,
  output  [32-1:0]  y_z_yc9_f4ppblmsch3z5, 
  output                         nmp2x4e8pl59l6he_f9_, 
  output                         yc7tq3wh6q569ueq7i07em, 
  output                         yfy18a1ju6mptqd0_u, 
  output                         gducqncehu9g7n4lydij_0, 
  output  [32-1:0]               dd_gpw58ph81_864rnspr,
  output  [4-1:0]                nhzg88_kzsk0fbtrtku,

  input                          ixpwz6oo67i61vepd74,
  output                         t7hb1k3tkjzooetwf,
  input                          da2pgeraioxt6edc  ,
  input  [32-1:0]                u2fwd1l2_bdiuiftn,

  output                         ooqxby68qkbvkc5xteznb_x,
  input                          zhr6liff5rm5wfulyyq,
  output  [32-1:0]  xlsvmbo_v42zk9mypgihxz, 
  output                         pzv82u11m6kxelyx220ilq5, 
  output                         yhhbbaf9pqjys_bjgq6h4gj, 
  output                         qbaqr2mf9nkictp7plgs, 
  output                         ijehxhtls_byykogg4h, 
  output  [32-1:0]       ylsn7ect00nktb3n8gy6,
  output  [4-1:0]    etkmv0abc25lclz_o85,
                               
  input                          txrvwlqb8aeb5k6eo4p0tb2,
  output                         q8mbpl9ben1u54xn_d,
  input                          igk23ds0cu4_sziqf  ,
  input   [32-1:0]       rsvzuajc8qp4__n0807,

  output                         sc9dq6vpj_vb3unfw0,
  input                          ni7lsi0fuchbbgfizw0l,
  output  [32-1:0]  cvmgqobwfiy_kwo814x, 
  output                         h_htd26ozpf1rjy0gsvy, 
  output                         gbzyzsndu75k8rua21_v9c, 
  output                         w2e5ixihsvl50pgq6b4, 
  output  [32-1:0]       tl_6em2dyajt9yrv4j794c,
  output  [4-1:0]    mf1rr9vurug23q2qsrv,
                               
  input                          m1vcvvn1ntgzmmwe1bse,
  output                         f20ikomgiyzoonhphcz,
  input                          q7emifz3jwxt_jv0_w  ,
  input   [32-1:0]       l1hbm4iglo7pz0pdg_ayjs,

  output                         x0i6aykuzxn1t7_hyw9s7r4to,
  input                          pbyudse8quydhisrzo9pbl4,
  output [16-1:0]   vapgj050raiah87lnzt_a, 
  output                         cvksl3f95u8b10a3rmr6qvom,
  output                         togorwkvhfveb6zwndvww,
  output                         i036i6j05gm5ht39aak7k,
  output                         xubhke6y45gk7d9bj7c1022icq,
  output                         nao0kbyh1yex0kg7uycyc,

  input                          c8u60qjfyfel53grl6lmf5_3, 
  input                          vhl77l_vrkmhgbq9nx8p8ix,   
  input  [64-1:0]        sedkfhar7baq5_wmvydzjmit2, 
  input                          sf4u33sbbh0akueinpc6j4ly8ue,   


  output                        bm7mey1b6dibd5i6lfpukeue,

  output                        a8h5u6ohzhowdrvqrnlllzd70h,
  input                         pz92yc3xo60c49ayrztvq18a,
  output [16-1:0]  pwzrcrecvxehn8htjdn3kv2d0, 
  output                        m5itqssum7ljklhpn5nvzvd93, 
  output [64-1:0]       kkk0rwd1njowzq01nvxke,
  output [8-1:0]    a2kttuidwhopy02uoajaf,
  output                        g4hx0dbyp7f7ou8x02a0,
  output                        zce_icdtm3r9hzeanwhlu3fv,
  output [1:0]                  jkp1oke9n1q9ikytwx_7k,
  output                        ksa323b46ngmxwazg70t76,
  output                        bs4xe3ath5_4_iwylkfwppp,
  output                        njyud2m27xz7r6j0g0ieq17m,

  input                         mu3ut_ezr05qz2bbi7_vc_aod,
  output                        sk3bm3yc69h4ac84pc4killh,
  input                         b7g_hkjxumf964flze01v6p  ,
  input                         cmtnwdaxz9zk1858kalga2vt  ,
  input  [64-1:0]        qjvmrd1013dapqkahq_f87b,



  output                         ndsqg7zrec89ncrv9yu3k,

  output                         eth8quxx9hhjhxr4u9k2s77f,
  input                          zw6mbnvv_8hcztypnytp87v_vy,
  output [16-1:0]   l_s_khzs83700pzjuq3_obo44, 
  output                         tcrjx_8vlmtrlqjvk3tu, 
  output [64-1:0]        y0jaju01t8mqh2ycz05limpxfu,
  output [8-1:0]      x88dy7qz1z117o2jmbslutlpm,
  output                         kykdx6vx9n3hm7k6oybv,
  output                         b59iokn7e2645ocyqifdk6sp1,
  output [1:0]                   xs2l1_f3yynnrl_rw2zbe,
  output                         kyvscpwy0vljnwysfxqxb,
  output                         sl5cpfvi658e8pl6nh2cm4,
  output                         tmqgi_fx924f3bq8ms4u8t0,

  input                          hf8rqlrzsk0e9ho4orde_r,
  output                         opns8_xijy8grr0gygeszh,
  input                          hng3_y3ldjtyu4a9n45  ,
  input                          y1ovf4ea_l0kgs84_pwk6czrs  ,
  input  [64-1:0]        n6fa00b9i708mtqu7yc9wjvxip,




  output                           v0bybbiepfqv4kc_cdg,  
  output                           i28_g1tt8nk7e30,  
  output [7-1:0] m_aqi5ytp0maje5sj, 
  output [54-1:0] e2iagwi42o6sun5_ykv9,          
  input  [54-1:0] wa_f05baz0i8dkq7t_4y,

  output                           hpf4dbs7lpgqzs89,  
  output                           hlpyb4rsu9gt28ml_u,  
  output [9-1:0] qh651fblp7os_lrh1rf5, 
  output [64-1:0] yalqjjffhlwhb4fi3re,          
  input  [64-1:0] s0j6brb1s7b0asp2o_4vmv0,

  output                           a9pfw7vdfvtnr1l89,  
  output                           qmlhx0ddtv5q5m65mb2,  
  output [7-1:0] gg035mahjzmwm_850rpfm, 
  output [54-1:0] faibzt_25z6u6lt9f,          
  input  [54-1:0] n_6989smoxxpesripwzs5,

  
  output                           pq_z6zyr2bjwut728ldr,  
  output                           p4ls8ac9eyqc7uznlkv,  
  output [9-1:0] utq6xdqs0m3irmvrgwe7, 
  output [64-1:0] tw7hzxhmmtptsxpzz1x9d17,          
  input  [64-1:0] tz_zq72t3w19dm7c3a0mu,




  input  f2qbwkn13kmm9hmrn159wahi,
  
  output                          mum8f1rtatle7p_55y84,  
  output [6-1:0]  pn5bpwlp5ijfako9m5ao,
  output                          g3s0qe2adsxsx8e6z ,
  output [24-1:0]  a1rl4lmhqp8ydyk07kqkn,          
  input  [24-1:0]  apnns9jlj7y3y5bg8ynz,
   
  output                          pmz7e4mgvbnmimqp0nghk,  
  output [6-1:0]  j61algpxjoycxbswhgsuf, 
  output                          omq1ehm8hp4q9jgp5n5vn ,
  output [24-1:0]  fbv1q6sraswzp91zcn,          
  input  [24-1:0]  jv8kv41vzuir6an4iod,


  
  
  output                          qgl4363n31jx6xjyo05zkn,  
  output [8-1:0] zec78nyllxlfwmpsgncluudf, 
  output [4-1:0] dwvnjl0vxqkgd8t6dtvg5z,
  output [32-1:0] gngmcj5c1jd85csel9ntru,          
  input  [32-1:0] tkt93y5lfluzkia5plvksp,
                                                
  output                          km7co8hqm563od8ga_03_g,  
  output [8-1:0] j4mas6g26o63wvnsdquh8c4p, 
  output [4-1:0] nniah5mh0cunkhyln9,
  output [32-1:0] rcy_v3911lf33nza5j,          
  input  [32-1:0] g4nfgu53_rgc0632w8z97,
                                                
  output                          xzgkclcxsgfuseg87,  
  output [8-1:0] djwlah5bo0r6myit6cal0t, 
  output [4-1:0] qu_ju3lv6nvkdbo8h11uf,
  output [32-1:0] dydwz9i6k80alqfarffop,          
  input  [32-1:0] ql1c7hzoj9kf__7r97krm,
                                                
  output                          kp2j8kv1p1cjcg0lerwm,  
  output [8-1:0] v4a7g1wh3ivw0esp7dye0oiz, 
  output [4-1:0] x9zuk21gpaj58uszvm5,
  output [32-1:0] n_h5oz0c5bo5rpevwjcu8,          
  input  [32-1:0] ryid4_99ns1jc83at_88x,



  output nv5a7f_68p9ebw,
  input  klwwlfrft,
  output bebngvg8sove,
  input  oi60pknul,

  input                                           moqs2k81l9fugde5v_581,
  output                                          i0acx70llka5qu09r5jd, 
  output                                          e44u8ctdv_z5u19to, 
  output                                          h7k_k0xxi7vktla, 
  output                                          v_vouzmjecsvtjxt, 
  output [66-1:0]               ef9y8yyld9onuy00de7o, 
  output [66-1:0]               ammhazyeeglt3ewt4p, 
  output [6-1:0]              xvwzwg7_3ek2tx, 
  input  [66-1:0]               y8sg6kbsyavoh4usiqn, 
  input  [66-1:0]               gnqkycbjc0k9k4_edoube, 



  
  input                             wh6iy6zpdqsnv2y,
  output                            bd6yatp5cqq,
  output [4-1:0]             fl1qsvyu,
  output [32-1:0]      b9889wezsu,
  output [7:0]                      an__mxugc4,
  output [2:0]                      poj6g8vw9e,
  output [1:0]                      dafaivw3ze9g3hi,
  output [1:0]                      q2c0d6fxz_1bw,
  output [3:0]                      wblesminvapwua,
  output [2:0]                      v3cim36gj8g,
  output [3:0]                      ss22f8fuy2uhr,
  output [3:0]                      hoaoalj5pcdnpnm0,
  output [1-1:0]               rh8f1e3jgg3xi,
  
  input                             roral7fym4h3_,
  output                            b_gwvq35iq0_yvk,
  output [4-1:0]             lqm2hm0cjm5zt,
  output [32-1:0]      f3n3tpjs44e0_,
  output [7:0]                      dmc59hxf352z,
  output [2:0]                      a63l3og_8qak5jy,
  output [1:0]                      m0wp58qmji79,
  output [1:0]                      c8qmnfk1vqai,
  output [3:0]                      pbov8g9yizcwr,
  output [2:0]                      t8qjehupeajtzjr,
  output [3:0]                      hhp1rh0x0jn,
  output [3:0]                      w9yptl69xj6p,
  output [1-1:0]               yvcpy_gyehs4lji, 

  input                             kted7ph0krq,
  output                            a93i3d2hji,
  output [4-1:0]             of5p5cb8p4,
  output [64-1:0]           g1bi1xzuv64,
  output [8-1:0]        gj6p5b5ik3r9p,
  output                            m1fmaas4oww6,
  
  output                            hjstsi51gm,
  input                             onpqhy0s69,
  input [4-1:0]              aw7xjbi,
  input [64-1:0]            z0cc2y_uzoh_,
  input [1:0]                       y8tc_vywu82ugn,
  input                             o2h9d51o6m6,
  
  output                            nneek3ep5xykwl,
  input                             g8khua4l0y77zjp,
  input [4-1:0]              wmlp1a2b,
  input [1:0]                       weop50xb_avne,

  input                            su81e8dxdzng9d,

 
  output [1:0]                   lueem7uei21mn66  ,  
  output                         vgodhub5af4gihqv5eef  ,  
  output [32-1:0]   lueqjwqinfpts52   ,  
  output [2:0]                   lv9moee8_5_8dsy5   ,  
  output [32-1:0]        ck0wbvgghs6n9j4  ,  
  output [3:0]                   uecfgtalcganlj42vmq   ,

  input  [32-1:0]        msxgfr_x73l96858p1s  ,  
  input  [1:0]                   tze074ath5y6h2m41   ,  
  input                          o752t3g6xbcxc6if88wi  ,  

  input                          nprvxoyk8ecm174bi8,


  output              wex3zbl1x6s4be1en,   
  output [1:0]        pszbl2iobld50k,   
  output              vfuu2l_7oof31qn0_a,   
  output [32    -1:0] bvy9o58rgxtbjz_xph,    
  output [2:0]        gcpthp2sfxb3cxo,
  output [2:0]        xzjdk5deciqs4l3my_l,
  output [3:0]        peug05ptx4vv93u4xc, 
  output [64    -1:0] dlg9f36umgj9xdv0wa,   
  input  [64    -1:0] yienty7ycnc25au,   
  input  [1:0]        rxlx2eq69oye0ba3,    
  input               j2amhrzbhku8dzd,  

  
  input                         fkm9up63o1aeauaqhjb,
  output                        to_1lv9wnb3vmu6tvz5rc,
  input  [32-1:0]  ju1kbeplcqy314lfj4, 
  input                         r985fbe5k7hgzaq9i, 
  input                         bb04gpwotp2s6c7_p1gqkq, 
  input                         sqmey185cu3mtixhl, 
  input                         rffcsd1o699ytclmx,
  input  [64-1:0]       lbr88vbqtg8rht7320frde,
  input  [8-1:0]    g7qq38mx3d58n1b15kcia,
  input                         demg_fwfkmaeawq30t,
  input                         grtb6ypa0px2gi1c,
  input  [1:0]                  f128d8ws0seoihu1,
  
  output                        m2r7mfmq3afdd1ine,
  input                         nhafiywg3hg_52kogwh,
  output                        xrqayy6vigrw66z8a  ,
  output                        jyy72ywt9nbo10f2jxupacld,
  output [64-1:0]       drz92qecqx_qtxwro,
  output                        st4f16aums5, 
  output                        p05ld2ghmwh, 


  input  [31:0]                  ij_sgq3rtvw2,
  input  [31:0]                  k9jntnqwqp,

  output bf61lpqg8z,
  input  dnl01g_,

  output wz_if_2q_23jhl2,
  input  n1wslu68m9v,

  output dyl5g2vgrvy4mb3,
  input  viuu21jzrv,

  output trtkzwpsx6l,
  input  h87jx93oz7,

  output emc_bywzarijbo,
  output h8xul8_er09on,
  output umnrzb6pv8dzc,
  output e592323mqvany, 

  output j4xe_w_yjq2,
  output j2t29hqv0s6c7,
  output aui65oshqn8b5_iz6,
  output jmoafuo8zb_i1t,
  output sa5of37yr6xn0s3e,
  input  o_dsdljul,
  input  juyzxopct4k03sl,
  input  qyqw_37_fxv8z,
  input  hyw0m71z3q3rpt1,
  input  fx_h7chccf02z,
  input  o5q5hev,
  input  c8fchlpwl,
  input  erv7j3wmd3gb_dp,
  input  fid1178x5nxb,
  input  dk2xhkj77a,

  input  gc4b3kdcan6do88ta_,
  input  ru_wi
  );


  wire xmbe_e4vm6ofjbn7lq;


  wire ifu_o_valid;
  wire ifu_o_ready;
  wire [32-1:0] ifu_o_ir;
  wire [64-1:0] ifu_o_pc;
  wire bcv5wwa3cpmh6o9d; 
  wire pbiupof7z_siv68x2; 
  wire eey8q1ex7jqqx0hm_; 
  wire hyzfgvg8iynh8zpa4; 
  wire mdfkn7idoni9xj; 
  wire v3pirqtitn2_xu9; 
  wire n0p5652lvx0qj1yuwu; 
  wire ddp4_khmuujfs; 
  wire m_7gx91ep6vkla; 
  wire iyoccmh9a_a2ov94o; 
  wire [5-1:0] s8mlhtj2pe58l;
  wire [5-1:0] eh7xldx93qn_e_ig;
  wire [5-1:0] mxxfa5sn2ahc21k;
  wire                         wp3ochi2x8_ljvjh;
  wire                         yzl1nx341x5d2p4;
  wire                         l11qpt1sf6a7;
  wire n3mz6a4lr36ftz11;
  wire [64-1:0] f2d4k4kxynjpd0gghqe140;
  wire [4*8-1:0] uuy2zpbrzrwdf432a7_g;
  wire [4*8-1:0] d4d7ru_yllps7en_tto;
  wire [7:0] ylmhlw32ex4fxli7;
  wire [7:0] n_lam8gs1mljgiq8zi;
  wire [2:0] v_97hsna5xll5n1xslwe3;
  wire [2:0] v2r90qa11qssvr5tq98dbi961;
  wire ba89afyz0al00;
  wire gkonom22e0fpa2_v3w0ab;
  wire [2-1:0] fxvpc9o9zl2t2nuwpg0;
  wire [2-1:0] gtvau5cygdmb10dr_makqf;
  wire qu31vl4s4x0pmeth2j_7neq1;
  wire himvp4q0erus0anat5;
  wire ps9l2wesoladg;

  wire y_0q8d40rrzolo1y6;
  wire ao17frh5wnr0wddz3;
  wire mmludd_fnt2yevok8a1a0;
  wire buwj9_8l8bwj80kkinq9p;

  wire hwpkcsh2atrq  ;
  wire v3e6l1k7eo9k3 ;
  wire hxrmt706n071lic0f7;
  wire tluzd_2baaw1fpd4o1td_h;
  wire agcvtek_6ocmw76d;
  wire [64-1:0] j0_nonyh_r387uiy;
  wire [9-1:0] p54semfzu2zyfb;
  wire [9-1:0] xosc7587i2hjow2yjw;
  wire zsgl59ydqwjln;
  wire b9yq2alidby7zgom1;


  wire tvqijouldcgiz2dxdco7;
  wire zkxlkidschdubxpkpm;
  wire xmcrni1qngfvh9pil9j;
  wire btkcf2uqr61gkiqhde0lai;
  wire [64-1:0] h01d94xsxbxe_req;  
  wire w1casjl7bz73brz;
  wire hjri7cufo9ckntq;
  wire yghffofulqa77bd7aw07badta1a;
  wire rrl7evvmayt1_vvp74iq9h6_cjf;
  wire [27-1:0] zddoxp22m1o11x30gbe;
  wire [16-1:0] hwfethpzkuauejcgtbl6o; 

  wire n3ak8l6cvn0s4;
  wire hsxh9536ho4bw8o;
  wire r_edve7v9jcr26q6zk;
  wire vrqfzuog2k4pos133;
  wire bmw2yi333716crywk;
  wire k2sr7sw1plcmnki5ajtscw;
  wire [64-1:0] jkzw_f9anx55;  
  wire t8muv9e6d7yk_whqa0;
  wire hzdfp71n6g3f5fsg5;
  wire lwdhmuzyvcvv14mjbl0h2a41z;
  wire xy48dugh009wtmazqug3kpy2a5h_;
  wire [27-1:0] l4ztejmt2__wxqm2rw;
  wire [16-1:0] s3ujdp2a8n69bm6engxok; 


  wire                                   gvkx7hystgemle; 
  wire                                   ii7h_yx8mmn1y82k; 
  wire [74-1:0] f71s92bjwuhpisqhx13nk; 
  wire                                   xrkn9p6pdpoya56pfoc6t; 
  wire [5:0]                             qqo7mp2z_os7tj0c4w6kf6y; 
  

  wire                                   mcfeo0u7nf9; 
  wire                                   sa3k3tsgxwqp8z; 
  wire [74-1:0] wfa5o72ctktgt55fgv2eo; 
  wire                                   igeg6alwzopr62ti9; 
  wire                                   g3e0lri_3krzlfxnnlo_2y82qf; 



  wire lln3b7iev7jpvogh964ro_9bc_3y;
  wire q97rqfy8n7ixfm2a5wev4nd5sylpcq3j;
  wire hujgg6hjnhtbspbkekuz5_u;
  wire v3pnt81kfrgbaanm1mhh51w;
  wire [64-1:0] i08eq60d_snxeq8si_ezod;
  wire y8wz7aud_fd6dfiakjtx2i0g;
  wire dgnjyd9xs8efyxm0tdlsvfq4eop;
  wire a3xib90kwk4_hm1;
  wire nfzexr8q9g893gi;
  wire [64-1:0] opkkwp3eg8g3448t;
  wire um28jgd2x4mbs;
  wire [64-1:0] l_imk5zs8ejjka;
  wire [64-1:0] lz3vnoxnz_z;
  wire yhbtmo4kyz_ewog3;
  wire cd4d2_i3rcc1_p;
  wire [5-1:0] wyu42gj62n994v0wo_;
  wire x9cmkt53yq483z1;
  wire cxmwxfttqy2t7ura   ;
  wire b5wruck8tj9sa   ;
  wire bxentpryfwb3d  ;
  wire o2a43mjdbgea1  ;

  wire dkmuhc79d2wm0wubp; 
  wire u2demhkod_er3kf6b; 
  wire uz7pt71lvqit85od; 
  wire [4-1:0] v3uvhtx7e5vbtvie;
  wire [64-1:0] tmqkgmlzi018;
  wire [64-1:0] lx_olubu7t8h;
  wire [64-1:0] dd1p3tnenmm9r;
  wire [3-1:0] l60zv02z95hlayri;
  wire l1xzyldaa9dr2q7mla;
  wire a5z_23_ryr_m29hhia_p ;

  wire vejdvgqormu727s;
  wire [64-1:0] ar9ro1ql86jzmq_p;
  wire [5-1:0] qz1gqv6vh5qturw6v1mz;

  wire y7rd1k0an54clel_5q6; 
  wire com03bquiktu249yb0; 
  wire [64-1:0] tzg0yjgx9bn98i;
  wire [5-1:0] x8_a2j7z3gz3l0tfjqp;
  wire [4 -1:0] c2mipfm_6z5ef4p3aoz;
  wire y3z8rf7c6hvsiux ; 

  wire xq0mj5mg2_512eu4; 
  wire e11m1298jo38qcwq9er2; 
  wire [64-1:0] ec94_mk193di7tj;
  wire [5-1:0] nodrapn01yl1vxle30p;
  wire [4 -1:0] m2sw40fca0wvnmy;
  wire ywhfwlbfro2dmuvf ;

  wire ex_g_cnadtiu1r9u;
  wire orzasugx5h5pio22_;
  wire [64-1:0] dxwtzud_wfj8jqk0;
  wire [5-1:0] dn074lh73rzchvrqzm8;
  wire [4 -1:0] gi8o690aydhqi8;
  wire zl1r9cfvuhltjq ;


  wire  rnx27onf2lbe  ;



  wire                         enwn0u48p2_ls5az80;
  wire                         miax48k27o484e8a;

  
  
  
  
  wire                                     moj77icm1kmex0900;                
  wire    [27-1:0]     hib0x0rvcjwnn75a;                
  wire    [1:0]                            cgmsm8wvxc5kg90xwvwq0cga;                
  
  wire                                     w9mx37ezcezieq_9__94o;          
  wire                                     hsnr3xtposirc7pmphtiko3xlz;     
  wire                                     k1jkhgd9bvypwrti7ietjp0n7_nyzu;   
  wire   [51-1:0]       qirelbyt49gkn46_f24yxtc;
  wire                                     jq4wiwydrozelhpru9snvs0;         
  wire                                     j6muxslh7pud3298q9d8lc2;         



  wire qo5p9t6s74zxpo;




































  wire                        x27lqkgq55knwoqsc6_bn0p;
  wire                        ud5ygg9b8pmm93drtbfk4l8hv;
  wire [64-1:0]   f_lrqmtz5mpqmbrhn6f05; 
  wire                        ss92bd8t5gyfjfl1_lp2;
  wire [2:0]                  z1beclu7k0_h4nn6njz05sbe1;
  wire [1:0]                  w1i6s2iwu2nnj7idywd;
  wire                        czjipv9hqkdx4jllt3ajsl;
  wire                        j92g3e8ublsg2d9sjj_i3;
  wire                        af3a5ot65per6f87crwmj;
  wire                        bjucsszqg5d1sc5etnwvf1;
  wire                        t37flu99i5ex1j3e_8   ;
  wire [1:0]                  wvjkzp74fi8ed7nnr7xlm3gt ;

  wire                        phzkntckzzbndu4wevf1o6;
  wire                        bpyef3a0dnkkyqdpymy  ;
  wire [64-1:0]       ba1ucnyekcm68i9wuqwmn;


  wire                                   bz8qao4o4xqslni1d3;
  wire  [27-1:0]           vpecdc5kos; 
  wire  [1:0]                            pccd7o463jfc_dpc5va; 
  wire                                   k5ovx8tintgvetip; 
  wire                                   f97le_hyejv7saw9vslna; 
  wire                                   yruel3nusosm39gnmb9ev_; 
  wire                                   oeux55k_cre0he7w7jip5b1; 
  wire   [55-1:0]     r8z2r_ud53zj8mrpk; 
  wire                                   bu1949pq_9946o1_e2q_uvr8p4; 
  wire                                   b4isf5u8b8pj34e09f72vxe38zg; 
  wire                                   kvpemhoim1tq5y8mzwvix5; 
  wire                                   docsdqb0rnb9fmmgf3; 
  wire                                   xyqctztl2_la5wbp2an04mw; 
  wire                                   du_nrgluldn3gf5tg1wa8slreks; 
  wire  [27-1:0]           w8mlksniwgqyojf1iy; 
  wire  [16-1:0]           vn9mhiqoo1jrmofqr4xn; 
  wire                                   b518xebdeds3frng6hy4g; 
  wire                                   z1l_kkshyf_56cwmaq2dm;
  wire                                   f1ofib7_3yq8rgwsltzwex = ~z1l_kkshyf_56cwmaq2dm;
  wire  [16-1:0]           w7u50np_chxy7wq5n9et_q;
  wire  [20-1:0]             l2dse4sd3runnrb1rcbydauc; 
  wire                                   kr1rhzlb5gr_wty1pe392s5oqet; 
  wire  [1:0]                            ox2ptuhum_e2aodz8wine6h; 
  wire                                   g_qmxgznvfin609fmm97kuc2dm02; 
  wire                                   i9oln6xm1pi9dzsd61s1kg4dmo7j; 
  wire  [1:0]                            hei_cs0rbwsv; 
  wire                                   yf_5vs18cke5xg660my; 
  wire                                   sneofd4rq3b0m9eu91r8;  

  wire                                   xib8tki1lzl05e71ry; 
  wire                                   hdle8ta5fimb1inf1z; 
  wire  [32-1:0]              trtxm7l0l_kp36i9y;
  wire  [1:0]                            p0akg_4worvsnfq_q36vp;
  
  wire                                   mqdc73rtez0bzh2_1;
  wire                                   vl5p5iump0rpm1hbr;
  wire                                   oj6rvjf7ujgb34264;
  wire                                   vjfz03uzu8p_0jhhvvev;
  wire                                   p1qeemcgwrrzzt73bl;
  wire                                   ertspxpg0txqgp9i6fx53;
  wire                                   z3xt8rx_qs6z0goo1;
  wire   [64-1:0]                ln7r12q36ofpcd6m6u;


  wire                         mfnb4b0       ;   
  wire                         edebnrit9_y77l ;   
  wire                         gbhvs__f9z_q97jj ;   
  wire                         hle5nop1tcht5cg ;   
  wire                         t7panq_mivym6dhmjp;   
  wire                         uaehep04469aadw4ga1;   
  wire                         op60_2nivpji1_v8upx;  
  wire [5-1:0] nzi6n_pc9q_5ybxyh;   
  wire [5-1:0] sqliqgffeni4u6uzs;   
  wire [5-1:0] gr8qapbswugbbkjl5;   


  wire n8mvs5sw2pw48loob7jv6nmjdds;
  wire dbzz2cu7abqy43de_ky433v;
  wire y3iin4ygz2ed73_84l91h73;
  wire gbb0bfnz8wqnjr5sufoh6ojt4pr;
  wire im70q80i1xh1y_5mo9ndr1 ;


  wire c4ughu0qm5sfai;

  wire w92a5o09fp9dg6   ;
  wire eglor15f7p2ivpny5dc   ;
  wire ous_emkpecrqhg5e7;
  wire doh50j3p7c7yl7uk9;
  wire s7eq8f6z1uyi2in;
  wire qbsr1jytrqtsbk4ttb8nz;

  w3yn55ly7roq dkjwc4tume0l(

    .s7eq8f6z1uyi2in   (s7eq8f6z1uyi2in),
    .qbsr1jytrqtsbk4ttb8nz(qbsr1jytrqtsbk4ttb8nz),

    .w92a5o09fp9dg6   (w92a5o09fp9dg6   ),
    .ous_emkpecrqhg5e7(ous_emkpecrqhg5e7),

    .c4ughu0qm5sfai   (c4ughu0qm5sfai),
    .tw5xnp59d8x     (tw5xnp59d8x   ),
    .aw82i964do       (aw82i964do),
    .y8_gkxsfle       (y8_gkxsfle),

    .pydatzxqqi     (pydatzxqqi),
    .enwn0u48p2_ls5az80    (enwn0u48p2_ls5az80),
    .miax48k27o484e8a    (miax48k27o484e8a),
      .pcr4upio7_tx37     (pcr4upio7_tx37   ), 
      .uzklqlncpqqm1rav  (uzklqlncpqqm1rav),
      .ortueunvnkx_l5m_j  (ortueunvnkx_l5m_j),
      .hwuhtb7ucto_utk56  (hwuhtb7ucto_utk56),
      .i1env2kmns7qvvuuc  (i1env2kmns7qvvuuc),
      .g3s3vpafvy3i  (g3s3vpafvy3i),

      .e1jv60iid34gonwyukkue                        (gvkx7hystgemle                          ),           
      .xz57o2ko5gkcbk8rq                       (f71s92bjwuhpisqhx13nk                     ),          
      .grv8y38uxakr22asia                      (ii7h_yx8mmn1y82k                          ),         
      .bvmb0d5jendar95w7nbnob8                  (xrkn9p6pdpoya56pfoc6t                ),           
      .h47i__o10wyo2sbyt58zq1_h5                   (qqo7mp2z_os7tj0c4w6kf6y                 ),           
      

      .vxwhhz9_cff6uy0x                           (f1ofib7_3yq8rgwsltzwex                 ), 
      .moj77icm1kmex0900                          (moj77icm1kmex0900                        ),                
      .hib0x0rvcjwnn75a                           (hib0x0rvcjwnn75a                         ),                 
      .cgmsm8wvxc5kg90xwvwq0cga                    (cgmsm8wvxc5kg90xwvwq0cga                  ),                 
      .w9mx37ezcezieq_9__94o                    (w9mx37ezcezieq_9__94o                  ),          
      .hsnr3xtposirc7pmphtiko3xlz               (hsnr3xtposirc7pmphtiko3xlz             ),     
      .k1jkhgd9bvypwrti7ietjp0n7_nyzu             (k1jkhgd9bvypwrti7ietjp0n7_nyzu           ),   
      .qirelbyt49gkn46_f24yxtc                     (qirelbyt49gkn46_f24yxtc                   ),           
      .jq4wiwydrozelhpru9snvs0                   (jq4wiwydrozelhpru9snvs0                 ),         
      .j6muxslh7pud3298q9d8lc2                   (j6muxslh7pud3298q9d8lc2                 ),         



    .h8xul8_er09on      (h8xul8_er09on),
    .wd9dvepxj        (wd9dvepxj),  





































    .x0i6aykuzxn1t7_hyw9s7r4to    (x0i6aykuzxn1t7_hyw9s7r4to  ),
    .pbyudse8quydhisrzo9pbl4    (pbyudse8quydhisrzo9pbl4  ),
    .vapgj050raiah87lnzt_a     (vapgj050raiah87lnzt_a   ),
    .cvksl3f95u8b10a3rmr6qvom    (cvksl3f95u8b10a3rmr6qvom  ),
    .togorwkvhfveb6zwndvww    (togorwkvhfveb6zwndvww  ),
    .i036i6j05gm5ht39aak7k    (i036i6j05gm5ht39aak7k  ),
    .xubhke6y45gk7d9bj7c1022icq    (xubhke6y45gk7d9bj7c1022icq  ),
	.nao0kbyh1yex0kg7uycyc      (nao0kbyh1yex0kg7uycyc    ),
                                                     
    .c8u60qjfyfel53grl6lmf5_3    (c8u60qjfyfel53grl6lmf5_3  ),
    .vhl77l_vrkmhgbq9nx8p8ix      (vhl77l_vrkmhgbq9nx8p8ix    ),
    .sedkfhar7baq5_wmvydzjmit2    (sedkfhar7baq5_wmvydzjmit2  ),
    .sf4u33sbbh0akueinpc6j4ly8ue   (sf4u33sbbh0akueinpc6j4ly8ue ), 
                                                    

    .ozt73ngxbaqnefsu        (rnx27onf2lbe        ), 

    .m6dcbta00ca03    (),
    .c06dvphgeptbqa    (),
    .t2e9t5kf8lqaa82dtg(),
    .viaoqex1en8ydnwh5(),
    .st9v6ljxhtiqln7(),
    .sehjrvl7lsqlkpl8js(),
    .owbvtem77_l_b4(),
    .crywtg_a3ctx3707n(),


    .h9zak9fmm8rw         (mfnb4b0       ),   
    .xvhg384tm4h76gdzx   (edebnrit9_y77l ), 
    .hdlty51ir9snk3qql9ow   (gbhvs__f9z_q97jj ), 
    .e0bgl8ntt8sp5j7o1yo   (hle5nop1tcht5cg ), 
    .ifg_e4rrluhhouqgceuo2  (t7panq_mivym6dhmjp), 
    .sz1c6k4c7y75fhzt1m81q  (uaehep04469aadw4ga1), 
    .y_g5vz_1yjpqe371ks  (op60_2nivpji1_v8upx), 
    .y88swlv8vqatvrurk392  (nzi6n_pc9q_5ybxyh), 
    .yx32lmcp5paz31u5hecbq  (sqliqgffeni4u6uzs), 
    .pktjjlrrkgnqgrqag  (gr8qapbswugbbkjl5), 








    .yoo3wc2tlwfyc6            (ifu_o_valid         ),
    .f78zm1o77tcsokzo            (ifu_o_ready         ),
    .z0o61mxkm788c               (ifu_o_ir            ),
    .pm7xlj7bu           (ifu_o_pc        ),
    .bcv5wwa3cpmh6o9d         (bcv5wwa3cpmh6o9d      ),
    .pbiupof7z_siv68x2         (pbiupof7z_siv68x2      ),
    .eey8q1ex7jqqx0hm_         (eey8q1ex7jqqx0hm_      ),
    .hyzfgvg8iynh8zpa4           (hyzfgvg8iynh8zpa4        ),
    .mdfkn7idoni9xj          (mdfkn7idoni9xj       ), 
    .v3pirqtitn2_xu9           (v3pirqtitn2_xu9        ), 
    .n0p5652lvx0qj1yuwu       (n0p5652lvx0qj1yuwu    ), 
    .ddp4_khmuujfs           (ddp4_khmuujfs        ), 
    .m_7gx91ep6vkla           (m_7gx91ep6vkla        ), 
    .iyoccmh9a_a2ov94o         (iyoccmh9a_a2ov94o      ), 
    .s8mlhtj2pe58l           (s8mlhtj2pe58l        ),
    .eh7xldx93qn_e_ig           (eh7xldx93qn_e_ig        ),
    .mxxfa5sn2ahc21k           (mxxfa5sn2ahc21k        ),
    .wp3ochi2x8_ljvjh            (wp3ochi2x8_ljvjh         ),
    .yzl1nx341x5d2p4            (yzl1nx341x5d2p4         ),
    .l11qpt1sf6a7            (l11qpt1sf6a7         ),
    .n3mz6a4lr36ftz11       (n3mz6a4lr36ftz11    ),
    .f2d4k4kxynjpd0gghqe140      (f2d4k4kxynjpd0gghqe140   ),
    .uuy2zpbrzrwdf432a7_g     (uuy2zpbrzrwdf432a7_g  ),
    .d4d7ru_yllps7en_tto     (d4d7ru_yllps7en_tto  ),
    .ylmhlw32ex4fxli7         (ylmhlw32ex4fxli7       ),
    .n_lam8gs1mljgiq8zi         (n_lam8gs1mljgiq8zi       ),
    .v_97hsna5xll5n1xslwe3    (v_97hsna5xll5n1xslwe3),
    .v2r90qa11qssvr5tq98dbi961  (v2r90qa11qssvr5tq98dbi961),
    .ba89afyz0al00          (ba89afyz0al00        ),  
    .gkonom22e0fpa2_v3w0ab       (gkonom22e0fpa2_v3w0ab     ),  
    .fxvpc9o9zl2t2nuwpg0      (fxvpc9o9zl2t2nuwpg0    ),  
    .gtvau5cygdmb10dr_makqf      (gtvau5cygdmb10dr_makqf    ),  
    .qu31vl4s4x0pmeth2j_7neq1  (qu31vl4s4x0pmeth2j_7neq1),
    .himvp4q0erus0anat5       (himvp4q0erus0anat5    ),
    .ps9l2wesoladg             (ps9l2wesoladg           ),

    .p0olq02_hyvx0           (y_0q8d40rrzolo1y6),
    .mneths0pu5slsnpiv           (ao17frh5wnr0wddz3),
    .hwpkcsh2atrq            (hwpkcsh2atrq  ),
    .v3e6l1k7eo9k3           (v3e6l1k7eo9k3 ),
    .hxrmt706n071lic0f7          (hxrmt706n071lic0f7),
    .v7rzl8qveorn2jg6659m69   (tluzd_2baaw1fpd4o1td_h),
    .v_k8ohy_e2e9vlp6az04    (agcvtek_6ocmw76d),
    .y_vw514j6xmphhfhc       (j0_nonyh_r387uiy),
    .p54semfzu2zyfb          (p54semfzu2zyfb),          
    .xosc7587i2hjow2yjw          (xosc7587i2hjow2yjw),          
    .zsgl59ydqwjln         (zsgl59ydqwjln      ),
    .b9yq2alidby7zgom1         (b9yq2alidby7zgom1      ),


    .tvqijouldcgiz2dxdco7    (tvqijouldcgiz2dxdco7),
    .zkxlkidschdubxpkpm    (zkxlkidschdubxpkpm),
    .xmcrni1qngfvh9pil9j    (xmcrni1qngfvh9pil9j),
    .btkcf2uqr61gkiqhde0lai    (btkcf2uqr61gkiqhde0lai),
    .h01d94xsxbxe_req          (h01d94xsxbxe_req),  
    .w1casjl7bz73brz      (w1casjl7bz73brz),
    .hjri7cufo9ckntq      (hjri7cufo9ckntq),
    .yghffofulqa77bd7aw07badta1a  (yghffofulqa77bd7aw07badta1a  ),
    .rrl7evvmayt1_vvp74iq9h6_cjf(rrl7evvmayt1_vvp74iq9h6_cjf),
    .zddoxp22m1o11x30gbe      (zddoxp22m1o11x30gbe      ),
    .hwfethpzkuauejcgtbl6o    (hwfethpzkuauejcgtbl6o    ),  

    .n3ak8l6cvn0s4           (n3ak8l6cvn0s4     ),
    .hsxh9536ho4bw8o           (hsxh9536ho4bw8o     ),
    .r_edve7v9jcr26q6zk      (r_edve7v9jcr26q6zk),
    .vrqfzuog2k4pos133      (vrqfzuog2k4pos133),
    .bmw2yi333716crywk      (bmw2yi333716crywk),
    .k2sr7sw1plcmnki5ajtscw      (k2sr7sw1plcmnki5ajtscw),
    .jkzw_f9anx55            (jkzw_f9anx55      ),
    .t8muv9e6d7yk_whqa0        (t8muv9e6d7yk_whqa0),
    .hzdfp71n6g3f5fsg5        (hzdfp71n6g3f5fsg5),
    .lwdhmuzyvcvv14mjbl0h2a41z  (lwdhmuzyvcvv14mjbl0h2a41z  ),
    .xy48dugh009wtmazqug3kpy2a5h_(xy48dugh009wtmazqug3kpy2a5h_),
    .l4ztejmt2__wxqm2rw      (l4ztejmt2__wxqm2rw      ),
    .s3ujdp2a8n69bm6engxok    (s3ujdp2a8n69bm6engxok    ),  

    .lln3b7iev7jpvogh964ro_9bc_3y  (lln3b7iev7jpvogh964ro_9bc_3y),
    .q97rqfy8n7ixfm2a5wev4nd5sylpcq3j (q97rqfy8n7ixfm2a5wev4nd5sylpcq3j),
    .hujgg6hjnhtbspbkekuz5_u         (hujgg6hjnhtbspbkekuz5_u),         
    .v3pnt81kfrgbaanm1mhh51w          (v3pnt81kfrgbaanm1mhh51w ),         
    .i08eq60d_snxeq8si_ezod         (i08eq60d_snxeq8si_ezod),
    .y8wz7aud_fd6dfiakjtx2i0g  (y8wz7aud_fd6dfiakjtx2i0g),
    .dgnjyd9xs8efyxm0tdlsvfq4eop (dgnjyd9xs8efyxm0tdlsvfq4eop),
    .a3xib90kwk4_hm1         (a3xib90kwk4_hm1),         
    .nfzexr8q9g893gi          (nfzexr8q9g893gi ),         
    .opkkwp3eg8g3448t         (opkkwp3eg8g3448t),

    .um28jgd2x4mbs             (um28jgd2x4mbs), 
    .l_imk5zs8ejjka              (l_imk5zs8ejjka    ),
    .lz3vnoxnz_z             (lz3vnoxnz_z   ),
    .yhbtmo4kyz_ewog3           (yhbtmo4kyz_ewog3 ),
    .cd4d2_i3rcc1_p          (cd4d2_i3rcc1_p),
    .wyu42gj62n994v0wo_          (wyu42gj62n994v0wo_),
    .x9cmkt53yq483z1         (x9cmkt53yq483z1),
    .cxmwxfttqy2t7ura            (cxmwxfttqy2t7ura   ),
    .b5wruck8tj9sa            (b5wruck8tj9sa   ),
    .bxentpryfwb3d           (bxentpryfwb3d  ),
    .o2a43mjdbgea1           (o2a43mjdbgea1  ),

    .svlxg92fk8wh7_jgsa8x    (svlxg92fk8wh7_jgsa8x),

    .ldqpjrsj9dp8yg3uc       (v0bybbiepfqv4kc_cdg   ),
    .s70e4xdis3p67ndpn6fbx       (i28_g1tt8nk7e30   ),
    .h9zlka3j3ih8ihpvwvky1     (m_aqi5ytp0maje5sj ),
    .tf_tmpul8i8qbm_djvtl5f      (e2iagwi42o6sun5_ykv9  ),        
    .qtsqtuxyont41a7h7i6     (wa_f05baz0i8dkq7t_4y ),
                                                
    .w0ve66vjdz8lzwws3ic       (hpf4dbs7lpgqzs89   ),
    .df775k2ts6dn4528iq_ce5       (hlpyb4rsu9gt28ml_u   ),
    .k3dychuj1pv4vw7cfj01ft8v     (qh651fblp7os_lrh1rf5 ),
    .jh4zf96qrsb31j072n      (yalqjjffhlwhb4fi3re  ),        
    .vfvtxk4jkkc3ql7_rqd     (s0j6brb1s7b0asp2o_4vmv0 ),
                                                
    .hv6xxz3oswj4wy4j46       (a9pfw7vdfvtnr1l89   ),
    .q6p7kcdd9o7j3e2c886       (qmlhx0ddtv5q5m65mb2   ),
    .ee_yaeclihal4dht69liwy6z     (gg035mahjzmwm_850rpfm ),
    .thl4cxcuzntax8hnsn9bl4      (faibzt_25z6u6lt9f  ),        
    .mysqpp41yovfcis6f2dza47     (n_6989smoxxpesripwzs5 ),
                                                
    .vp3x08mx4e27x4k26n       (pq_z6zyr2bjwut728ldr   ),
    .a7b829uahvy2i28yzgg       (p4ls8ac9eyqc7uznlkv   ),
    .kzxrmeg90fb06oya08h1     (utq6xdqs0m3irmvrgwe7 ),
    .kl5wycr14v5ukl7oqfhwe6      (tw7hzxhmmtptsxpzz1x9d17  ),        
    .wt6c82_zmqgmt7if41t698     (tz_zq72t3w19dm7c3a0mu ),
 
                                            
 
    .i_x3a8jgmo8qd81tcr (i_x3a8jgmo8qd81tcr),


    .wz_if_2q_23jhl2 (wz_if_2q_23jhl2),
    .n1wslu68m9v    (n1wslu68m9v   ),

    .x27lqkgq55knwoqsc6_bn0p    (x27lqkgq55knwoqsc6_bn0p), 
    .ud5ygg9b8pmm93drtbfk4l8hv    (ud5ygg9b8pmm93drtbfk4l8hv),
    .f_lrqmtz5mpqmbrhn6f05     (f_lrqmtz5mpqmbrhn6f05 ),
    .ss92bd8t5gyfjfl1_lp2     (ss92bd8t5gyfjfl1_lp2 ),
    .czjipv9hqkdx4jllt3ajsl    (czjipv9hqkdx4jllt3ajsl),
    .j92g3e8ublsg2d9sjj_i3    (j92g3e8ublsg2d9sjj_i3),
    .af3a5ot65per6f87crwmj    (af3a5ot65per6f87crwmj),
    .t37flu99i5ex1j3e_8       (t37flu99i5ex1j3e_8   ),
    .wvjkzp74fi8ed7nnr7xlm3gt     (wvjkzp74fi8ed7nnr7xlm3gt ),
    .bjucsszqg5d1sc5etnwvf1    (bjucsszqg5d1sc5etnwvf1),
    .z1beclu7k0_h4nn6njz05sbe1    (z1beclu7k0_h4nn6njz05sbe1),
    .w1i6s2iwu2nnj7idywd     (w1i6s2iwu2nnj7idywd ),

    .phzkntckzzbndu4wevf1o6    (phzkntckzzbndu4wevf1o6), 
    .bpyef3a0dnkkyqdpymy      (bpyef3a0dnkkyqdpymy  ),
    .ba1ucnyekcm68i9wuqwmn    (ba1ucnyekcm68i9wuqwmn),

    .j8cjhcuf0m6xjvemdaz       (gbb0bfnz8wqnjr5sufoh6ojt4pr), 
    .umc_2tn6um_9xaiy7_ksg0w     (n8mvs5sw2pw48loob7jv6nmjdds), 
    .uiyh4da4134sjv7gnmc     (dbzz2cu7abqy43de_ky433v), 
    .q7ru87fmzxczveihcxcwh     (y3iin4ygz2ed73_84l91h73), 
    .s_eowfyzlvx7gjv542upo      (im70q80i1xh1y_5mo9ndr1 ), 

    .d40pep591l63yhmefp7i        (kvpemhoim1tq5y8mzwvix5      ),

    .t57d026x085pay         (docsdqb0rnb9fmmgf3       ),
    .k5th293qdrtsytaehbsk        (b518xebdeds3frng6hy4g      ),
    .g6gwjq519o1w1m3csgrrf3    (xyqctztl2_la5wbp2an04mw  ),
    .lo_2ny7_v71by78q3          (w8mlksniwgqyojf1iy        ),
    .hbdj3fcr8qkfkgzq58o1o2ozh  (du_nrgluldn3gf5tg1wa8slreks),
    .m_k_n75bb0f_im9fu_        (vn9mhiqoo1jrmofqr4xn      ),

    .bf61lpqg8z (bf61lpqg8z),
    .dnl01g_    (dnl01g_   ),

    .gc4b3kdcan6do88ta_         (gc4b3kdcan6do88ta_),
    .o5q5hev                (o5q5hev  ),
    .ru_wi                  (ru_wi         ) 
  );

  
  
  
  
  
  
  
  
  wire  [48-1:0] k9lv9ppimt14qx3d7rj;  
  wire  [64-1:0] llskuqv0ehm60atlo;
  wire  oug11blpzcta8zyu0ya;
  wire  zr1pc8tfxyljdj7a8a3eh5;
  wire  qg9g70jgx5r5l_wpc7;
  wire  o_qquv0pnx4zpz4h3gwxgl3;
  wire  j1fek3jzmt5bhhpnhvrmgt;
  wire  ds75nafgmrespy002qvcsb8;
  wire [5-1:0] jc4yg1pkylr2gonwcd;   
  wire [5-1:0] nd3cgvec1pogf2;   
  wire [5-1:0] f7crsrzernrwgmepy;   

  wire [64-1:0] vwxjizbv8c62_r6sf;
  wire [64-1:0] ft8qpl2cvbar7ci;
  wire [64-1:0] fi80hkldjwlh4v;

  wire [64-1:0] j7em0nbya;
  wire [64-1:0] ofkuwn9yg;

  wire                           rclkn1q60a3cbgtn67g ;
  wire [48-1:0] zamt9z8_hsjwlky8aktxv6;  
  wire [64-1:0]          ofmr0b7vez483r8wl ;
  wire [64-1:0]          zgn_d2n28xfn1zff ;
  wire [64-1:0]          ceewyf1unn6p7peejem ;
  wire [64-1:0]          oegl6jlhw01xkqeetu5y ;




  re1ncz9e2e3zo oiptvueshb9o(
    

    .k9lv9ppimt14qx3d7rj    (k9lv9ppimt14qx3d7rj  ),  
    .llskuqv0ehm60atlo     (llskuqv0ehm60atlo   ),
    .oug11blpzcta8zyu0ya   (oug11blpzcta8zyu0ya ),
    .zr1pc8tfxyljdj7a8a3eh5   (zr1pc8tfxyljdj7a8a3eh5 ),
    .qg9g70jgx5r5l_wpc7   (qg9g70jgx5r5l_wpc7 ),
    .o_qquv0pnx4zpz4h3gwxgl3  (o_qquv0pnx4zpz4h3gwxgl3),
    .j1fek3jzmt5bhhpnhvrmgt  (j1fek3jzmt5bhhpnhvrmgt),
    .ds75nafgmrespy002qvcsb8  (ds75nafgmrespy002qvcsb8),

    .rclkn1q60a3cbgtn67g     (rclkn1q60a3cbgtn67g  ) ,
    .zamt9z8_hsjwlky8aktxv6   (zamt9z8_hsjwlky8aktxv6),
    .ofmr0b7vez483r8wl    (ofmr0b7vez483r8wl ),
    .zgn_d2n28xfn1zff    (zgn_d2n28xfn1zff ),
    .ceewyf1unn6p7peejem    (ceewyf1unn6p7peejem ),
    .oegl6jlhw01xkqeetu5y    (oegl6jlhw01xkqeetu5y ),


    .ehq614orwiy4ww5(jc4yg1pkylr2gonwcd),
    .hgg2w2ca4wsixuj(nd3cgvec1pogf2),
    .lgv405vv46(f7crsrzernrwgmepy),

    .vwxjizbv8c62_r6sf(vwxjizbv8c62_r6sf),
    .ft8qpl2cvbar7ci(ft8qpl2cvbar7ci),
    .fi80hkldjwlh4v(fi80hkldjwlh4v),

    
    
    



    .dkmuhc79d2wm0wubp   (dkmuhc79d2wm0wubp ),
    .u2demhkod_er3kf6b (u2demhkod_er3kf6b ),
    .uz7pt71lvqit85od (uz7pt71lvqit85od ),
    .v3uvhtx7e5vbtvie  (v3uvhtx7e5vbtvie  ),
    .tmqkgmlzi018        (tmqkgmlzi018       ),
    .lx_olubu7t8h        (lx_olubu7t8h       ),
    .dd1p3tnenmm9r        (dd1p3tnenmm9r       ),
    .l60zv02z95hlayri      (l60zv02z95hlayri     ),
    .l1xzyldaa9dr2q7mla      (l1xzyldaa9dr2q7mla     ),
    .a5z_23_ryr_m29hhia_p (a5z_23_ryr_m29hhia_p),
                                        
    .vejdvgqormu727s  (vejdvgqormu727s  ),
    .ar9ro1ql86jzmq_p (ar9ro1ql86jzmq_p ),
    .qz1gqv6vh5qturw6v1mz(qz1gqv6vh5qturw6v1mz),

    .y7rd1k0an54clel_5q6   (y7rd1k0an54clel_5q6), 
    .com03bquiktu249yb0   (com03bquiktu249yb0), 
    .tzg0yjgx9bn98i    (tzg0yjgx9bn98i ),
    .x8_a2j7z3gz3l0tfjqp   (x8_a2j7z3gz3l0tfjqp),
    .c2mipfm_6z5ef4p3aoz    (c2mipfm_6z5ef4p3aoz ),
    .y3z8rf7c6hvsiux     (y3z8rf7c6hvsiux  ), 
 
    .xq0mj5mg2_512eu4   (xq0mj5mg2_512eu4), 
    .e11m1298jo38qcwq9er2   (e11m1298jo38qcwq9er2), 
    .ec94_mk193di7tj    (ec94_mk193di7tj ),
    .nodrapn01yl1vxle30p   (nodrapn01yl1vxle30p),
    .m2sw40fca0wvnmy    (m2sw40fca0wvnmy ),
    .ywhfwlbfro2dmuvf     (ywhfwlbfro2dmuvf  ), 

    .ex_g_cnadtiu1r9u   (ex_g_cnadtiu1r9u),
    .orzasugx5h5pio22_   (orzasugx5h5pio22_),
    .dxwtzud_wfj8jqk0    (dxwtzud_wfj8jqk0 ),
    .dn074lh73rzchvrqzm8   (dn074lh73rzchvrqzm8),
    .gi8o690aydhqi8    (gi8o690aydhqi8 ),
    .zl1r9cfvuhltjq     (zl1r9cfvuhltjq  ),
                      
    .xsn02pxoid_pw25   (j7em0nbya),
    .llv_dny70d   (ofkuwn9yg),



    .gc4b3kdcan6do88ta_        (gc4b3kdcan6do88ta_),
    .j4xe_w_yjq2       (j4xe_w_yjq2),
    .aui65oshqn8b5_iz6   (aui65oshqn8b5_iz6),
    .jmoafuo8zb_i1t   (jmoafuo8zb_i1t),
    .sa5of37yr6xn0s3e   (sa5of37yr6xn0s3e),
    .o_dsdljul          (o_dsdljul   ),
    .juyzxopct4k03sl      (juyzxopct4k03sl),
    .qyqw_37_fxv8z      (qyqw_37_fxv8z),
    .hyw0m71z3q3rpt1      (hyw0m71z3q3rpt1),
    
    .o5q5hev          (o5q5hev   ),
    .fx_h7chccf02z       (fx_h7chccf02z   ),
    .ru_wi            (ru_wi  ) 
  );


  wire                         f0jwv0n5olimpf4vnvqpb4hs;
  wire                         k8qtud5yr1e98g; 
  wire                         mw1zdgavbul7ic; 
  wire [64-1:0]        covjtr51ggzngufqow;
  wire [4 -1:0] qfhwjs9ygxr4e0rg86a;
  wire                         r86mhhg0562g6n9sah0z ; 
  wire                         aqz_nh46x0w0rdwc83s7c ; 
  wire                         oor8acg0u_d09e0moah ; 
  wire                         drgmlg58l2czwg2ijhc;
  wire                         hvgjjhizbfp9km9dd;
  wire [64 -1:0]  nd1hj8zlmdgys5obof18pe;
  wire [64 -1:0]  oe3uwa3e_ggymrc7ri;
  wire [4:0]                   a51im30isjous61asad1lrg5;

  wire                         z5vf_v21veoi10ybi; 
  wire [64-1:0]        tq4dt8fbx7xch3x4b;
  wire [4 -1:0] ip_8jolx6gnp;

  wire                         kzfv878bfk6iooqik; 
  wire                         o3cx5caf3g3nzd0pu; 
  wire [64-1:0]        woxzhk095h66amt5;
  wire [4 -1:0] n4bind2sncm8mh;
  wire                         wtw3apxzccvxdx8 ; 
  wire                         qfx1o1rp7psuvaq ; 
  wire                         zckohvd58ff_pyuth ; 
  wire                         j11k71dn8a;
  wire                         fov_crsecs;
  wire [64 -1:0]  avaoxa8z58nyr0g127g;
  wire [64 -1:0]  yc8cklg0l;
  wire [4:0]                   mb94n_xsixgup9p0;
  wire                         b0ylmw5xa8oytsw3j6n;










  wire                         flcopog5zzpohfautwy; 
  wire                         gtb8f_h0g28itdr8k; 
  wire                         wf15djwi2hw25nz_  ; 
  wire                         t1q5qmk9jzpf6glng4y;
  wire [64-1:0]        xsmx4zoewhbt07jxq;

  wire                         f5jobxqu5r8tdcgp9dz_; 
  wire                         hfh_n8b2_6ltn5lve4_271m; 
  wire                         xiy2xcok2j1vz3hdn21fq8us4e; 
  wire [32-1:0]   ezq9pnmedz815gxhjrvk5x; 
  wire                         k250aa9_7n16_xye3p__d4ew7; 
  wire                         p4_cbhjumvsd2_nee5pbvt1; 
  wire                         m63kr3yu_6uz_m3_yti5_e9; 
  wire                         rykqnjd3sew6zqm077moncthemet9; 
  wire                         z2oi9osh3p0wy7vb2sr69u07; 
  wire                         n1ko5ud3mahcu4f2t8; 
  wire                         gs8s9g8gtij6u619m3tcdcvnd;   
  wire                         i36cd1y8_65k09dz0thns;   
  wire                         wb6ynztvqw_c7jt0r60z0a3;   

  wire [64-1:0]        at3xavrqfa9vpvz2wfl28m2; 
  wire [8-1:0]     zawrb3vcmuri8b2986t8n2f; 
  wire [1:0]                   y_nw0z1jiz_z1j47b284ciw;
  wire                         sxokdo7nllqwvltwlem22uf5;
  wire [4 -1:0] z_l3eykrjali3v1mh46uf5mt;
  wire                         jis_avsh9dp0zny0zshz7;
  wire [4:0]                   tudsip00rgu_1pit8jhrmcjt35cbx; 

  wire  z_rab_1o8tf_6vir    ;
  wire  p9or1fzh0lqhmmmlo  ;
  wire  hj050gyk784wqb85v  ;


  wire                           y5qvboneeuu7u9c6ex2k32;
  wire                           r0b984qp4dbimt7m049jn;
  wire [4-1:0]       eq0u1926xaldb_6z8t8xdam;

  wire                           o4tmdwuwe0a_icm5c4xc3pnm0;
  wire                           vhfqvbg0i9tkhk8b7_1xw94s_n3h;
  wire [4-1:0]       hn6ha7kpsoxids4i7ilrw;
  wire [64-1:0]          qelk6ys1izwqop2178az43;

  wire                           wt6jy410rpokxn04lscbst6uo7;
  wire                           pdl18ljotymfj543wtjh49b_r;

  wire [4-1:0]       kavx5xx6zd8f9hqjq1s;
  wire [64-1:0]          z8hscmi55sjt_ufebya9e;

  wire                         o21b8ypt1xiu5ml63d; 
  wire                         badsf4ksbp3k6p_p5hnj2i; 
  wire                         vrsqde4muadsevgpemk; 
  wire                         ed4kcy8s9nrisftgx_q; 
  wire [32-1:0]   bdqo1tgw2_bpi2e8alini; 
  wire                         zdpamqgv7ddf1n3x5t2q; 
  wire                         wpsukhyqhl92dzoam7cm; 
  wire                         v3oo69y614hgiemyyld; 
  wire                         p648zxn2luyxy8mt992a; 
  wire                         uxlldm0w_h7kicit8gvhqv2; 
  wire                         yvu98r_7ji4o250r_u; 
  wire                         jp5nha2l14e7kx2jzpke;   
  wire                         za9xg3zsqni_aeqmke;   
  wire                         c1gmncmorg16sachdas;   
  wire [64-1:0]        a4a48egkdkec8d9b_9; 
  wire [8-1:0]     xwfmltfzahuj4qfn4qf2; 
  wire [1:0]                   ggxoqcj7ytp1a4pjf7ee;
  wire                         l3c127qdc9a2mfc13;
  wire [4 -1:0] oq9b5zfhza9yvdoj;
  wire                         sg33s7pt45jp_;
  wire                         g9i9mf8jq7sc699j;
  wire [4:0]                   szrgf24or2mbt7w_yleh_vt; 


  wire  yixt0a_xmh   ;
  wire  bp9qt1h52k23  ;
  wire  t6ehcvrshdj  ;
  wire  rm1dxjejhq7dh3q5m;
  wire  rvr30vvllni;


  wire n3zlo14nquu5l7zf3;

  wire a_1o1o8345o28hui ;
  wire t8p1kh0tvb2ej56s  ;
  wire                   p7ah58va5_2njbtv; 
  wire [64-1:0]  u981qrwkgi5h0e72b__gg19w;  
  wire                   p0i2i3v3j1tclelx51;
  
  
  
  
  
  
  
  

  
  
  



  wire r5hpbriny8m67sv9e_ylgo1;


  pxp_0xj1  u_ux607_exu(

    .ollg7               (ollg7),
    .d3n7pwgwcgze9cr4  (d3n7pwgwcgze9cr4),
    .amc4c8vcbecv1i     (amc4c8vcbecv1i   ),  
    .pby60vfdze02     (pby60vfdze02),
    .vm3pyzc9nt95     (vm3pyzc9nt95),
    .rbz4pv_atxqopdwt     (rbz4pv_atxqopdwt),
    .qs1xgat7r8xow     (qs1xgat7r8xow),


    .av1w8ld09cfofn     (av1w8ld09cfofn    ),
    .im2b5l0h98avl6t4sj (im2b5l0h98avl6t4sj),
    .bw65wl7fvekfymd8vqx  (bw65wl7fvekfymd8vqx ),
    .pecbpcoa04vq      (pecbpcoa04vq     ),
    .tb_snaxyfs       (tb_snaxyfs      ),
    .zc4mldgm25r      (zc4mldgm25r     ),
    .d23wb5yh1iyvf      (d23wb5yh1iyvf     ),
    .srim3bfnzhve       (srim3bfnzhve      ),
    .cy3nuhzm_v2p73mt  (cy3nuhzm_v2p73mt ),
    .fvqwdz2hdbb      (fvqwdz2hdbb     ),

     .a02zzbowpjn06h (a02zzbowpjn06h),
	.st4f16aums5        (st4f16aums5       ), 
	.p05ld2ghmwh        (p05ld2ghmwh       ), 

    .s7eq8f6z1uyi2in   (s7eq8f6z1uyi2in),
    .qbsr1jytrqtsbk4ttb8nz(qbsr1jytrqtsbk4ttb8nz),

    .w92a5o09fp9dg6   (w92a5o09fp9dg6   ),
    .eglor15f7p2ivpny5dc   (eglor15f7p2ivpny5dc   ),
    .ous_emkpecrqhg5e7(ous_emkpecrqhg5e7),
    .doh50j3p7c7yl7uk9(doh50j3p7c7yl7uk9),
    .wd9dvepxj        (wd9dvepxj),  
    .rm1dxjejhq7dh3q5m    (rm1dxjejhq7dh3q5m),
    .rvr30vvllni      (rvr30vvllni  ),
    .aw82i964do          (aw82i964do),
    .y8_gkxsfle          (y8_gkxsfle),

      .pcr4upio7_tx37     (pcr4upio7_tx37   ), 
      .uzklqlncpqqm1rav  (uzklqlncpqqm1rav),
      .ortueunvnkx_l5m_j  (ortueunvnkx_l5m_j),
      .hwuhtb7ucto_utk56  (hwuhtb7ucto_utk56),
      .i1env2kmns7qvvuuc  (i1env2kmns7qvvuuc),
      .g3s3vpafvy3i  (g3s3vpafvy3i),



      .uc5qxb4d2b28ye5          (uc5qxb4d2b28ye5),
      .o2qkf90r783          (o2qkf90r783),

      .habgbg2jn3qi     (habgbg2jn3qi),
      .dg4hzu_          (dg4hzu_     ),
      .h7fseh5_df0hbx     (h7fseh5_df0hbx),

    .bz8qao4o4xqslni1d3              (bz8qao4o4xqslni1d3                ),
    .vpecdc5kos                      (vpecdc5kos                        ), 
    .pccd7o463jfc_dpc5va               (pccd7o463jfc_dpc5va                 ), 
    .k5ovx8tintgvetip                    (k5ovx8tintgvetip                      ), 
    .f97le_hyejv7saw9vslna               (f97le_hyejv7saw9vslna                 ), 
    .yruel3nusosm39gnmb9ev_              (yruel3nusosm39gnmb9ev_                ), 
    .oeux55k_cre0he7w7jip5b1            (oeux55k_cre0he7w7jip5b1              ), 
    .r8z2r_ud53zj8mrpk               (r8z2r_ud53zj8mrpk                 ), 
    .bu1949pq_9946o1_e2q_uvr8p4         (bu1949pq_9946o1_e2q_uvr8p4           ), 
    .b4isf5u8b8pj34e09f72vxe38zg         (b4isf5u8b8pj34e09f72vxe38zg           ), 
    .kvpemhoim1tq5y8mzwvix5             (kvpemhoim1tq5y8mzwvix5               ), 
    .z1l_kkshyf_56cwmaq2dm           (z1l_kkshyf_56cwmaq2dm             ), 
    .w7u50np_chxy7wq5n9et_q           (w7u50np_chxy7wq5n9et_q             ), 
    .l2dse4sd3runnrb1rcbydauc            (l2dse4sd3runnrb1rcbydauc              ),  
    .kr1rhzlb5gr_wty1pe392s5oqet        (kr1rhzlb5gr_wty1pe392s5oqet          ), 
    .ox2ptuhum_e2aodz8wine6h         (ox2ptuhum_e2aodz8wine6h           ), 
    .g_qmxgznvfin609fmm97kuc2dm02         (g_qmxgznvfin609fmm97kuc2dm02           ), 
    .i9oln6xm1pi9dzsd61s1kg4dmo7j         (i9oln6xm1pi9dzsd61s1kg4dmo7j           ), 
    .hei_cs0rbwsv                    (hei_cs0rbwsv                      ), 
    .yf_5vs18cke5xg660my              (yf_5vs18cke5xg660my                ), 
    .deo3wn_907tw886r                 (sneofd4rq3b0m9eu91r8                   ),










    .dyl5g2vgrvy4mb3         (dyl5g2vgrvy4mb3         ),
    .r5hpbriny8m67sv9e_ylgo1   (r5hpbriny8m67sv9e_ylgo1         ),

    .umnrzb6pv8dzc (umnrzb6pv8dzc),


    .x8rpm78rvvycis(gvkx7hystgemle), 
    .h7lpiwlxyb79qyr06(ii7h_yx8mmn1y82k), 
    .canacnkc7zibtkn418i(f71s92bjwuhpisqhx13nk), 
    .bkkiffh6ob85nh79doya_(xrkn9p6pdpoya56pfoc6t), 
    .qhqqh0lyehgtfop1tc(qqo7mp2z_os7tj0c4w6kf6y), 
    

    .sxhicsqvufwfbnk0(mcfeo0u7nf9), 
    .c5wzn6bil69i9toc(sa3k3tsgxwqp8z), 
    .x03ux1utw4qem5kk3c(wfa5o72ctktgt55fgv2eo), 
    .pjic5x84bqxpvdduy4r2s(igeg6alwzopr62ti9), 
    .w5az87bw32r0tjbo0tdrv2ouvx(g3e0lri_3krzlfxnnlo_2y82qf),












    .enwn0u48p2_ls5az80          (enwn0u48p2_ls5az80),
    .f_i1959b4xizzq9jea     (f_i1959b4xizzq9jea),
    .b4lwcgm6l21pi          (b4lwcgm6l21pi),
    .hjrk_rwjkqj3zk_b         (hjrk_rwjkqj3zk_b),
    .zwcbp7zqfei5xz         (zwcbp7zqfei5xz),
    .znzjygllppv1s0a8cqub3c    (znzjygllppv1s0a8cqub3c), 
    .dxi_ue3gf5zqqqxwgq2a    (dxi_ue3gf5zqqqxwgq2a),
    .ix299qulxi5            (ix299qulxi5    ),
    .jjj61w03m77lv           (jjj61w03m77lv    ),
    .gfy3zost37aq8qmr          (gfy3zost37aq8qmr),
    .dz0zrf512290tvcy4q       (dz0zrf512290tvcy4q),
    .dn8riluj40uunvq5        (dn8riluj40uunvq5),
    .miax48k27o484e8a        (miax48k27o484e8a),
    .fzdb65fcrotwcaccus_cwo    (fzdb65fcrotwcaccus_cwo ),
    .tcy_87vt9vet39knuw     (tcy_87vt9vet39knuw  ),
    .fc_4ns_w1nh4h02z_dgg   (fc_4ns_w1nh4h02z_dgg),
    .jqsukc5b5drcc1e78       (jqsukc5b5drcc1e78    ),
    .gnn46rd7vvofruqij       (gnn46rd7vvofruqij    ),
    
    

    .qo5p9t6s74zxpo            (qo5p9t6s74zxpo),


    .gc4b3kdcan6do88ta_              (gc4b3kdcan6do88ta_),
    .tw5xnp59d8x               (tw5xnp59d8x),
    .um8zsjyxn_4p     (um8zsjyxn_4p   ),

    .emc_bywzarijbo             (emc_bywzarijbo),


    .v09gw6e6rfjf05qg           (v09gw6e6rfjf05qg),
    .fcjh1nct4r                (fcjh1nct4r),
    .x_cq40qmp6a            (x_cq40qmp6a),
    .z1l80uwh6vyyg34          (z1l80uwh6vyyg34),
    .rn1o3sl83              (rn1o3sl83),
    .zz5wo47gw146x4             (zz5wo47gw146x4),
    .fgr486jx5kevbua             (fgr486jx5kevbua),
    .pvfk1_6o89lmby              (pvfk1_6o89lmby),
    .xx87vzbpchg              (xx87vzbpchg),



    .k405wpjt       (mfnb4b0       ),   
    .epi4op2w5ban9o (edebnrit9_y77l ),   
    .heqeu11d07lcg2ss (gbhvs__f9z_q97jj ),   
    .exzr5we0sujvtby (hle5nop1tcht5cg ),   
    .anvecdxcx1ouoa0(t7panq_mivym6dhmjp),   
    .x240tjzbog6i9q(uaehep04469aadw4ga1),   
    .uimia9sdhaq9x(op60_2nivpji1_v8upx),   
    .bq9_5ksloh67_2ti(nzi6n_pc9q_5ybxyh),   
    .qosgyc25p4fzq8b4(sqliqgffeni4u6uzs),   
    .cqk3fh13g1cxf9j(gr8qapbswugbbkjl5),   





    .zscjnjl4ffiey84zel2    (k9lv9ppimt14qx3d7rj  ),  
    .qy0ycb_z4ngy2ll8pqo     (llskuqv0ehm60atlo   ),
    .nb2chelz4_ijwumv9murokla   (oug11blpzcta8zyu0ya ),
    .bcrcin74qehflgu36ch9ghyv   (zr1pc8tfxyljdj7a8a3eh5 ),
    .fbzipldpa3ewvv31mgr   (qg9g70jgx5r5l_wpc7 ),
    .nlptjpg_zybrljgsnky1iwvhf  (o_qquv0pnx4zpz4h3gwxgl3),
    .zgv8w7jqb5wr6l2elow5znmm  (j1fek3jzmt5bhhpnhvrmgt),
    .rpceina94e3bcz2ov7g1t_iom  (ds75nafgmrespy002qvcsb8),


    .c4i0yanuek7va0ztp     (rclkn1q60a3cbgtn67g  ) ,
    .ajk1fk4kecwsdaeiybv    (oegl6jlhw01xkqeetu5y ),
    .n5x33q1l9ewebt6692qaofd8   (zamt9z8_hsjwlky8aktxv6),  
    .eqhoch739wo4sqhno2u    (ofmr0b7vez483r8wl ),
    .qj1fn7kk041c_7kez4t2fkt    (zgn_d2n28xfn1zff ),
    .q2qa0la3s98x10a2aqsb73g    (ceewyf1unn6p7peejem ),


    .cjo14q6bim0c           (jc4yg1pkylr2gonwcd ),
    .yqawr6m8r98vjx73           (nd3cgvec1pogf2 ),
    .wuzzw7m7hpf4p6q31           (f7crsrzernrwgmepy ),

    .ndn228hd1n2x           (vwxjizbv8c62_r6sf),
    .kwk_z0jwwa2r           (ft8qpl2cvbar7ci),
    .fnbi_cp8jq6t9ropn           (fi80hkldjwlh4v),




    .er2ibckhm98h98(j7em0nbya),
    .tmi776v7orl(ofkuwn9yg),
    .uzevp4zrbs9gi (rnx27onf2lbe), 

    .dkmuhc79d2wm0wubp     (dkmuhc79d2wm0wubp ),
    .u2demhkod_er3kf6b   (u2demhkod_er3kf6b ),
    .uz7pt71lvqit85od   (uz7pt71lvqit85od ),
    .v3uvhtx7e5vbtvie    (v3uvhtx7e5vbtvie  ),
    .tmqkgmlzi018        (tmqkgmlzi018       ),
    .lx_olubu7t8h        (lx_olubu7t8h       ),
    .dd1p3tnenmm9r        (dd1p3tnenmm9r       ),
    .l60zv02z95hlayri      (l60zv02z95hlayri     ),
    .l1xzyldaa9dr2q7mla      (l1xzyldaa9dr2q7mla     ),
    .a5z_23_ryr_m29hhia_p (a5z_23_ryr_m29hhia_p),
                                        
    .vejdvgqormu727s  (vejdvgqormu727s  ),
    .ar9ro1ql86jzmq_p (ar9ro1ql86jzmq_p ),
    .qz1gqv6vh5qturw6v1mz(qz1gqv6vh5qturw6v1mz),
    .ptyuk4efbbdu9asp0b8cmreeh(j2t29hqv0s6c7),

    .y7rd1k0an54clel_5q6   (y7rd1k0an54clel_5q6), 
    .com03bquiktu249yb0   (com03bquiktu249yb0), 
    .tzg0yjgx9bn98i    (tzg0yjgx9bn98i ),
    .x8_a2j7z3gz3l0tfjqp   (x8_a2j7z3gz3l0tfjqp),
    .c2mipfm_6z5ef4p3aoz    (c2mipfm_6z5ef4p3aoz ),
    .y3z8rf7c6hvsiux     (y3z8rf7c6hvsiux  ), 
   
    .xq0mj5mg2_512eu4   (xq0mj5mg2_512eu4), 
    .e11m1298jo38qcwq9er2   (e11m1298jo38qcwq9er2), 
    .ec94_mk193di7tj    (ec94_mk193di7tj ),
    .nodrapn01yl1vxle30p   (nodrapn01yl1vxle30p),
    .m2sw40fca0wvnmy    (m2sw40fca0wvnmy ),
    .ywhfwlbfro2dmuvf     (ywhfwlbfro2dmuvf  ), 
                    
    .ex_g_cnadtiu1r9u   (ex_g_cnadtiu1r9u),
    .orzasugx5h5pio22_   (orzasugx5h5pio22_),
    .dxwtzud_wfj8jqk0    (dxwtzud_wfj8jqk0 ),
    .dn074lh73rzchvrqzm8   (dn074lh73rzchvrqzm8),
    .gi8o690aydhqi8    (gi8o690aydhqi8 ),
    .zl1r9cfvuhltjq     (zl1r9cfvuhltjq  ),
                      
    .f71k3zhdtjavw19c52g45  (e592323mqvany),


    .c5ewdqztjw9za                (c5ewdqztjw9za),
    .rn2mt6nngsc9w5cz        (rn2mt6nngsc9w5cz),

    .qeb3z0x5                (qeb3z0x5        ),
    .ibhfuwrztbm8p4gg            (ibhfuwrztbm8p4gg    ),
    .i8_5wt0vppx             (i8_5wt0vppx     ),
    .osv2437qj_3nuf         (osv2437qj_3nuf ),


    .b7g_vsn0zoewh6g1    (b7g_vsn0zoewh6g1),
    .onnv64ydiajl        (onnv64ydiajl    ),
    .r21i4by0bu3ks       (r21i4by0bu3ks   ),
    .hn85hkp2yav       (hn85hkp2yav),

    .j0qaxhuqtdi       (j0qaxhuqtdi     ),
    .pbzpk52jinfscit4mm     (pbzpk52jinfscit4mm   ),
    .gwj6ow6qvbhs0tc31     (gwj6ow6qvbhs0tc31   ),
    .iwdkm52x_w4hpak_a2_w  (iwdkm52x_w4hpak_a2_w),
    .mm0ssgy582fv_j       (mm0ssgy582fv_j     ),
    .ir2913p9xpmq_1bvfd1  (ir2913p9xpmq_1bvfd1),
    .bsjo0v5e0t556pph  (bsjo0v5e0t556pph),
    .mwegg_7inaca6povsw(mwegg_7inaca6povsw),
    .wnkp7091zrsevkbl  (wnkp7091zrsevkbl),


    .azll7rq5fab5ou      (azll7rq5fab5ou      ),
    .n6a0r_0zddzrme8      (n6a0r_0zddzrme8      ),
    .ns0i7siujgkrghjpqv6(ns0i7siujgkrghjpqv6),
                                     
    .pydatzxqqi               (pydatzxqqi  ),
    .t5trf35s8vy             (t5trf35s8vy),
    .zbac123pv78sbz3          (zbac123pv78sbz3),
    .z4e_m564fxae0kpbjr          (z4e_m564fxae0kpbjr),
    .zmwq3e9oijvo7d7          (zmwq3e9oijvo7d7),
    .hixy2y36a1pn0          (hixy2y36a1pn0),
    .ozwene1gdpatk6g             (ozwene1gdpatk6g   ),
    .sxvvsxtbhyvt             (sxvvsxtbhyvt   ),

    .c4ughu0qm5sfai           (c4ughu0qm5sfai),

    .jjzotrbn                (ifu_o_valid         ),
    .hw1_k1jmu                (ifu_o_ready         ),
    .j3oz8j2                   (ifu_o_ir            ),
    .bwjyqadn                   (ifu_o_pc        ),
    .u2k4dyp52s_m                (bcv5wwa3cpmh6o9d      ),
    .djvj1e_                (pbiupof7z_siv68x2      ),
    .bktu0z1mk56                (eey8q1ex7jqqx0hm_      ),
    .ipht6ss_sh6h               (hyzfgvg8iynh8zpa4        ),
    .piwiqvrjoq              (mdfkn7idoni9xj       ), 
    .al4xeg8mukgfg               (v3pirqtitn2_xu9        ), 
    .ryc6z1c7rmzrnlno           (n0p5652lvx0qj1yuwu    ), 
    .rhufxsnopy0n               (ddp4_khmuujfs        ), 
    .wbhvg_1r9435               (m_7gx91ep6vkla        ), 
    .s1woka0byzgo             (iyoccmh9a_a2ov94o      ), 
    .cpt0qfwiz               (s8mlhtj2pe58l        ),
    .vf7a_1kae4zv5               (eh7xldx93qn_e_ig        ),
    .djv9nstr               (mxxfa5sn2ahc21k        ),
    .gy5zhpbrnl                (wp3ochi2x8_ljvjh         ),
    .qv70a7n8p                (yzl1nx341x5d2p4         ),
    .anlbkc8jny                (l11qpt1sf6a7         ),
    .qhyq467foflgyn5y           (n3mz6a4lr36ftz11    ),
    .binjv97px9r7dt04h0          (f2d4k4kxynjpd0gghqe140   ),
    .jt4l0g4njcsrt720n         (uuy2zpbrzrwdf432a7_g  ),
    .w7uciar2_6p9xc5mc         (d4d7ru_yllps7en_tto  ),
    .m9cdnl05ykr_3p             (ylmhlw32ex4fxli7       ),
    .ex6ixmgf331             (n_lam8gs1mljgiq8zi       ),
    .akh3h7anvh7892ugn        (v_97hsna5xll5n1xslwe3),
    .vfu1cc_k9n55lt38g_vii       (v2r90qa11qssvr5tq98dbi961),  
    .o_d157fc5_l              (ba89afyz0al00        ),
    .texy7g6tpvcgwtyd           (gkonom22e0fpa2_v3w0ab     ),
    .oypxxr_e_rms7ai          (fxvpc9o9zl2t2nuwpg0    ),
    .gkps1gyqdwgzcvr0c          (gtvau5cygdmb10dr_makqf    ),
    .s68_9qhgnb_o              (xosc7587i2hjow2yjw        ),
    .q52oeddgdt76b              (p54semfzu2zyfb        ),
    .ajl4tppx98ihuirj_mxih      (qu31vl4s4x0pmeth2j_7neq1),
    .sa2f4h4xeakpfnunl           (himvp4q0erus0anat5    ),
    .nrebzehsuam                 (ps9l2wesoladg           ),

    .y_0q8d40rrzolo1y6       (y_0q8d40rrzolo1y6),
    .ao17frh5wnr0wddz3       (ao17frh5wnr0wddz3),
    .mmludd_fnt2yevok8a1a0       (mmludd_fnt2yevok8a1a0),
    .buwj9_8l8bwj80kkinq9p       (buwj9_8l8bwj80kkinq9p),

    .hwpkcsh2atrq            (hwpkcsh2atrq  ),
    .v3e6l1k7eo9k3           (v3e6l1k7eo9k3 ),
    .hxrmt706n071lic0f7          (hxrmt706n071lic0f7),
    .gfod0nmy6eta29jeeg6mr2     (tluzd_2baaw1fpd4o1td_h),
    .n4soswat5yihd74b        (agcvtek_6ocmw76d),
    .if0fog4bug_zkykpi         (j0_nonyh_r387uiy),
    .lln3b7iev7jpvogh964ro_9bc_3y  (lln3b7iev7jpvogh964ro_9bc_3y),
    .q97rqfy8n7ixfm2a5wev4nd5sylpcq3j (q97rqfy8n7ixfm2a5wev4nd5sylpcq3j),
    .hujgg6hjnhtbspbkekuz5_u        (hujgg6hjnhtbspbkekuz5_u),
    .v3pnt81kfrgbaanm1mhh51w         (v3pnt81kfrgbaanm1mhh51w),
    .i08eq60d_snxeq8si_ezod        (i08eq60d_snxeq8si_ezod),
    .y8wz7aud_fd6dfiakjtx2i0g  (y8wz7aud_fd6dfiakjtx2i0g),
    .dgnjyd9xs8efyxm0tdlsvfq4eop (dgnjyd9xs8efyxm0tdlsvfq4eop),
    .a3xib90kwk4_hm1        (a3xib90kwk4_hm1),
    .nfzexr8q9g893gi         (nfzexr8q9g893gi),
    .opkkwp3eg8g3448t        (opkkwp3eg8g3448t),
    .zsgl59ydqwjln         (zsgl59ydqwjln      ),
    .b9yq2alidby7zgom1         (b9yq2alidby7zgom1      ),


    .tvqijouldcgiz2dxdco7    (tvqijouldcgiz2dxdco7),
    .zkxlkidschdubxpkpm    (zkxlkidschdubxpkpm),
    .xmcrni1qngfvh9pil9j    (xmcrni1qngfvh9pil9j),
    .btkcf2uqr61gkiqhde0lai    (btkcf2uqr61gkiqhde0lai),
    .h01d94xsxbxe_req          (h01d94xsxbxe_req),  
    .w1casjl7bz73brz      (w1casjl7bz73brz),
    .hjri7cufo9ckntq      (hjri7cufo9ckntq),
    .yghffofulqa77bd7aw07badta1a  (yghffofulqa77bd7aw07badta1a  ),
    .rrl7evvmayt1_vvp74iq9h6_cjf(rrl7evvmayt1_vvp74iq9h6_cjf),
    .zddoxp22m1o11x30gbe      (zddoxp22m1o11x30gbe      ),
    .hwfethpzkuauejcgtbl6o    (hwfethpzkuauejcgtbl6o    ),  
    .n3ak8l6cvn0s4           (n3ak8l6cvn0s4     ),
    .hsxh9536ho4bw8o           (hsxh9536ho4bw8o     ),
    .r_edve7v9jcr26q6zk      (r_edve7v9jcr26q6zk),
    .vrqfzuog2k4pos133      (vrqfzuog2k4pos133),
    .bmw2yi333716crywk      (bmw2yi333716crywk),
    .k2sr7sw1plcmnki5ajtscw      (k2sr7sw1plcmnki5ajtscw),
    .jkzw_f9anx55            (jkzw_f9anx55      ),
    .t8muv9e6d7yk_whqa0        (t8muv9e6d7yk_whqa0),
    .hzdfp71n6g3f5fsg5        (hzdfp71n6g3f5fsg5),
    .lwdhmuzyvcvv14mjbl0h2a41z  (lwdhmuzyvcvv14mjbl0h2a41z  ),
    .xy48dugh009wtmazqug3kpy2a5h_(xy48dugh009wtmazqug3kpy2a5h_),
    .l4ztejmt2__wxqm2rw      (l4ztejmt2__wxqm2rw      ),
    .s3ujdp2a8n69bm6engxok    (s3ujdp2a8n69bm6engxok    ),  


    .vz63qkw5s3m8urb9        (z5vf_v21veoi10ybi ),
    .iojqlhtwx45_siz         (tq4dt8fbx7xch3x4b  ),
    .ydtm1yuxqj7fmxvqc         (ip_8jolx6gnp  ),

    .o4qff84vfbn            (kzfv878bfk6iooqik   ),
    .x74_jhmpouk            (o3cx5caf3g3nzd0pu   ),
    .z5tnbveujliw633sxlb8        (woxzhk095h66amt5    ),
    .l8ng5e_pa1fg07__37        (n4bind2sncm8mh    ),
    .erdoc9bbdnq8065yw         (wtw3apxzccvxdx8     ),
    .rqy9v1_k_o74etonfc       (zckohvd58ff_pyuth     ),
    .ro93aearv5754gz9w       (qfx1o1rp7psuvaq     ),
    .zqx1cj9lvt0e           (j11k71dn8a),
    .zsxgccndqw2suf6           (fov_crsecs),
    .y9389ymcyh2ia2082yx1_      (avaoxa8z58nyr0g127g     ),
    .uiu4_g7j41kz           (yc8cklg0l),
    .ytp8_jsqr2sjmu08gdn       (mb94n_xsixgup9p0),
    .b0ylmw5xa8oytsw3j6n      (b0ylmw5xa8oytsw3j6n),

    .f0jwv0n5olimpf4vnvqpb4hs  (f0jwv0n5olimpf4vnvqpb4hs),

    .flcopog5zzpohfautwy     (flcopog5zzpohfautwy ),
    .gtb8f_h0g28itdr8k     (gtb8f_h0g28itdr8k ),
    .wf15djwi2hw25nz_       (wf15djwi2hw25nz_   ),
    .t1q5qmk9jzpf6glng4y   (t1q5qmk9jzpf6glng4y),
    .xsmx4zoewhbt07jxq     (xsmx4zoewhbt07jxq),
    .xmbe_e4vm6ofjbn7lq        (xmbe_e4vm6ofjbn7lq),

    .o21b8ypt1xiu5ml63d        (f5jobxqu5r8tdcgp9dz_     ),

    .yixt0a_xmh               (z_rab_1o8tf_6vir  ), 
    .ej7frm_ut9j6y           (p9or1fzh0lqhmmmlo), 
    .izjeme5aukvcc           (hj050gyk784wqb85v), 

    .badsf4ksbp3k6p_p5hnj2i      (hfh_n8b2_6ltn5lve4_271m   ),
    .ed4kcy8s9nrisftgx_q      (xiy2xcok2j1vz3hdn21fq8us4e   ),
    .bdqo1tgw2_bpi2e8alini       (ezq9pnmedz815gxhjrvk5x    ),
    .zdpamqgv7ddf1n3x5t2q      (k250aa9_7n16_xye3p__d4ew7   ),
    .wpsukhyqhl92dzoam7cm      (p4_cbhjumvsd2_nee5pbvt1   ),
    .v3oo69y614hgiemyyld      (m63kr3yu_6uz_m3_yti5_e9   ),
    .p648zxn2luyxy8mt992a   (rykqnjd3sew6zqm077moncthemet9 ),
    .uxlldm0w_h7kicit8gvhqv2     (z2oi9osh3p0wy7vb2sr69u07 ),
    .yvu98r_7ji4o250r_u         (n1ko5ud3mahcu4f2t8),
    .jp5nha2l14e7kx2jzpke       (gs8s9g8gtij6u619m3tcdcvnd    ),
    .za9xg3zsqni_aeqmke       (i36cd1y8_65k09dz0thns    ),
    .c1gmncmorg16sachdas       (wb6ynztvqw_c7jt0r60z0a3    ),
    .a4a48egkdkec8d9b_9      (at3xavrqfa9vpvz2wfl28m2   ),
    .xwfmltfzahuj4qfn4qf2      (zawrb3vcmuri8b2986t8n2f   ),
    .ggxoqcj7ytp1a4pjf7ee       (y_nw0z1jiz_z1j47b284ciw    ),
    .l3c127qdc9a2mfc13      (sxokdo7nllqwvltwlem22uf5   ),
    .oq9b5zfhza9yvdoj       (z_l3eykrjali3v1mh46uf5mt    ),
    .sg33s7pt45jp_           (jis_avsh9dp0zny0zshz7        ),
    .szrgf24or2mbt7w_yleh_vt (tudsip00rgu_1pit8jhrmcjt35cbx), 


    .p1kjflyurzeuxj      (y5qvboneeuu7u9c6ex2k32),
    .yvjlu1e9eng5_5tme     (r0b984qp4dbimt7m049jn),
    .hh8nc68zrpki2m9r    (eq0u1926xaldb_6z8t8xdam),
    .v8wv99vga5gkl8xhk7x9in  (o4tmdwuwe0a_icm5c4xc3pnm0),
    .ahfx5rs9jkdyw3b8ztscfx (vhfqvbg0i9tkhk8b7_1xw94s_n3h),
    .ts3_k4ergzh8upz7     (hn6ha7kpsoxids4i7ilrw),
    .ktqya1x1mfi5j3q7      (qelk6ys1izwqop2178az43),
    .z6njhanl_m_hv48x5i9y  (wt6jy410rpokxn04lscbst6uo7),
    .dvm_h24fnflt11prmyvme (pdl18ljotymfj543wtjh49b_r),
    .uvyubcp0tbk9yirhz     (kavx5xx6zd8f9hqjq1s),
    .ivoui15mvw3de5ds44      (z8hscmi55sjt_ufebya9e),

    .n3zlo14nquu5l7zf3   (n3zlo14nquu5l7zf3),

    .a_1o1o8345o28hui      (a_1o1o8345o28hui),
    .t8p1kh0tvb2ej56s    (t8p1kh0tvb2ej56s ),
    .p7ah58va5_2njbtv     (p7ah58va5_2njbtv     ),
    .u981qrwkgi5h0e72b__gg19w(u981qrwkgi5h0e72b__gg19w),
    .p0i2i3v3j1tclelx51    (p0i2i3v3j1tclelx51    ),
    
    
    
    
    
    
    
    
    
    
    
    


    .um28jgd2x4mbs             (um28jgd2x4mbs    ),
    .l_imk5zs8ejjka              (l_imk5zs8ejjka     ),
    .lz3vnoxnz_z             (lz3vnoxnz_z    ),
    .yhbtmo4kyz_ewog3           (yhbtmo4kyz_ewog3  ),
    .cd4d2_i3rcc1_p          (cd4d2_i3rcc1_p ),
    .wyu42gj62n994v0wo_          (wyu42gj62n994v0wo_ ),
    .x9cmkt53yq483z1         (x9cmkt53yq483z1),
    .cxmwxfttqy2t7ura            (cxmwxfttqy2t7ura   ),
    .b5wruck8tj9sa            (b5wruck8tj9sa   ),
    .bxentpryfwb3d           (bxentpryfwb3d  ),
    .o2a43mjdbgea1           (o2a43mjdbgea1  ),


    .ij_sgq3rtvw2                (ij_sgq3rtvw2),
    .k9jntnqwqp               (k9jntnqwqp),

    .dk2xhkj77a                (dk2xhkj77a),
    .gf33atgy                    (c8fchlpwl),
    .stlp3kak                 (erv7j3wmd3gb_dp),
    .ru_wi                  (ru_wi  ) 
  );

  assign sfyn3seo6gs = ifu_o_valid;
  assign sgthjbo1oq1kw1e6 = ifu_o_ready;

  wire                        cv0k9k_ijjnnylw1s7b_0d;

  wire                        swpk4h0gei3t_34xogbqncbo4;

  wire                        u9qmfl3rwx0dhr92z875vx7q;
  wire [32-1:0]  unu_x_i6jmr33nz0yitzk; 
  wire                        bei3qhdtd0euq2emblogsu_x; 
  wire [64-1:0]       bf0_ynb648lqi7s93eieo0ln;
  wire [8-1:0]    wf8o7p9_qfthhoxs747wyeuwkky;
  wire [2:0]                  ygro7xue7x7rtdafkj3o4q4;
  wire [1:0]                  drrly3q0ocg8d4pwh3m9o77;
  wire                        g654a6a9cesbee7xs6_uu9lu5;
  wire                        x7fex0jf9da6a5v1c28upl72t;
  wire [1:0]                  ege0_1ufqm8i68zo4il6cwe46d;
  wire                        ngyxf4n1cpcgks_s2zmgfb260;
  wire                        c7m50uaw8lmp_iv4ci38q2;
  wire                        m04a1mtbabwezldp1crh4rg6z;
  wire                        hwjq1ubtaei44lpk609fm2hb8;
  wire                        e28p_fu1k484ncul0p85ko;

  wire                        bvg_3t_ujbpur7b_h7f63jse;

  wire                        m5l6wu3uz_jfqasz8e3tsvrm;
  wire                        g9so28ythfl0q7xnk66p1  ;
  wire                        e66wluxk71p2ldu3a1qk994bq  ;
  wire [64-1:0]       ig2roj0y08x8_ntp3knz9rd;

  wire                        a0_d_zdz9h9fgk46e8arf;

  wire                        twr9y24wxhs3qj2z9f2hzpaig6;

  wire                        w8b46r9cof57xvd5zo1u4zh8;
  wire [32-1:0]  wn1l4cmih7rwce1rb7wk3f9wy; 
  wire                        cgnzbuo_1yz6v42seb25duv; 
  wire [64-1:0]       zopev7f487spn9mwvuowqo;
  wire [8-1:0]    p32jk0lb8g31kqlpvmllo75qim;
  wire [2:0]                  g973rcaou05i456suvk_89dm;
  wire [1:0]                  wflv6rhfdwyxttak111v1l;
  wire                        ggsmt4nzx8pwlowehinqvk60f;
  wire                        xu8494ii8ectqb91224uuer;
  wire [1:0]                  r6rk128ijo839ougen9stbe;
  wire                        xo6ciibewn8p8xey97jcsqi5;
  wire                        evz1w_girwszyfnlcg4mwvtjo;
  wire                        ju5f9fb1erjep_bv8gpfn6;
  wire                        hadi1_f3quoaotjv5758x8kksot2;
  wire                        bdi4gjlb0po4ejcztowoqil7;

  wire                        m7tq_t57mr5bovbb9ghffl4k;

  wire                        gpcgdcri3e6_fxrw8wwtysoqqr;
  wire                        a6s4kxg1ibr6mntc85jik  ;
  wire                        hizzalmpwr8cqkxqi80wvbt65x  ;




  wire                        g1jacxqkf1oj5l4jvp9a7qacc3;
  wire                        nj35btypmlzn6n67k5a3sbxlz_;
  wire [32-1:0]   vknrn2pdsorktjh1khqd1o5u; 
  wire                        otv_22s88_efzve7t9aewczn; 
  wire [32-1:0]        huhgp41uzpgntu1igqiuh8bpy;
  wire [4-1:0]      glmsykv9_w4rhlqnh8qmvqcu3n;
  wire                        y69op1rhrojqmwt2zvwvt6_w1v;
  wire                        qya9tage13i6s6ij4c93w406f;
  wire [1:0]                  kbs9xq0ed1rv9h4kn8c9l7v8_c;
  wire                        kul32yktlkh84fqkeuiasdj4c;
  wire                        a0711e1j5ewmq9032iiam6zd;
  wire                        yxxau7egbjhe86w26b64yf;
  wire                        u4pdpnruu01ssoo78t_r;
  wire                        wpa_w8k78vc5tscpvglay54t;
  wire                        j_xo5pr2yvkxhr8c7fcp5m;
  wire                        o7cx0ajdhtouycxdeb8ly50;
  wire                        xjpj_prxqbclz5urycgi1vv;
  
  
  wire                        n71nv9q2skeheb436zhxyw8iy;
  wire                        ah736xwkrzyalnwp8ow6mi1z;
  wire                        pn6t3ogf6fkiu3lq50zejhq2_  ;
  wire                        nyapu28mzy38j3qnbv84wn19w;
  wire [32-1:0]        lfg1njvjoj4o9aupkvjol5f;


  neplroszbk3r28 gdqagtg556cxpg(

    .f5jobxqu5r8tdcgp9dz_     (f5jobxqu5r8tdcgp9dz_     ),
    .hfh_n8b2_6ltn5lve4_271m   (hfh_n8b2_6ltn5lve4_271m ),
    .xiy2xcok2j1vz3hdn21fq8us4e   (xiy2xcok2j1vz3hdn21fq8us4e ),
    .ezq9pnmedz815gxhjrvk5x    (ezq9pnmedz815gxhjrvk5x  ),
    .k250aa9_7n16_xye3p__d4ew7   (k250aa9_7n16_xye3p__d4ew7 ),
    .p4_cbhjumvsd2_nee5pbvt1   (p4_cbhjumvsd2_nee5pbvt1 ),
    .m63kr3yu_6uz_m3_yti5_e9   (m63kr3yu_6uz_m3_yti5_e9 ),
    .rykqnjd3sew6zqm077moncthemet9 (rykqnjd3sew6zqm077moncthemet9 ),
    .z2oi9osh3p0wy7vb2sr69u07  (z2oi9osh3p0wy7vb2sr69u07 ),
    .n1ko5ud3mahcu4f2t8      (n1ko5ud3mahcu4f2t8),
    .gs8s9g8gtij6u619m3tcdcvnd    (gs8s9g8gtij6u619m3tcdcvnd  ),
    .i36cd1y8_65k09dz0thns    (i36cd1y8_65k09dz0thns  ),
    .wb6ynztvqw_c7jt0r60z0a3    (wb6ynztvqw_c7jt0r60z0a3  ),
    .at3xavrqfa9vpvz2wfl28m2   (at3xavrqfa9vpvz2wfl28m2 ),
    .zawrb3vcmuri8b2986t8n2f   (zawrb3vcmuri8b2986t8n2f ),
    .y_nw0z1jiz_z1j47b284ciw    (y_nw0z1jiz_z1j47b284ciw  ),

    .sxokdo7nllqwvltwlem22uf5   (sxokdo7nllqwvltwlem22uf5),
    .z_l3eykrjali3v1mh46uf5mt    (z_l3eykrjali3v1mh46uf5mt),
    .jis_avsh9dp0zny0zshz7        (jis_avsh9dp0zny0zshz7),


    .tudsip00rgu_1pit8jhrmcjt35cbx(tudsip00rgu_1pit8jhrmcjt35cbx), 

    .z_rab_1o8tf_6vir            (z_rab_1o8tf_6vir          ),  
    .as_mlum8anvtnrny9tls        (p9or1fzh0lqhmmmlo        ), 
    .fd8f2gq4oaalsv4p_j        (hj050gyk784wqb85v        ), 


  .y5qvboneeuu7u9c6ex2k32 (y5qvboneeuu7u9c6ex2k32),
  .r0b984qp4dbimt7m049jn (r0b984qp4dbimt7m049jn),
  .eq0u1926xaldb_6z8t8xdam (eq0u1926xaldb_6z8t8xdam),
  .o4tmdwuwe0a_icm5c4xc3pnm0 (o4tmdwuwe0a_icm5c4xc3pnm0),
  .vhfqvbg0i9tkhk8b7_1xw94s_n3h (vhfqvbg0i9tkhk8b7_1xw94s_n3h),
  .hn6ha7kpsoxids4i7ilrw (hn6ha7kpsoxids4i7ilrw),
  .qelk6ys1izwqop2178az43 (qelk6ys1izwqop2178az43),
  .wt6jy410rpokxn04lscbst6uo7 (wt6jy410rpokxn04lscbst6uo7),
  .pdl18ljotymfj543wtjh49b_r (pdl18ljotymfj543wtjh49b_r),
  .kavx5xx6zd8f9hqjq1s (kavx5xx6zd8f9hqjq1s),
  .z8hscmi55sjt_ufebya9e (z8hscmi55sjt_ufebya9e),



  .slk31s106jz  (n3zlo14nquu5l7zf3),

    .yixt0a_xmh            (yixt0a_xmh          ), 
    .fgnb7mhn1254le9        (bp9qt1h52k23        ), 
    .okt7c24tca9ji6pw        (t6ehcvrshdj        ), 
    .o21b8ypt1xiu5ml63d        (o21b8ypt1xiu5ml63d     ),

    .badsf4ksbp3k6p_p5hnj2i   (badsf4ksbp3k6p_p5hnj2i ),
    .vrsqde4muadsevgpemk   (vrsqde4muadsevgpemk ),
    .ed4kcy8s9nrisftgx_q   (ed4kcy8s9nrisftgx_q ),
    .bdqo1tgw2_bpi2e8alini    (bdqo1tgw2_bpi2e8alini  ),
    .zdpamqgv7ddf1n3x5t2q   (zdpamqgv7ddf1n3x5t2q ),
    .wpsukhyqhl92dzoam7cm   (wpsukhyqhl92dzoam7cm ),
    .v3oo69y614hgiemyyld   (v3oo69y614hgiemyyld ),
    .p648zxn2luyxy8mt992a (p648zxn2luyxy8mt992a ),
    .uxlldm0w_h7kicit8gvhqv2  (uxlldm0w_h7kicit8gvhqv2 ),
    .yvu98r_7ji4o250r_u      (yvu98r_7ji4o250r_u),
    .jp5nha2l14e7kx2jzpke    (jp5nha2l14e7kx2jzpke  ),
    .za9xg3zsqni_aeqmke    (za9xg3zsqni_aeqmke  ),
    .c1gmncmorg16sachdas    (c1gmncmorg16sachdas  ),
    .a4a48egkdkec8d9b_9   (a4a48egkdkec8d9b_9 ),
    .xwfmltfzahuj4qfn4qf2   (xwfmltfzahuj4qfn4qf2 ),
    .ggxoqcj7ytp1a4pjf7ee    (ggxoqcj7ytp1a4pjf7ee  ),

    .l3c127qdc9a2mfc13   (l3c127qdc9a2mfc13),
    .oq9b5zfhza9yvdoj    (oq9b5zfhza9yvdoj),
    .sg33s7pt45jp_        (sg33s7pt45jp_),
    .g9i9mf8jq7sc699j           (g9i9mf8jq7sc699j        ),


    .szrgf24or2mbt7w_yleh_vt(szrgf24or2mbt7w_yleh_vt), 

  .f0jwv0n5olimpf4vnvqpb4hs (f0jwv0n5olimpf4vnvqpb4hs),

  .gf33atgy   (c8fchlpwl),
  .ru_wi (ru_wi) 
  );

  dkh50cge16y  irl6exrcvz(
  .rm1dxjejhq7dh3q5m(rm1dxjejhq7dh3q5m),
  .sxvvsxtbhyvt  (sxvvsxtbhyvt),

  .pcr4upio7_tx37   (pcr4upio7_tx37   ), 
  .uzklqlncpqqm1rav(uzklqlncpqqm1rav),
  .ortueunvnkx_l5m_j(ortueunvnkx_l5m_j),
  .hwuhtb7ucto_utk56(hwuhtb7ucto_utk56),
  .i1env2kmns7qvvuuc(i1env2kmns7qvvuuc),
  .g3s3vpafvy3i(g3s3vpafvy3i),
                            
  .rvr30vvllni  (rvr30vvllni  ),


    .dn8riluj40uunvq5       (dn8riluj40uunvq5),
    .w92a5o09fp9dg6        (w92a5o09fp9dg6), 
    .eglor15f7p2ivpny5dc        (eglor15f7p2ivpny5dc), 
    .qo5p9t6s74zxpo         (qo5p9t6s74zxpo),


    .umnrzb6pv8dzc          (umnrzb6pv8dzc),
    .o4qff84vfbn         (k8qtud5yr1e98g),
    .x74_jhmpouk         (mw1zdgavbul7ic),
    .z5tnbveujliw633sxlb8     (covjtr51ggzngufqow),
    .l8ng5e_pa1fg07__37     (qfhwjs9ygxr4e0rg86a),
    .erdoc9bbdnq8065yw      (r86mhhg0562g6n9sah0z ),
    .rqy9v1_k_o74etonfc    (oor8acg0u_d09e0moah),
    .ro93aearv5754gz9w    (aqz_nh46x0w0rdwc83s7c),
    .zqx1cj9lvt0e        (drgmlg58l2czwg2ijhc),
    .zsxgccndqw2suf6        (hvgjjhizbfp9km9dd),
    .y9389ymcyh2ia2082yx1_   (nd1hj8zlmdgys5obof18pe),
    .uiu4_g7j41kz        (oe3uwa3e_ggymrc7ri),
    .ytp8_jsqr2sjmu08gdn    (a51im30isjous61asad1lrg5),

    .flcopog5zzpohfautwy     (flcopog5zzpohfautwy ),
    .gtb8f_h0g28itdr8k     (gtb8f_h0g28itdr8k ),
    .wf15djwi2hw25nz_       (wf15djwi2hw25nz_   ),
    .t1q5qmk9jzpf6glng4y   (t1q5qmk9jzpf6glng4y),
    .xsmx4zoewhbt07jxq     (xsmx4zoewhbt07jxq),

    .yixt0a_xmh            (yixt0a_xmh          ), 
    .fgnb7mhn1254le9        (bp9qt1h52k23        ), 
    .okt7c24tca9ji6pw        (t6ehcvrshdj        ), 
    .o21b8ypt1xiu5ml63d        (o21b8ypt1xiu5ml63d     ),

    .badsf4ksbp3k6p_p5hnj2i   (badsf4ksbp3k6p_p5hnj2i ),
    .vrsqde4muadsevgpemk   (1'b0 ),
    .ed4kcy8s9nrisftgx_q   (ed4kcy8s9nrisftgx_q ),
    .bdqo1tgw2_bpi2e8alini    (bdqo1tgw2_bpi2e8alini  ),
    .zdpamqgv7ddf1n3x5t2q   (zdpamqgv7ddf1n3x5t2q ),
    .wpsukhyqhl92dzoam7cm   (wpsukhyqhl92dzoam7cm ),
    .v3oo69y614hgiemyyld   (v3oo69y614hgiemyyld ),
    .p648zxn2luyxy8mt992a (p648zxn2luyxy8mt992a ),
    .uxlldm0w_h7kicit8gvhqv2  (uxlldm0w_h7kicit8gvhqv2 ),
    .yvu98r_7ji4o250r_u      (yvu98r_7ji4o250r_u),
    .jp5nha2l14e7kx2jzpke    (jp5nha2l14e7kx2jzpke  ),
    .za9xg3zsqni_aeqmke    (c1gmncmorg16sachdas  ),
    .c1gmncmorg16sachdas    (za9xg3zsqni_aeqmke  ),
    .a4a48egkdkec8d9b_9   (a4a48egkdkec8d9b_9 ),
    .xwfmltfzahuj4qfn4qf2   (xwfmltfzahuj4qfn4qf2 ),
    .ggxoqcj7ytp1a4pjf7ee    (ggxoqcj7ytp1a4pjf7ee  ),

    .l3c127qdc9a2mfc13   (l3c127qdc9a2mfc13),
    .oq9b5zfhza9yvdoj    (oq9b5zfhza9yvdoj),
    .sg33s7pt45jp_        (sg33s7pt45jp_),
    .g9i9mf8jq7sc699j           (g9i9mf8jq7sc699j        ),


    .szrgf24or2mbt7w_yleh_vt(szrgf24or2mbt7w_yleh_vt), 


    .cxrbvs1hde7j8ziudd4ar          (xib8tki1lzl05e71ry   ), 
    .dmzxpdd5dgmp_2ip6h3_6          (hdle8ta5fimb1inf1z   ), 
    .piv1ndd8n8dlaqx9           (trtxm7l0l_kp36i9y    ),
    .dycy3iz66xw6yj5ea           (p0akg_4worvsnfq_q36vp    ),
    .zqnzorh6g9hnwsot5zr         (1'b0 ),  
	.sp2wnouu73ujsanhkn0           (1'b0 ),
	.n5w05rcecv47nvnfkkw5           (1'b0 ),
	.r3rgwuaokuw68zin           (1'b1 ),
	.p1g5jbgswdsx9v1j01103          (64'b0),
	.zmrmpw_9vyme3rakn8br8e          (8'b0),
    .fd_1f891ni339pnyzw63mg          (vl5p5iump0rpm1hbr   ),  
    .m2aue5rcrjkbzdwbqvlzvr          (oj6rvjf7ujgb34264   ),  
    .u7a8_cbg_zi4w4b4slc08          (vjfz03uzu8p_0jhhvvev   ),  
    .wic6t212ob4tfa             (mqdc73rtez0bzh2_1      ),  

    .ro76scx3ggmfi4xp2bjx          (p1qeemcgwrrzzt73bl   ),
    .t9yh0n7ay27ft001vimu6          (ertspxpg0txqgp9i6fx53   ),
    .gpjxeoxkmf35ldn            (z3xt8rx_qs6z0goo1     ),
	.owde01ai01h2x5kn3_ng        (),
    .atur2zwqwk4mnbtz68l2          (ln7r12q36ofpcd6m6u    ),


	.fkm9up63o1aeauaqhjb   (fkm9up63o1aeauaqhjb),
	.to_1lv9wnb3vmu6tvz5rc   (to_1lv9wnb3vmu6tvz5rc),
	.ju1kbeplcqy314lfj4    (ju1kbeplcqy314lfj4 ), 
	.r985fbe5k7hgzaq9i    (r985fbe5k7hgzaq9i ), 
	.bb04gpwotp2s6c7_p1gqkq   (bb04gpwotp2s6c7_p1gqkq), 
	.sqmey185cu3mtixhl   (sqmey185cu3mtixhl), 
	.rffcsd1o699ytclmx   (rffcsd1o699ytclmx),
	.lbr88vbqtg8rht7320frde   (lbr88vbqtg8rht7320frde),
	.g7qq38mx3d58n1b15kcia   (g7qq38mx3d58n1b15kcia),
	.demg_fwfkmaeawq30t    (demg_fwfkmaeawq30t ),
	.grtb6ypa0px2gi1c    (grtb6ypa0px2gi1c ),
	.f128d8ws0seoihu1    (f128d8ws0seoihu1 ),

	.m2r7mfmq3afdd1ine   (m2r7mfmq3afdd1ine),
	.nhafiywg3hg_52kogwh   (nhafiywg3hg_52kogwh),
	.xrqayy6vigrw66z8a     (xrqayy6vigrw66z8a  ),
	.jyy72ywt9nbo10f2jxupacld (jyy72ywt9nbo10f2jxupacld),
	.drz92qecqx_qtxwro   (drz92qecqx_qtxwro),
    .hr7la0400ty0hiwk5d0  (g1jacxqkf1oj5l4jvp9a7qacc3),
    .y1ipzdhzcfq282ups6ja  (nj35btypmlzn6n67k5a3sbxlz_),
    .lqv5bv6hq78ov_prb97v5z   (vknrn2pdsorktjh1khqd1o5u ),
    .o15lm7no18top00l32ra  (kul32yktlkh84fqkeuiasdj4c),
    .ly1y__c5rzaa9xv_9_m1ppr  (a0711e1j5ewmq9032iiam6zd),
    .f1msmreidlchd7rf9w625  (yxxau7egbjhe86w26b64yf),
    .uarhtvlb5te5hc2g3   (otv_22s88_efzve7t9aewczn ),
    .g9ayxf51lhjl44vvw62u3  (huhgp41uzpgntu1igqiuh8bpy),
    .qfoijjxktg6dht3klxhyw5g  (glmsykv9_w4rhlqnh8qmvqcu3n),
    .gao2lzva86gawlwp2   (y69op1rhrojqmwt2zvwvt6_w1v ),
    .xpt7vgmhw7tamcpv2l   (qya9tage13i6s6ij4c93w406f ),
    .lrh4lctjvrz1rhm6b9oh   (kbs9xq0ed1rv9h4kn8c9l7v8_c ),
    .pyfc_rgr3cwwvo34pf    (u4pdpnruu01ssoo78t_r),
    .krh62hs2scfnb76m67a    (wpa_w8k78vc5tscpvglay54t),
    .u6xj18ku9lj1890n7   (j_xo5pr2yvkxhr8c7fcp5m),
    .s3lwpy5def9adgbbvx9ct   (o7cx0ajdhtouycxdeb8ly50),
    .q96vjidg4x6ohxl7    (xjpj_prxqbclz5urycgi1vv),
   
    .b6m1vcd7bmemxnu99_zke  (n71nv9q2skeheb436zhxyw8iy),
    .vqld30a8qt13mzhwoc  (ah736xwkrzyalnwp8ow6mi1z),
    .jpa5gwkjwqz_j0a3cy1    (pn6t3ogf6fkiu3lq50zejhq2_  ),
    .kjxe2fpsacp9bx2_0fah36ij(nyapu28mzy38j3qnbv84wn19w  ),
    .xsw8oz2ni13z6vac1tn61  (lfg1njvjoj4o9aupkvjol5f),

    .cv0k9k_ijjnnylw1s7b_0d    (cv0k9k_ijjnnylw1s7b_0d),

    .swpk4h0gei3t_34xogbqncbo4  (swpk4h0gei3t_34xogbqncbo4),

    .u9qmfl3rwx0dhr92z875vx7q  (u9qmfl3rwx0dhr92z875vx7q),
    .unu_x_i6jmr33nz0yitzk   (unu_x_i6jmr33nz0yitzk ),
    .bei3qhdtd0euq2emblogsu_x   (bei3qhdtd0euq2emblogsu_x ),
    .bf0_ynb648lqi7s93eieo0ln  (bf0_ynb648lqi7s93eieo0ln),
    .wf8o7p9_qfthhoxs747wyeuwkky  (wf8o7p9_qfthhoxs747wyeuwkky),
    .ygro7xue7x7rtdafkj3o4q4  (ygro7xue7x7rtdafkj3o4q4),
    .drrly3q0ocg8d4pwh3m9o77   (drrly3q0ocg8d4pwh3m9o77),
    .g654a6a9cesbee7xs6_uu9lu5   (g654a6a9cesbee7xs6_uu9lu5 ),
    .x7fex0jf9da6a5v1c28upl72t   (x7fex0jf9da6a5v1c28upl72t ),
    .ege0_1ufqm8i68zo4il6cwe46d   (ege0_1ufqm8i68zo4il6cwe46d ),
    .ngyxf4n1cpcgks_s2zmgfb260  (ngyxf4n1cpcgks_s2zmgfb260),
    .c7m50uaw8lmp_iv4ci38q2  (c7m50uaw8lmp_iv4ci38q2),
    .m04a1mtbabwezldp1crh4rg6z  (m04a1mtbabwezldp1crh4rg6z),
    .hwjq1ubtaei44lpk609fm2hb8 (hwjq1ubtaei44lpk609fm2hb8),
    .e28p_fu1k484ncul0p85ko     (e28p_fu1k484ncul0p85ko),

    .bvg_3t_ujbpur7b_h7f63jse  (bvg_3t_ujbpur7b_h7f63jse),

    .m5l6wu3uz_jfqasz8e3tsvrm  (m5l6wu3uz_jfqasz8e3tsvrm),
    .g9so28ythfl0q7xnk66p1    (g9so28ythfl0q7xnk66p1  ),
    .e66wluxk71p2ldu3a1qk994bq(e66wluxk71p2ldu3a1qk994bq),
    .ig2roj0y08x8_ntp3knz9rd  (ig2roj0y08x8_ntp3knz9rd),

    .a0_d_zdz9h9fgk46e8arf    (a0_d_zdz9h9fgk46e8arf),

    .twr9y24wxhs3qj2z9f2hzpaig6  (twr9y24wxhs3qj2z9f2hzpaig6),

    .w8b46r9cof57xvd5zo1u4zh8  (w8b46r9cof57xvd5zo1u4zh8),
    .wn1l4cmih7rwce1rb7wk3f9wy   (wn1l4cmih7rwce1rb7wk3f9wy ),
    .cgnzbuo_1yz6v42seb25duv   (cgnzbuo_1yz6v42seb25duv ),
    .zopev7f487spn9mwvuowqo  (zopev7f487spn9mwvuowqo),
    .p32jk0lb8g31kqlpvmllo75qim  (p32jk0lb8g31kqlpvmllo75qim),
    .g973rcaou05i456suvk_89dm  (g973rcaou05i456suvk_89dm),
    .wflv6rhfdwyxttak111v1l   (wflv6rhfdwyxttak111v1l),
    .ggsmt4nzx8pwlowehinqvk60f   (ggsmt4nzx8pwlowehinqvk60f ),
    .xu8494ii8ectqb91224uuer   (xu8494ii8ectqb91224uuer ),
    .r6rk128ijo839ougen9stbe   (r6rk128ijo839ougen9stbe ),
    .xo6ciibewn8p8xey97jcsqi5  (xo6ciibewn8p8xey97jcsqi5),
    .evz1w_girwszyfnlcg4mwvtjo  (evz1w_girwszyfnlcg4mwvtjo),
    .ju5f9fb1erjep_bv8gpfn6  (ju5f9fb1erjep_bv8gpfn6),
    .hadi1_f3quoaotjv5758x8kksot2 (hadi1_f3quoaotjv5758x8kksot2),
    .bdi4gjlb0po4ejcztowoqil7     (bdi4gjlb0po4ejcztowoqil7),

    .m7tq_t57mr5bovbb9ghffl4k  (m7tq_t57mr5bovbb9ghffl4k),

    .gpcgdcri3e6_fxrw8wwtysoqqr  (gpcgdcri3e6_fxrw8wwtysoqqr),
    .a6s4kxg1ibr6mntc85jik    (a6s4kxg1ibr6mntc85jik  ),
    .hizzalmpwr8cqkxqi80wvbt65x(hizzalmpwr8cqkxqi80wvbt65x),


    
    
    
    
    
    
    
    
    
    
    
    


    .p7ah58va5_2njbtv         (p7ah58va5_2njbtv     ),
    .u981qrwkgi5h0e72b__gg19w    (u981qrwkgi5h0e72b__gg19w),
    .p0i2i3v3j1tclelx51        (p0i2i3v3j1tclelx51    ),

                       
                           .mum8f1rtatle7p_55y84     (mum8f1rtatle7p_55y84  ),   
                           .pn5bpwlp5ijfako9m5ao   (pn5bpwlp5ijfako9m5ao),
                           .g3s0qe2adsxsx8e6z     (g3s0qe2adsxsx8e6z  ),
                           .a1rl4lmhqp8ydyk07kqkn    (a1rl4lmhqp8ydyk07kqkn ),       
                           .apnns9jlj7y3y5bg8ynz   (apnns9jlj7y3y5bg8ynz),
                                                                      
                           .pmz7e4mgvbnmimqp0nghk     (pmz7e4mgvbnmimqp0nghk  ),
                           .j61algpxjoycxbswhgsuf   (j61algpxjoycxbswhgsuf),
                           .omq1ehm8hp4q9jgp5n5vn     (omq1ehm8hp4q9jgp5n5vn  ),
                           .fbv1q6sraswzp91zcn    (fbv1q6sraswzp91zcn ),       
                           .jv8kv41vzuir6an4iod   (jv8kv41vzuir6an4iod),
                                                                      
                                                                      
                           .qgl4363n31jx6xjyo05zkn     (qgl4363n31jx6xjyo05zkn  ),
                           .zec78nyllxlfwmpsgncluudf   (zec78nyllxlfwmpsgncluudf),
                           .dwvnjl0vxqkgd8t6dtvg5z    (dwvnjl0vxqkgd8t6dtvg5z ),
                           .gngmcj5c1jd85csel9ntru    (gngmcj5c1jd85csel9ntru ),       
                           .tkt93y5lfluzkia5plvksp   (tkt93y5lfluzkia5plvksp),
                                                                      
                           .km7co8hqm563od8ga_03_g     (km7co8hqm563od8ga_03_g  ),
                           .j4mas6g26o63wvnsdquh8c4p   (j4mas6g26o63wvnsdquh8c4p),
                           .nniah5mh0cunkhyln9    (nniah5mh0cunkhyln9 ),
                           .rcy_v3911lf33nza5j    (rcy_v3911lf33nza5j ),       
                           .g4nfgu53_rgc0632w8z97   (g4nfgu53_rgc0632w8z97),
                                                                      
                           .xzgkclcxsgfuseg87     (xzgkclcxsgfuseg87  ),
                           .djwlah5bo0r6myit6cal0t   (djwlah5bo0r6myit6cal0t),
                           .qu_ju3lv6nvkdbo8h11uf    (qu_ju3lv6nvkdbo8h11uf ),
                           .dydwz9i6k80alqfarffop    (dydwz9i6k80alqfarffop ),       
                           .ql1c7hzoj9kf__7r97krm   (ql1c7hzoj9kf__7r97krm),
                                                                      
                           .kp2j8kv1p1cjcg0lerwm     (kp2j8kv1p1cjcg0lerwm  ),
                           .v4a7g1wh3ivw0esp7dye0oiz   (v4a7g1wh3ivw0esp7dye0oiz),
                           .x9zuk21gpaj58uszvm5    (x9zuk21gpaj58uszvm5 ),
                           .n_h5oz0c5bo5rpevwjcu8    (n_h5oz0c5bo5rpevwjcu8 ),       
                           .ryid4_99ns1jc83at_88x   (ryid4_99ns1jc83at_88x),

    .indfp6mwqdqamez0mex (f2qbwkn13kmm9hmrn159wahi),
    .tia1md5dyh6kj4     (doh50j3p7c7yl7uk9),
    .c4ughu0qm5sfai (c4ughu0qm5sfai),

    .dyl5g2vgrvy4mb3 (dyl5g2vgrvy4mb3),
    .r5hpbriny8m67sv9e_ylgo1   (r5hpbriny8m67sv9e_ylgo1         ),

    .n8mvs5sw2pw48loob7jv6nmjdds(n8mvs5sw2pw48loob7jv6nmjdds),
    .dbzz2cu7abqy43de_ky433v(dbzz2cu7abqy43de_ky433v),
    .y3iin4ygz2ed73_84l91h73(y3iin4ygz2ed73_84l91h73),
    .gbb0bfnz8wqnjr5sufoh6ojt4pr(gbb0bfnz8wqnjr5sufoh6ojt4pr),
    .im70q80i1xh1y_5mo9ndr1 (im70q80i1xh1y_5mo9ndr1 ),

    .mmludd_fnt2yevok8a1a0    (mmludd_fnt2yevok8a1a0),
    .buwj9_8l8bwj80kkinq9p    (buwj9_8l8bwj80kkinq9p),

    .viuu21jzrv          (viuu21jzrv),



    .c0x_72w8ddbpt17fn      (bm7mey1b6dibd5i6lfpukeue),

    .tw0yf9aln_vu06k8l    (a8h5u6ohzhowdrvqrnlllzd70h  ),
    .q84eo09gg53r2jj5a5xn    (pz92yc3xo60c49ayrztvq18a  ),
    .ss4cm882613f24kdjqsyl     (pwzrcrecvxehn8htjdn3kv2d0   ),
    .zm9uosdggg7ntkh97elw    (ksa323b46ngmxwazg70t76  ),
    .g_ahl2zik6mj75atnp_hej    (bs4xe3ath5_4_iwylkfwppp  ),
    .bjl40q8m35dwdn_mn9    (njyud2m27xz7r6j0g0ieq17m  ),
    .oefdpb9h9kx627r_0y5     (m5itqssum7ljklhpn5nvzvd93   ),
    .fh1jm1za5zvqmvdloi    (kkk0rwd1njowzq01nvxke  ),
    .sp_0hv_ae5rrl9vagusi    (a2kttuidwhopy02uoajaf  ),
    .b4oh48a9a0g269ybrm     (g4hx0dbyp7f7ou8x02a0   ),
    .r5s3ykb7_xkl6t12oucf     (zce_icdtm3r9hzeanwhlu3fv   ),
    .ssswxj_bpfx_ebsbj     (jkp1oke9n1q9ikytwx_7k   ),
                                                   
    .fsj22rallxmhdrvuwenpq    (mu3ut_ezr05qz2bbi7_vc_aod  ),
    .yign8d_dhrow0i5wjts4bd    (sk3bm3yc69h4ac84pc4killh  ),
    .hhlfu4md9k5v7naf1qt      (b7g_hkjxumf964flze01v6p    ),
    .j8m9s_du9fk99idlbh80  (cmtnwdaxz9zk1858kalga2vt), 
    .aapsfpke41r7dyya4ah    (qjvmrd1013dapqkahq_f87b  ),

    .y1rlahaedj99shvl6uc      (ndsqg7zrec89ncrv9yu3k    ),

    .rqf8b5xxbw0n1_qaw    (eth8quxx9hhjhxr4u9k2s77f  ),
    .ocwcf75wgxfb1bawe    (zw6mbnvv_8hcztypnytp87v_vy  ),
    .holgl43_yucp7f7l     (l_s_khzs83700pzjuq3_obo44   ),
    .oyev1ipmdflkvxygwr    (kyvscpwy0vljnwysfxqxb  ),
    .ihknw7_lm_572tv6s    (sl5cpfvi658e8pl6nh2cm4  ),
    .o31l03k34sdhwt4lkazfa5    (tmqgi_fx924f3bq8ms4u8t0  ),
    .gy2sgn_1bpkac7msq3     (tcrjx_8vlmtrlqjvk3tu   ),
    .r_1u6q2lzkfus3o9nfl    (y0jaju01t8mqh2ycz05limpxfu  ),
    .yff7wf8wth2vjkdjpr    (x88dy7qz1z117o2jmbslutlpm  ),
    .lppjhpov_5lgvx7n7fm4g     (kykdx6vx9n3hm7k6oybv   ),
    .sdfg9zykj79rz_7thf9k     (b59iokn7e2645ocyqifdk6sp1   ),
    .wt4e4tlh0u_4cljr2j5f9     (xs2l1_f3yynnrl_rw2zbe   ),
  
    .o4wuryrcvw13y2v5m6b6u    (hf8rqlrzsk0e9ho4orde_r  ),
    .bt4howrm5xnf6u4fuwrum6    (opns8_xijy8grr0gygeszh  ),
    .vnqegbzme0jutvf      (hng3_y3ldjtyu4a9n45    ),
    .jdj122rbumyogtin6xpg97  (y1ovf4ea_l0kgs84_pwk6czrs), 
    .p9mcc6npaw32uigcp6    (n6fa00b9i708mtqu7yc9wjvxip  ),


  .ysnexkrvlg2s55ajc5g69tm      (mcfeo0u7nf9     ),           
  .p7832rg37bbm7_ssxunhcj7     (wfa5o72ctktgt55fgv2eo),          
  .t1xtkdoie_8djygqlt1br56pwt    (sa3k3tsgxwqp8z     ),         
  .w33zvryieg8hhgy58581ny437h9 (igeg6alwzopr62ti9),           
  .lv96t6re1w44borcb7do83ndua3vjy (g3e0lri_3krzlfxnnlo_2y82qf),      



    .gf33atgy           (fid1178x5nxb ),
    .ru_wi         (ru_wi        ) 
  );

  urpfdi55wfwmmi3i n_wbwq9kmmbxh (
    .k8qtud5yr1e98g            (k8qtud5yr1e98g   ),
    .mw1zdgavbul7ic            (mw1zdgavbul7ic   ),
    .covjtr51ggzngufqow        (covjtr51ggzngufqow    ),
    .qfhwjs9ygxr4e0rg86a        (qfhwjs9ygxr4e0rg86a    ),
    .r86mhhg0562g6n9sah0z         (r86mhhg0562g6n9sah0z     ),
    .oor8acg0u_d09e0moah       (oor8acg0u_d09e0moah     ),
    .aqz_nh46x0w0rdwc83s7c       (aqz_nh46x0w0rdwc83s7c     ),
    .drgmlg58l2czwg2ijhc           (drgmlg58l2czwg2ijhc),
    .hvgjjhizbfp9km9dd           (hvgjjhizbfp9km9dd),
    .nd1hj8zlmdgys5obof18pe      (nd1hj8zlmdgys5obof18pe     ),
    .oe3uwa3e_ggymrc7ri           (oe3uwa3e_ggymrc7ri),
    .a51im30isjous61asad1lrg5       (a51im30isjous61asad1lrg5),


    .eapsrdy52u                 (a_1o1o8345o28hui     ),
    .slk31s106jz               (t8p1kh0tvb2ej56s  ),



    .vz63qkw5s3m8urb9           (z5vf_v21veoi10ybi   ),
    .iojqlhtwx45_siz            (tq4dt8fbx7xch3x4b   ),
    .ydtm1yuxqj7fmxvqc            (ip_8jolx6gnp   ),

    .jfsrn6g5wjvu1s            (kzfv878bfk6iooqik),
    .a726ykhkw2fkfxd            (o3cx5caf3g3nzd0pu),
    .sml00v8pmuueefw             (woxzhk095h66amt5),
    .ewg8titgu69y7lmx0j             (n4bind2sncm8mh),
    .hz3c9eiwgzw2hb              (wtw3apxzccvxdx8 ),
    .p4pen8le4jxeud_b           (zckohvd58ff_pyuth),
    .mxu7x8rtlq0kewjvcl           (qfx1o1rp7psuvaq),
    .xbzkx8ucmech               (j11k71dn8a),
    .ehkpciu6l7p               (fov_crsecs),
    .jm0nv8cdtqhyk5t2ddht          (avaoxa8z58nyr0g127g),
    .oo04o1rrd2a               (yc8cklg0l),
    .eqedamf6p97lmc2ywq            (mb94n_xsixgup9p0),
    .b0ylmw5xa8oytsw3j6n        (b0ylmw5xa8oytsw3j6n),
















    .gf33atgy           (c8fchlpwl ),
    .ru_wi         (ru_wi ) 
  );



 u52cit50_7l ryz1p9vyh_azra(

    .xmbe_e4vm6ofjbn7lq        (xmbe_e4vm6ofjbn7lq),

    .nv5a7f_68p9ebw             (nv5a7f_68p9ebw),
    .cv0k9k_ijjnnylw1s7b_0d (cv0k9k_ijjnnylw1s7b_0d),
    .swpk4h0gei3t_34xogbqncbo4 (swpk4h0gei3t_34xogbqncbo4),
    .u9qmfl3rwx0dhr92z875vx7q (u9qmfl3rwx0dhr92z875vx7q),
    .unu_x_i6jmr33nz0yitzk (unu_x_i6jmr33nz0yitzk), 
    .bei3qhdtd0euq2emblogsu_x (bei3qhdtd0euq2emblogsu_x), 
    .bf0_ynb648lqi7s93eieo0ln (bf0_ynb648lqi7s93eieo0ln),
    .wf8o7p9_qfthhoxs747wyeuwkky (wf8o7p9_qfthhoxs747wyeuwkky),
    .ygro7xue7x7rtdafkj3o4q4 (ygro7xue7x7rtdafkj3o4q4),
    .drrly3q0ocg8d4pwh3m9o77 (drrly3q0ocg8d4pwh3m9o77),
    .g654a6a9cesbee7xs6_uu9lu5 (g654a6a9cesbee7xs6_uu9lu5),
    .x7fex0jf9da6a5v1c28upl72t (x7fex0jf9da6a5v1c28upl72t),
    .ege0_1ufqm8i68zo4il6cwe46d (ege0_1ufqm8i68zo4il6cwe46d),
    .ngyxf4n1cpcgks_s2zmgfb260 (ngyxf4n1cpcgks_s2zmgfb260), 
    .c7m50uaw8lmp_iv4ci38q2 (c7m50uaw8lmp_iv4ci38q2), 
    .m04a1mtbabwezldp1crh4rg6z (m04a1mtbabwezldp1crh4rg6z), 
    .hwjq1ubtaei44lpk609fm2hb8 (hwjq1ubtaei44lpk609fm2hb8), 
    .e28p_fu1k484ncul0p85ko (e28p_fu1k484ncul0p85ko), 
    .a0_d_zdz9h9fgk46e8arf (a0_d_zdz9h9fgk46e8arf),
    .twr9y24wxhs3qj2z9f2hzpaig6 (twr9y24wxhs3qj2z9f2hzpaig6),
    .w8b46r9cof57xvd5zo1u4zh8 (w8b46r9cof57xvd5zo1u4zh8),
    .wn1l4cmih7rwce1rb7wk3f9wy (wn1l4cmih7rwce1rb7wk3f9wy), 
    .cgnzbuo_1yz6v42seb25duv (cgnzbuo_1yz6v42seb25duv), 
    .zopev7f487spn9mwvuowqo (zopev7f487spn9mwvuowqo),
    .p32jk0lb8g31kqlpvmllo75qim (p32jk0lb8g31kqlpvmllo75qim),
    .g973rcaou05i456suvk_89dm (g973rcaou05i456suvk_89dm),
    .wflv6rhfdwyxttak111v1l (wflv6rhfdwyxttak111v1l),
    .ggsmt4nzx8pwlowehinqvk60f (ggsmt4nzx8pwlowehinqvk60f),
    .xu8494ii8ectqb91224uuer (xu8494ii8ectqb91224uuer),
    .r6rk128ijo839ougen9stbe (r6rk128ijo839ougen9stbe),
    .xo6ciibewn8p8xey97jcsqi5 (xo6ciibewn8p8xey97jcsqi5), 
    .evz1w_girwszyfnlcg4mwvtjo (evz1w_girwszyfnlcg4mwvtjo), 
    .ju5f9fb1erjep_bv8gpfn6 (ju5f9fb1erjep_bv8gpfn6), 
    .hadi1_f3quoaotjv5758x8kksot2 (hadi1_f3quoaotjv5758x8kksot2), 
    .bdi4gjlb0po4ejcztowoqil7 (bdi4gjlb0po4ejcztowoqil7), 
    .bvg_3t_ujbpur7b_h7f63jse (bvg_3t_ujbpur7b_h7f63jse),
    .m5l6wu3uz_jfqasz8e3tsvrm (m5l6wu3uz_jfqasz8e3tsvrm),
    .g9so28ythfl0q7xnk66p1   (g9so28ythfl0q7xnk66p1  ),
    .e66wluxk71p2ldu3a1qk994bq (e66wluxk71p2ldu3a1qk994bq),
    .ig2roj0y08x8_ntp3knz9rd (ig2roj0y08x8_ntp3knz9rd), 
    .m7tq_t57mr5bovbb9ghffl4k (m7tq_t57mr5bovbb9ghffl4k),
    .gpcgdcri3e6_fxrw8wwtysoqqr (gpcgdcri3e6_fxrw8wwtysoqqr),
    .a6s4kxg1ibr6mntc85jik   (a6s4kxg1ibr6mntc85jik  ),
    .hizzalmpwr8cqkxqi80wvbt65x (hizzalmpwr8cqkxqi80wvbt65x),


































    .rsgiw0g_vwk7sxen_4zrphe7    (x27lqkgq55knwoqsc6_bn0p), 
    .ghredfib76bt_a9caiytel4    (ud5ygg9b8pmm93drtbfk4l8hv),
    .neuurwim9m_f3o_6nal7q7ft     (f_lrqmtz5mpqmbrhn6f05[32-1:0] ),
    .i0bh8gwxh68vtael53ff2y_ir5x    (czjipv9hqkdx4jllt3ajsl),
    .e41m_8qgi_o4t4e2_v4c6pxn5g4    (j92g3e8ublsg2d9sjj_i3),
    .rkkjbx03o1tifh3uilzkztfkb    (af3a5ot65per6f87crwmj),
    .gzq7xf16ajsco5h0qj7civq    (bjucsszqg5d1sc5etnwvf1),
    .lpf8x_t3lmkkdri3nbex80     (ss92bd8t5gyfjfl1_lp2 ),
    .si54q2nl6njfvmi6thon6_0    (64'b0),
    .ppe31c4mhmxn9qqmpibp3ohumo2h    ({8{1'b0}}),
    .dp41iy8ngtqmissjqvvy10ihu     (1'b0 ),
    .aum4efqs_h1yct3n53gypfa     (1'b0 ),
    .rpje1avuaivhahlv82bint       (t37flu99i5ex1j3e_8   ),
    .j_iw8afyzfudhp5xe0v8v231     (wvjkzp74fi8ed7nnr7xlm3gt),
    .smpikn1zm93setxcwgrzoiybl8    (z1beclu7k0_h4nn6njz05sbe1),
    .a6jqkrqyut1oz9lpndklbhv     (w1i6s2iwu2nnj7idywd ),

    .bygw_825g7_dt283loevm5zym41e    (phzkntckzzbndu4wevf1o6), 
    .ir3fzbymkf93yhmjzi8gfgeq0    (1'b1), 
    .c0st8ve3a3f8xhdx147o8      (bpyef3a0dnkkyqdpymy  ),
    .h4r65p765_t877awntcuf03d6d3    (ba1ucnyekcm68i9wuqwmn),
    .wglnz1ixornvjx16dv6bvtdx6zpf  (),


    .wex3zbl1x6s4be1en    (wex3zbl1x6s4be1en    ),   
	.pszbl2iobld50k    (pszbl2iobld50k    ),
	.vfuu2l_7oof31qn0_a    (vfuu2l_7oof31qn0_a    ),
	.bvy9o58rgxtbjz_xph     (bvy9o58rgxtbjz_xph     ),
	.gcpthp2sfxb3cxo     (gcpthp2sfxb3cxo     ),
	.xzjdk5deciqs4l3my_l    (xzjdk5deciqs4l3my_l    ),
	.dlg9f36umgj9xdv0wa    (dlg9f36umgj9xdv0wa    ),
	.peug05ptx4vv93u4xc     (peug05ptx4vv93u4xc     ),
	.yienty7ycnc25au    (yienty7ycnc25au    ),
	.j2amhrzbhku8dzd    (j2amhrzbhku8dzd    ),
	.rxlx2eq69oye0ba3     (rxlx2eq69oye0ba3     ),




     .wh6iy6zpdqsnv2y (wh6iy6zpdqsnv2y),
     .bd6yatp5cqq (bd6yatp5cqq),
     .fl1qsvyu (fl1qsvyu),
     .b9889wezsu (b9889wezsu),
     .an__mxugc4 (an__mxugc4),
     .poj6g8vw9e (poj6g8vw9e),
     .dafaivw3ze9g3hi (dafaivw3ze9g3hi),
     .q2c0d6fxz_1bw (q2c0d6fxz_1bw),
     .wblesminvapwua (wblesminvapwua),
     .v3cim36gj8g (v3cim36gj8g),
     .ss22f8fuy2uhr (ss22f8fuy2uhr),
     .hoaoalj5pcdnpnm0 (hoaoalj5pcdnpnm0),
     .rh8f1e3jgg3xi (rh8f1e3jgg3xi),
     .roral7fym4h3_ (roral7fym4h3_),
     .b_gwvq35iq0_yvk (b_gwvq35iq0_yvk),
     .lqm2hm0cjm5zt (lqm2hm0cjm5zt),
     .f3n3tpjs44e0_ (f3n3tpjs44e0_),
     .dmc59hxf352z (dmc59hxf352z),
     .a63l3og_8qak5jy (a63l3og_8qak5jy),
     .m0wp58qmji79 (m0wp58qmji79),
     .c8qmnfk1vqai (c8qmnfk1vqai),
     .pbov8g9yizcwr (pbov8g9yizcwr),
     .t8qjehupeajtzjr (t8qjehupeajtzjr),
     .hhp1rh0x0jn (hhp1rh0x0jn),
     .w9yptl69xj6p (w9yptl69xj6p),
     .yvcpy_gyehs4lji (yvcpy_gyehs4lji), 
     .kted7ph0krq (kted7ph0krq),
     .a93i3d2hji (a93i3d2hji),
     .of5p5cb8p4 (of5p5cb8p4),
     .g1bi1xzuv64 (g1bi1xzuv64),
     .gj6p5b5ik3r9p (gj6p5b5ik3r9p),
     .m1fmaas4oww6 (m1fmaas4oww6),
     .hjstsi51gm (hjstsi51gm),
     .onpqhy0s69 (onpqhy0s69),
     .aw7xjbi (aw7xjbi),
     .z0cc2y_uzoh_ (z0cc2y_uzoh_),
     .y8tc_vywu82ugn (y8tc_vywu82ugn),
     .o2h9d51o6m6 (o2h9d51o6m6),
     .nneek3ep5xykwl (nneek3ep5xykwl),
     .g8khua4l0y77zjp (g8khua4l0y77zjp),
     .wmlp1a2b (wmlp1a2b),
     .weop50xb_avne (weop50xb_avne),
     .su81e8dxdzng9d (su81e8dxdzng9d),

    .gf33atgy                    (klwwlfrft ),
    .ru_wi                  (ru_wi ) 
  );

  xsz0s4xbnv9 hci4safv376(

    .bebngvg8sove         (bebngvg8sove),

    .g1jacxqkf1oj5l4jvp9a7qacc3  (g1jacxqkf1oj5l4jvp9a7qacc3),
    .nj35btypmlzn6n67k5a3sbxlz_  (nj35btypmlzn6n67k5a3sbxlz_),
    .vknrn2pdsorktjh1khqd1o5u   (vknrn2pdsorktjh1khqd1o5u ),
    .kul32yktlkh84fqkeuiasdj4c  (kul32yktlkh84fqkeuiasdj4c),
    .a0711e1j5ewmq9032iiam6zd  (a0711e1j5ewmq9032iiam6zd),
    .yxxau7egbjhe86w26b64yf  (yxxau7egbjhe86w26b64yf),
    .otv_22s88_efzve7t9aewczn   (otv_22s88_efzve7t9aewczn ),
    .huhgp41uzpgntu1igqiuh8bpy  (huhgp41uzpgntu1igqiuh8bpy),
    .glmsykv9_w4rhlqnh8qmvqcu3n  (glmsykv9_w4rhlqnh8qmvqcu3n),
    .y69op1rhrojqmwt2zvwvt6_w1v   (y69op1rhrojqmwt2zvwvt6_w1v ),
    .qya9tage13i6s6ij4c93w406f   (qya9tage13i6s6ij4c93w406f ),
    .kbs9xq0ed1rv9h4kn8c9l7v8_c   (kbs9xq0ed1rv9h4kn8c9l7v8_c ),
    .rqfuzid60p8me07wm6bsjailb  (3'b000),
    .fsro6vxjx57ptgecek7dolel   (2'b0 ),
    .wpa_w8k78vc5tscpvglay54t    (wpa_w8k78vc5tscpvglay54t),
    .u4pdpnruu01ssoo78t_r    (u4pdpnruu01ssoo78t_r),
    .j_xo5pr2yvkxhr8c7fcp5m    (j_xo5pr2yvkxhr8c7fcp5m),
    .o7cx0ajdhtouycxdeb8ly50    (o7cx0ajdhtouycxdeb8ly50),
    .xjpj_prxqbclz5urycgi1vv    (xjpj_prxqbclz5urycgi1vv),

    .n71nv9q2skeheb436zhxyw8iy  (n71nv9q2skeheb436zhxyw8iy),
    .ah736xwkrzyalnwp8ow6mi1z  (ah736xwkrzyalnwp8ow6mi1z),
    .pn6t3ogf6fkiu3lq50zejhq2_    (pn6t3ogf6fkiu3lq50zejhq2_  ),
    .nyapu28mzy38j3qnbv84wn19w(nyapu28mzy38j3qnbv84wn19w),
    .lfg1njvjoj4o9aupkvjol5f  (lfg1njvjoj4o9aupkvjol5f),




    .lueem7uei21mn66 (lueem7uei21mn66) ,  
    .vgodhub5af4gihqv5eef (vgodhub5af4gihqv5eef) ,  
    .lueqjwqinfpts52  (lueqjwqinfpts52 ) ,  
    .lv9moee8_5_8dsy5  (lv9moee8_5_8dsy5 ) ,  
    .ck0wbvgghs6n9j4 (ck0wbvgghs6n9j4) ,  
    .uecfgtalcganlj42vmq  (uecfgtalcganlj42vmq ) ,
    .msxgfr_x73l96858p1s (msxgfr_x73l96858p1s) ,  
    .tze074ath5y6h2m41  (tze074ath5y6h2m41 ) ,  
    .o752t3g6xbcxc6if88wi (o752t3g6xbcxc6if88wi) , 

    .nprvxoyk8ecm174bi8 (nprvxoyk8ecm174bi8) , 





    .ooqxby68qkbvkc5xteznb_x     (ooqxby68qkbvkc5xteznb_x),
    .zhr6liff5rm5wfulyyq     (zhr6liff5rm5wfulyyq),
    .xlsvmbo_v42zk9mypgihxz      (xlsvmbo_v42zk9mypgihxz ),
    .pzv82u11m6kxelyx220ilq5     (pzv82u11m6kxelyx220ilq5),
    .yhhbbaf9pqjys_bjgq6h4gj     (yhhbbaf9pqjys_bjgq6h4gj),
    .qbaqr2mf9nkictp7plgs     (qbaqr2mf9nkictp7plgs),
    .ijehxhtls_byykogg4h      (ijehxhtls_byykogg4h ),
    .ylsn7ect00nktb3n8gy6     (ylsn7ect00nktb3n8gy6),
    .etkmv0abc25lclz_o85     (etkmv0abc25lclz_o85),
    .cdpiwio563kpzebanibgl9      (),
    .r7w0ije3_ym7bdontco40e      (),
    .z8dedxyz7e4q36qmy70p      (),
    .y6swa_2gtejyczns_62cex     (),
    .urjwk5dc302d8z5nlzwb      (),
    
    .txrvwlqb8aeb5k6eo4p0tb2     (txrvwlqb8aeb5k6eo4p0tb2),
    .q8mbpl9ben1u54xn_d     (q8mbpl9ben1u54xn_d),
    .igk23ds0cu4_sziqf       (igk23ds0cu4_sziqf  ),
    .jkzbkg87eqm75wurn5snetjvg   (1'b0),
    .rsvzuajc8qp4__n0807     (rsvzuajc8qp4__n0807),

    .sc9dq6vpj_vb3unfw0     (sc9dq6vpj_vb3unfw0),
    .ni7lsi0fuchbbgfizw0l     (ni7lsi0fuchbbgfizw0l),
    .cvmgqobwfiy_kwo814x      (cvmgqobwfiy_kwo814x ),
    .h_htd26ozpf1rjy0gsvy     (h_htd26ozpf1rjy0gsvy),
    .gbzyzsndu75k8rua21_v9c     (gbzyzsndu75k8rua21_v9c),
    .w2e5ixihsvl50pgq6b4      (w2e5ixihsvl50pgq6b4 ),
    .tl_6em2dyajt9yrv4j794c     (tl_6em2dyajt9yrv4j794c),
    .mf1rr9vurug23q2qsrv     (mf1rr9vurug23q2qsrv),
    .ob4qe7emnlqe4zaoqvitt      (),
    .gmquwxhk5rxcr7xq57zcn      (),
    .nqeg1hcgcuxu2idsy840      (),
    .q0wbro_xv81_o_wumr3x5     (),
    .dessj2xl2_xq3mvaz438      (),
    
    .m1vcvvn1ntgzmmwe1bse     (m1vcvvn1ntgzmmwe1bse),
    .f20ikomgiyzoonhphcz     (f20ikomgiyzoonhphcz),
    .q7emifz3jwxt_jv0_w       (q7emifz3jwxt_jv0_w  ),
    .qc2wdr75ushg0r17szgvi9   (1'b0),
    .l1hbm4iglo7pz0pdg_ayjs     (l1hbm4iglo7pz0pdg_ayjs),

    .l9z66pxhit_o_1iyjp     (l9z66pxhit_o_1iyjp),
    .jdh22q4xq9e7wiznv     (jdh22q4xq9e7wiznv),
    .y_z_yc9_f4ppblmsch3z5      (y_z_yc9_f4ppblmsch3z5 ),
    .yc7tq3wh6q569ueq7i07em     (yc7tq3wh6q569ueq7i07em),
    .yfy18a1ju6mptqd0_u     (yfy18a1ju6mptqd0_u),
    .gducqncehu9g7n4lydij_0     (gducqncehu9g7n4lydij_0),
    .nmp2x4e8pl59l6he_f9_      (nmp2x4e8pl59l6he_f9_ ),
    .dd_gpw58ph81_864rnspr     (dd_gpw58ph81_864rnspr),
    .nhzg88_kzsk0fbtrtku     (nhzg88_kzsk0fbtrtku),
    .ar4vri2lev87gi9oug      (),
    .tzz1dn20stpsz4u3v      (),
    .meku6m0blkiklu01zs      (),
    .epjio2a09p_ymmxo_a     (),
    .uyh1mgy24c2cjlh4      (),
    
    .ixpwz6oo67i61vepd74     (ixpwz6oo67i61vepd74),
    .t7hb1k3tkjzooetwf     (t7hb1k3tkjzooetwf),
    .da2pgeraioxt6edc       (da2pgeraioxt6edc  ),
    .rf5x6hqfa2yhnqvhegzhfkh   (1'b0),
    .u2fwd1l2_bdiuiftn     (u2fwd1l2_bdiuiftn),

    .gf33atgy                    (oi60pknul ),
    .ru_wi                  (ru_wi ) 
  );





xnkv2ixv6wqo  gzynxggryaz6cnb(
    .ru_wi                           (ru_wi                             ),
    .gf33atgy                             (h87jx93oz7                           ),
    .g3ljqli3ukatw2132ssx              (moqs2k81l9fugde5v_581              ),
    .trtkzwpsx6l                      (trtkzwpsx6l                        ),
    .qhne8m65goz1y091ss8              (bz8qao4o4xqslni1d3                ),
    .z83wiqsi0hgv                      (vpecdc5kos                        ), 
    .r6p4z7df65i25fz                    (pccd7o463jfc_dpc5va                 ), 
    .mqi6hv3p07axtj                    (k5ovx8tintgvetip                      ), 
    .zgpvz622wmbpuyplhsxe2y               (f97le_hyejv7saw9vslna                 ), 
    .h7x7oqrhyprsd9fpyf7ukcq              (yruel3nusosm39gnmb9ev_                ), 
    .q4u0u5t961_a5u67h7zrv            (oeux55k_cre0he7w7jip5b1              ), 
    .qn5go609a7uekpxe4               (r8z2r_ud53zj8mrpk                 ), 
    .uxqm4y8nwwoy7a4manunpmrxz2a         (bu1949pq_9946o1_e2q_uvr8p4           ), 
    .tjdyq2su0gawzvcig32cszgu749r         (b4isf5u8b8pj34e09f72vxe38zg           ), 
    .qjkug4xiqzawij13384vr4              (docsdqb0rnb9fmmgf3                ), 
    .pb3pms28fol8dfr0gr8dkit         (xyqctztl2_la5wbp2an04mw           ), 
    .cj92o34fmt9lj4qchqzk6arhow       (du_nrgluldn3gf5tg1wa8slreks         ), 
    .qr21q8rwg0cu                    (vn9mhiqoo1jrmofqr4xn               ), 
    .g1400sa7kyme0jubnk7du               (w8mlksniwgqyojf1iy                 ), 
    .l875nvn0_y6wu72ui7ogut             (b518xebdeds3frng6hy4g               ), 
    .j9xmer7ue4wnuw7ba9gy              (moj77icm1kmex0900                    ), 
    .kqjz41lwlrrv                      (hib0x0rvcjwnn75a                     ),
    .ha7j195sl8e_t5                    (cgmsm8wvxc5kg90xwvwq0cga              ),                 
    .t0xxoojg_0iodq0py               (w9mx37ezcezieq_9__94o              ), 
    .mm9g9a4egd29oz9vvgscmya              (hsnr3xtposirc7pmphtiko3xlz         ), 
    .qouo17x2sfmp8hi9d3pto43t1            (k1jkhgd9bvypwrti7ietjp0n7_nyzu       ), 
    .l5xpteag34o1wqsgx               (qirelbyt49gkn46_f24yxtc               ), 
    .g2vry3iwllflk3zzplwitn3eq7gc         (jq4wiwydrozelhpru9snvs0             ),
    .ilj8lhiujxv57r4qqghj0_nntz         (j6muxslh7pud3298q9d8lc2             ), 
    .z1l_kkshyf_56cwmaq2dm           (z1l_kkshyf_56cwmaq2dm             ), 
    .w7u50np_chxy7wq5n9et_q           (w7u50np_chxy7wq5n9et_q             ), 
    .l2dse4sd3runnrb1rcbydauc            (l2dse4sd3runnrb1rcbydauc              ),  
    .kr1rhzlb5gr_wty1pe392s5oqet        (kr1rhzlb5gr_wty1pe392s5oqet          ), 
    .ox2ptuhum_e2aodz8wine6h         (ox2ptuhum_e2aodz8wine6h           ), 
    .g_qmxgznvfin609fmm97kuc2dm02         (g_qmxgznvfin609fmm97kuc2dm02           ), 
    .i9oln6xm1pi9dzsd61s1kg4dmo7j         (i9oln6xm1pi9dzsd61s1kg4dmo7j           ), 
   
    .yf_5vs18cke5xg660my              (yf_5vs18cke5xg660my                ), 
    .sneofd4rq3b0m9eu91r8                 (sneofd4rq3b0m9eu91r8                   ),
    .d6vb8lyc7vlnm0o3arpqw68r            (uzklqlncpqqm1rav                      ), 
    .pxmnhz1pxp2i2mmdb6540            (ortueunvnkx_l5m_j                      ), 
    .pfeolrpx0uzt9jq1ndjruu_            (hwuhtb7ucto_utk56                      ), 
    .xa286l0j7185h2h8cym8            (i1env2kmns7qvvuuc                      ), 
    .vs6zhd0u5jdq_fconvsekj            (g3s3vpafvy3i                      ), 
    .n9tjosvoxai4p0sj6mb                 (pcr4upio7_tx37                         ), 
    .i0acx70llka5qu09r5jd                 (i0acx70llka5qu09r5jd                   ),
    .e44u8ctdv_z5u19to                 (e44u8ctdv_z5u19to                   ), 
    .h7k_k0xxi7vktla                 (h7k_k0xxi7vktla                   ), 
    .v_vouzmjecsvtjxt                 (v_vouzmjecsvtjxt                   ), 
    .ef9y8yyld9onuy00de7o              (ef9y8yyld9onuy00de7o                ), 
    .ammhazyeeglt3ewt4p              (ammhazyeeglt3ewt4p                ), 
    .xvwzwg7_3ek2tx                   (xvwzwg7_3ek2tx                     ), 
    .y8sg6kbsyavoh4usiqn               (y8sg6kbsyavoh4usiqn                 ), 
    .gnqkycbjc0k9k4_edoube               (gnqkycbjc0k9k4_edoube                 ), 
    .xib8tki1lzl05e71ry               (xib8tki1lzl05e71ry                 ), 
    .hdle8ta5fimb1inf1z               (hdle8ta5fimb1inf1z                 ), 
    .trtxm7l0l_kp36i9y                (trtxm7l0l_kp36i9y                  ),
    .p0akg_4worvsnfq_q36vp                (p0akg_4worvsnfq_q36vp                  ),
    .mqdc73rtez0bzh2_1                  (mqdc73rtez0bzh2_1                    ), 
    .vl5p5iump0rpm1hbr               (vl5p5iump0rpm1hbr                 ), 
    .oj6rvjf7ujgb34264               (oj6rvjf7ujgb34264                 ), 
    .vjfz03uzu8p_0jhhvvev               (vjfz03uzu8p_0jhhvvev                 ), 
    .p1qeemcgwrrzzt73bl               (p1qeemcgwrrzzt73bl                 ),
    .ertspxpg0txqgp9i6fx53               (ertspxpg0txqgp9i6fx53                 ),
    .z3xt8rx_qs6z0goo1                 (z3xt8rx_qs6z0goo1                   ),
    .ln7r12q36ofpcd6m6u                (ln7r12q36ofpcd6m6u                  )
);






    assign u_ll4hq1b12s2i1 = w41ourymsjpvm8q1e;


endmodule                                      























module xsz0s4xbnv9(

  output                         bebngvg8sove,
  
  
  
  input                          g1jacxqkf1oj5l4jvp9a7qacc3,
  output                         nj35btypmlzn6n67k5a3sbxlz_,
  input  [32-1:0]   vknrn2pdsorktjh1khqd1o5u, 
  input                          otv_22s88_efzve7t9aewczn, 
  input  [32-1:0]        huhgp41uzpgntu1igqiuh8bpy,
  input  [4-1:0]      glmsykv9_w4rhlqnh8qmvqcu3n,
  input  [2:0]                   rqfuzid60p8me07wm6bsjailb,
  input  [1:0]                   fsro6vxjx57ptgecek7dolel,
  input                          y69op1rhrojqmwt2zvwvt6_w1v,
  input                          qya9tage13i6s6ij4c93w406f,
  input  [1:0]                   kbs9xq0ed1rv9h4kn8c9l7v8_c,
  input                          kul32yktlkh84fqkeuiasdj4c, 
  input                          a0711e1j5ewmq9032iiam6zd, 
  input                          yxxau7egbjhe86w26b64yf, 
  input                          u4pdpnruu01ssoo78t_r, 
  input                          j_xo5pr2yvkxhr8c7fcp5m, 
  input                          o7cx0ajdhtouycxdeb8ly50,
  input                          wpa_w8k78vc5tscpvglay54t, 
  input                          xjpj_prxqbclz5urycgi1vv, 
  
  output                         n71nv9q2skeheb436zhxyw8iy,
  input                          ah736xwkrzyalnwp8ow6mi1z,
  output                         pn6t3ogf6fkiu3lq50zejhq2_  ,
  output                         nyapu28mzy38j3qnbv84wn19w,
  output [32-1:0]        lfg1njvjoj4o9aupkvjol5f,

    
  
  output                         l9z66pxhit_o_1iyjp,
  input                          jdh22q4xq9e7wiznv,
  output [32-1:0]   y_z_yc9_f4ppblmsch3z5, 
  output                         nmp2x4e8pl59l6he_f9_, 
  output [32-1:0]        dd_gpw58ph81_864rnspr,
  output [4-1:0]      nhzg88_kzsk0fbtrtku,
  output [2:0]                   epjio2a09p_ymmxo_a,
  output [1:0]                   uyh1mgy24c2cjlh4,
  output                         ar4vri2lev87gi9oug,
  output                         tzz1dn20stpsz4u3v,
  output [1:0]                   meku6m0blkiklu01zs,
  output                         yc7tq3wh6q569ueq7i07em, 
  output                         yfy18a1ju6mptqd0_u, 
  output                         gducqncehu9g7n4lydij_0, 
  
  
  input                          ixpwz6oo67i61vepd74,
  output                         t7hb1k3tkjzooetwf,
  input                          da2pgeraioxt6edc  ,
  input                          rf5x6hqfa2yhnqvhegzhfkh,
  input  [32-1:0]        u2fwd1l2_bdiuiftn,

      
  
  output                         ooqxby68qkbvkc5xteznb_x,
  input                          zhr6liff5rm5wfulyyq,
  output [32-1:0]   xlsvmbo_v42zk9mypgihxz, 
  output                         ijehxhtls_byykogg4h, 
  output [32-1:0]        ylsn7ect00nktb3n8gy6,
  output [4-1:0]      etkmv0abc25lclz_o85,
  output [2:0]                   y6swa_2gtejyczns_62cex,
  output [1:0]                   urjwk5dc302d8z5nlzwb,
  output                         cdpiwio563kpzebanibgl9,
  output                         r7w0ije3_ym7bdontco40e,
  output [1:0]                   z8dedxyz7e4q36qmy70p,
  output                         pzv82u11m6kxelyx220ilq5, 
  output                         yhhbbaf9pqjys_bjgq6h4gj, 
  output                         qbaqr2mf9nkictp7plgs, 
  
  
  input                          txrvwlqb8aeb5k6eo4p0tb2,
  output                         q8mbpl9ben1u54xn_d,
  input                          igk23ds0cu4_sziqf  ,
  input                          jkzbkg87eqm75wurn5snetjvg,
  input  [32-1:0]        rsvzuajc8qp4__n0807,


      
  
  output                         sc9dq6vpj_vb3unfw0,
  input                          ni7lsi0fuchbbgfizw0l,
  output [32-1:0]   cvmgqobwfiy_kwo814x, 
  output                         w2e5ixihsvl50pgq6b4, 
  output [32-1:0]        tl_6em2dyajt9yrv4j794c,
  output [4-1:0]      mf1rr9vurug23q2qsrv,
  output [2:0]                   q0wbro_xv81_o_wumr3x5,
  output [1:0]                   dessj2xl2_xq3mvaz438,
  output                         ob4qe7emnlqe4zaoqvitt,
  output                         gmquwxhk5rxcr7xq57zcn,
  output [1:0]                   nqeg1hcgcuxu2idsy840,
  output                         h_htd26ozpf1rjy0gsvy, 
  output                         gbzyzsndu75k8rua21_v9c, 
  
  
  input                          m1vcvvn1ntgzmmwe1bse,
  output                         f20ikomgiyzoonhphcz,
  input                          q7emifz3jwxt_jv0_w  ,
  input                          qc2wdr75ushg0r17szgvi9,
  input  [32-1:0]        l1hbm4iglo7pz0pdg_ayjs,

  
  
  
  


  output [1:0]                   lueem7uei21mn66  ,  
  output                         vgodhub5af4gihqv5eef  ,  
  output [32-1:0]   lueqjwqinfpts52   ,  
  output [2:0]                   lv9moee8_5_8dsy5   ,  
  output [32-1:0]        ck0wbvgghs6n9j4  ,  
  output [3:0]                   uecfgtalcganlj42vmq   ,

  input  [32-1:0]        msxgfr_x73l96858p1s  ,  
  input  [1:0]                   tze074ath5y6h2m41   ,  
  input                          o752t3g6xbcxc6if88wi  ,  

  input                          nprvxoyk8ecm174bi8,


  input  gf33atgy,
  input  ru_wi
  );

  wire                         pz0q76ea_yiq3saws0z;
  wire                         af1vxcl5oex51d4gyi;
  wire [32-1:0]   ls7uc9xf_3_8qydto9c; 
  wire                         nnrcvgi4rjznrrjwsmfil; 
  wire [32-1:0]        xlr_1ussy71yinbg7iq;
  wire [4-1:0]      tcx5fhw92rxev45vp_eu;
  wire [2:0]                   irkxveoohccdbiuan0j;
  wire [1:0]                   sju7tc0kopo4lzwi_p1;
  wire                         fogsi4b5xwfjpe40xo96;
  wire                         wqooosnjio96iiecemj5;
  wire [1:0]                   fca60sudk287naxrfp;
  wire                         ybuoa7610v5vhluwnr6; 
  wire                         sje1v6_k812gs7c8vi4xhl; 
  wire                         p1z2bh3236unk7cfygp3; 
  
  wire                         fgp78l66kwouy_i3u;
  wire                         b7hycfm6whjnvn1zfcash6;
  wire                         plc0t8yx2zh5r1guqv  ;
  wire                         i7w52vtyh_v977qowyu_ju = 1'b0;
  wire [32-1:0]        ysrx86ke5yal46xmk;

























  localparam uc1_xpj8fyv3o5 = 0;

  localparam nfv2_7mn_l8sejrk = (uc1_xpj8fyv3o5 + 1);

  localparam x7g6e_ye_nr3yy = (nfv2_7mn_l8sejrk + 1);

  localparam lco1nzyasf1przhj = (x7g6e_ye_nr3yy + 1);


  localparam f7wqn6iss2tplp4a = (lco1nzyasf1przhj + 1);

  localparam tgongp9jmy57cyf = f7wqn6iss2tplp4a;

  localparam k_18vva78gwxfmb93wt = 2;


  localparam s3xvyho = 8;
  localparam y61y499cunmtec= 0;
  localparam a69a9ho1_kmpwc58n= 1;
  localparam kmj83muj1f9gt  = 2;
  localparam iqktc22qa2x4xf0zy  = 3;
  localparam vu69rf8t84hai  = 4;
  localparam ksdqvndai1tu41  = 5;
  localparam h4xfhp090mye  = 6;
  localparam qn77zdua2lv05_= 7;

  wire [s3xvyho-1:0] o5g1fg0iksctvgahi118;
  assign o5g1fg0iksctvgahi118[y61y499cunmtec] = yxxau7egbjhe86w26b64yf; 
  assign o5g1fg0iksctvgahi118[a69a9ho1_kmpwc58n] = kul32yktlkh84fqkeuiasdj4c;
  assign o5g1fg0iksctvgahi118[qn77zdua2lv05_] = a0711e1j5ewmq9032iiam6zd;

  assign o5g1fg0iksctvgahi118[kmj83muj1f9gt  ] = u4pdpnruu01ssoo78t_r;

  assign o5g1fg0iksctvgahi118[iqktc22qa2x4xf0zy  ] = j_xo5pr2yvkxhr8c7fcp5m;
                                           
  assign o5g1fg0iksctvgahi118[vu69rf8t84hai  ] = o7cx0ajdhtouycxdeb8ly50;
                                           
  assign o5g1fg0iksctvgahi118[h4xfhp090mye  ] = wpa_w8k78vc5tscpvglay54t;
                                           

  assign o5g1fg0iksctvgahi118[ksdqvndai1tu41  ] = 1'b0;
                                           

  wire c6kkvm_h8s0mvx4ftuhp;
  wire hrbp69rjgu_d2z82pu;
  wire [32-1:0] w_pgye9mqq713nhkax;
  wire schp22no0ojsdix6_p;
  wire [32-1:0] v7wulnc5uiem1r_nope;
  wire [4-1:0] ecvhc6gcpfteg133dys6;
  wire [2:0] mroyh40g9dv1yei_fz;
  wire [1:0] vf1q5jg437v0wixmm;
  wire zt4adl9qxxedlvknaqi58;
  wire yr0c7ctrmhb_movc;
  wire [1:0] ho91hs321kw4nilurz89;
  wire [s3xvyho-1:0] no3in967u5raf7fs9kl;


  wire xln1wnk65jj86mqgmi;
  wire m9qvkyy1wrqn4dhpgl_jq;
  wire q30nvrqaexwf_wontxwn;
  wire hd9f4_dsbj2z8sjxpcuemku;
  wire [32-1:0] m9pi4njc3tc3c0qjgurmsa;

  wire zmzpuim70lsljt2ccu2c1;

  ux607_gnrl_icb_buffer # (
    .OUTS_CNT_W   (4),
    .AW    (32),
    .DW    (32), 
    .CMD_DP(1),
    .RSP_DP(0),
      
      
      
    .RSP_ALWAYS_READY (0),

    .CMD_CUT_READY (0),
    .RSP_CUT_READY (0),
    .USR_W (s3xvyho)
  )l6zy02rbz_ljdt8b_ng(
    .bus_clk_en (1'b1),
    .icb_buffer_active      (zmzpuim70lsljt2ccu2c1),
    .i_icb_cmd_valid        (g1jacxqkf1oj5l4jvp9a7qacc3),
    .i_icb_cmd_ready        (nj35btypmlzn6n67k5a3sbxlz_),
    .i_icb_cmd_read         (otv_22s88_efzve7t9aewczn ),
    .i_icb_cmd_addr         (vknrn2pdsorktjh1khqd1o5u ),
    .i_icb_cmd_wdata        (huhgp41uzpgntu1igqiuh8bpy),
    .i_icb_cmd_wmask        (glmsykv9_w4rhlqnh8qmvqcu3n),
    .i_icb_cmd_lock         (y69op1rhrojqmwt2zvwvt6_w1v ),
    .i_icb_cmd_excl         (qya9tage13i6s6ij4c93w406f ),
    .i_icb_cmd_size         (kbs9xq0ed1rv9h4kn8c9l7v8_c ),
    .i_icb_cmd_burst        (rqfuzid60p8me07wm6bsjailb),
    .i_icb_cmd_beat         (fsro6vxjx57ptgecek7dolel ),
    .i_icb_cmd_usr          (o5g1fg0iksctvgahi118  ),
                     
    .i_icb_rsp_valid        (n71nv9q2skeheb436zhxyw8iy),
    .i_icb_rsp_ready        (ah736xwkrzyalnwp8ow6mi1z),
    .i_icb_rsp_err          (pn6t3ogf6fkiu3lq50zejhq2_  ),
    .i_icb_rsp_excl_ok      (nyapu28mzy38j3qnbv84wn19w),
    .i_icb_rsp_rdata        (lfg1njvjoj4o9aupkvjol5f),
    .i_icb_rsp_usr          (),
    
    .o_icb_cmd_valid        (c6kkvm_h8s0mvx4ftuhp),
    .o_icb_cmd_ready        (hrbp69rjgu_d2z82pu),
    .o_icb_cmd_read         (schp22no0ojsdix6_p ),
    .o_icb_cmd_addr         (w_pgye9mqq713nhkax ),
    .o_icb_cmd_wdata        (v7wulnc5uiem1r_nope),
    .o_icb_cmd_wmask        (ecvhc6gcpfteg133dys6),
    .o_icb_cmd_lock         (zt4adl9qxxedlvknaqi58 ),
    .o_icb_cmd_excl         (yr0c7ctrmhb_movc ),
    .o_icb_cmd_size         (ho91hs321kw4nilurz89 ),
    .o_icb_cmd_burst        (mroyh40g9dv1yei_fz),
    .o_icb_cmd_beat         (vf1q5jg437v0wixmm ),
    .o_icb_cmd_usr          (no3in967u5raf7fs9kl),
                         
    .o_icb_rsp_valid        (xln1wnk65jj86mqgmi),
    .o_icb_rsp_ready        (m9qvkyy1wrqn4dhpgl_jq),
    .o_icb_rsp_err          (q30nvrqaexwf_wontxwn  ),
    .o_icb_rsp_excl_ok      (hd9f4_dsbj2z8sjxpcuemku),
    .o_icb_rsp_rdata        (m9pi4njc3tc3c0qjgurmsa),
    .o_icb_rsp_usr          ({s3xvyho{1'b0}}  ),

    .clk                    (gf33atgy  ),
    .rst_n                  (ru_wi)
  );

 localparam mp26klefy4v2f = (32 + 2);


 
      
      
 wire                  zxvzk3_vgha5csgrrci6;
 wire                  gra9m8aonyccam2vtm6;
 wire                  gve831mbnld8ehisxrlrzk  ;
 wire                  lfd_p_beayl64b7h_g1h06dxs7;
 wire [32-1:0] d3ope9_k74q0c5awum24;

 wire [mp26klefy4v2f-1:0]a4fqa0u_cepdttsvjrtf0;
 wire [mp26klefy4v2f-1:0]q_9sg5nf6yh37omtsfxb;

  assign a4fqa0u_cepdttsvjrtf0 = {
                          i7w52vtyh_v977qowyu_ju,
                          plc0t8yx2zh5r1guqv,
                          ysrx86ke5yal46xmk
                          };

  assign {
                          lfd_p_beayl64b7h_g1h06dxs7,
                          gve831mbnld8ehisxrlrzk,
                          d3ope9_k74q0c5awum24
                          } = q_9sg5nf6yh37omtsfxb;


















assign q_9sg5nf6yh37omtsfxb = a4fqa0u_cepdttsvjrtf0;
assign zxvzk3_vgha5csgrrci6 = fgp78l66kwouy_i3u;
assign b7hycfm6whjnvn1zfcash6 = gra9m8aonyccam2vtm6;





  wire [s3xvyho-1:0] cc6x6p9zm9w_vfzqo_;
  wire [s3xvyho-1:0] tcv8dplxxgphst24g3s9;
  wire [s3xvyho-1:0] fyk4yj3a2b33ox73va9k;
  wire [s3xvyho-1:0] fnuyvj6i24mxzajq;

  assign gducqncehu9g7n4lydij_0 = cc6x6p9zm9w_vfzqo_[y61y499cunmtec];
  assign yc7tq3wh6q569ueq7i07em = cc6x6p9zm9w_vfzqo_[a69a9ho1_kmpwc58n];
  assign yfy18a1ju6mptqd0_u = cc6x6p9zm9w_vfzqo_[qn77zdua2lv05_];
  assign qbaqr2mf9nkictp7plgs = tcv8dplxxgphst24g3s9[y61y499cunmtec];
  assign pzv82u11m6kxelyx220ilq5 = tcv8dplxxgphst24g3s9[a69a9ho1_kmpwc58n];
  assign yhhbbaf9pqjys_bjgq6h4gj = tcv8dplxxgphst24g3s9[qn77zdua2lv05_];
  assign gbzyzsndu75k8rua21_v9c = fyk4yj3a2b33ox73va9k[y61y499cunmtec];
  assign h_htd26ozpf1rjy0gsvy = fyk4yj3a2b33ox73va9k[a69a9ho1_kmpwc58n];
  assign p1z2bh3236unk7cfygp3 = fnuyvj6i24mxzajq[y61y499cunmtec];
  assign ybuoa7610v5vhluwnr6 = fnuyvj6i24mxzajq[a69a9ho1_kmpwc58n];
  assign sje1v6_k812gs7c8vi4xhl = fnuyvj6i24mxzajq[qn77zdua2lv05_];

  wire [tgongp9jmy57cyf*1-1:0] fgaj26ic3vlyw4_j9cd2e9iw5e5;
  wire [tgongp9jmy57cyf*1-1:0] fo2e9fa1xtekqy_rau1jvp;
  wire [tgongp9jmy57cyf*32-1:0] yn3_ae3lzkj5xi4qm4r12;
  wire [tgongp9jmy57cyf*1-1:0] oo66a5i9yj7eu97xzyjljzo4m;
  wire [tgongp9jmy57cyf*32-1:0] t0xc_soqbh3onidnjvuak5;
  wire [tgongp9jmy57cyf*4-1:0] hb58z51gm9p0robvubcqsio45n7;
  wire [tgongp9jmy57cyf*3-1:0] k6_7qe0217bxabwti931g5pf;
  wire [tgongp9jmy57cyf*2-1:0] mqpao8z9f30uq2rzuys2zt;
  wire [tgongp9jmy57cyf*1-1:0] j016rws5wewra_ent6uzmgq8;
  wire [tgongp9jmy57cyf*1-1:0] ubwy6_856dlynocswg3b0h3;
  wire [tgongp9jmy57cyf*2-1:0] ujjmevva2mtja2eiajfdu;
  wire [tgongp9jmy57cyf*s3xvyho-1:0] ous1ovavtg25yc9cmar2;

  wire [tgongp9jmy57cyf*1-1:0] zw0jju5nmyaae6lkudb1rc8zsh;
  wire [tgongp9jmy57cyf*1-1:0] hjab85nvos0ly5k7d5qc0a3n;
  wire [tgongp9jmy57cyf*1-1:0] eihugo5lxty1ao1uxvhn68jh;
  wire [tgongp9jmy57cyf*1-1:0] ph3072ol08mqn_adsird67uf1;
  wire [tgongp9jmy57cyf*32-1:0] qzru8eufkdrjwbh5j3iayridl0j;

  wire tw05v8cq;
  wire stl2dyg;
  wire gep6mi;
  wire vvzkx7j;
  wire vp658_;
  wire fszy_tyz45;
  wire kzwqi4u2o;
  wire vb6z8hdlvds;
  wire yqtyvnmn35;
  wire tqf0jhuhh3;
  wire n41ts9l;
  wire uyb_dpr4jei;
  wire rsvim4n7wky;
  wire yq4gyp3pb7p;
  wire ct3ez8g;
  wire kjfys9rmr7;
  wire o09x3joq73tu;

  
  assign {tw05v8cq
                           , ooqxby68qkbvkc5xteznb_x
                           , sc9dq6vpj_vb3unfw0
                           , l9z66pxhit_o_1iyjp
                           , pz0q76ea_yiq3saws0z
                           } = {1'b0,fgaj26ic3vlyw4_j9cd2e9iw5e5};


  assign {stl2dyg
                           , xlsvmbo_v42zk9mypgihxz
                           , cvmgqobwfiy_kwo814x
                           , y_z_yc9_f4ppblmsch3z5
                           , ls7uc9xf_3_8qydto9c
                           } = {1'b0,yn3_ae3lzkj5xi4qm4r12};

  assign {gep6mi
                           , ijehxhtls_byykogg4h
                           , w2e5ixihsvl50pgq6b4
                           , nmp2x4e8pl59l6he_f9_
                           , nnrcvgi4rjznrrjwsmfil
                           } = {1'b0,oo66a5i9yj7eu97xzyjljzo4m};

  assign {vvzkx7j
                           , ylsn7ect00nktb3n8gy6
                           , tl_6em2dyajt9yrv4j794c
                           , dd_gpw58ph81_864rnspr
                           , xlr_1ussy71yinbg7iq
                           } = {1'b0,t0xc_soqbh3onidnjvuak5};

  assign {vp658_
                           , etkmv0abc25lclz_o85
                           , mf1rr9vurug23q2qsrv
                           , nhzg88_kzsk0fbtrtku
                           , tcx5fhw92rxev45vp_eu
                           } = {1'b0,hb58z51gm9p0robvubcqsio45n7};
                         
  assign {fszy_tyz45
                           , y6swa_2gtejyczns_62cex
                           , q0wbro_xv81_o_wumr3x5
                           , epjio2a09p_ymmxo_a
                           , irkxveoohccdbiuan0j
                           } = {1'b0,k6_7qe0217bxabwti931g5pf};
                         
  assign {kzwqi4u2o
                           , urjwk5dc302d8z5nlzwb
                           , dessj2xl2_xq3mvaz438
                           , uyh1mgy24c2cjlh4
                           , sju7tc0kopo4lzwi_p1
                           } = {1'b0,mqpao8z9f30uq2rzuys2zt};
                         
  assign {vb6z8hdlvds
                           , cdpiwio563kpzebanibgl9
                           , ob4qe7emnlqe4zaoqvitt
                           , ar4vri2lev87gi9oug
                           , fogsi4b5xwfjpe40xo96
                           } = {1'b0,j016rws5wewra_ent6uzmgq8};

  assign {yqtyvnmn35
                           , r7w0ije3_ym7bdontco40e
                           , gmquwxhk5rxcr7xq57zcn
                           , tzz1dn20stpsz4u3v
                           , wqooosnjio96iiecemj5
                           } = {1'b0,ubwy6_856dlynocswg3b0h3};
                           
  assign {tqf0jhuhh3
                           , z8dedxyz7e4q36qmy70p
                           , nqeg1hcgcuxu2idsy840
                           , meku6m0blkiklu01zs
                           , fca60sudk287naxrfp
                           } = {1'b0,ujjmevva2mtja2eiajfdu};

  assign {n41ts9l
                           , tcv8dplxxgphst24g3s9
                           , fyk4yj3a2b33ox73va9k
                           , cc6x6p9zm9w_vfzqo_
                           , fnuyvj6i24mxzajq
                           } = {1'b0,ous1ovavtg25yc9cmar2};

  assign {uyb_dpr4jei,fo2e9fa1xtekqy_rau1jvp} = {1'b0
                           , zhr6liff5rm5wfulyyq
                           , ni7lsi0fuchbbgfizw0l
                           , jdh22q4xq9e7wiznv
                           , af1vxcl5oex51d4gyi
                           };

  
  assign {rsvim4n7wky,zw0jju5nmyaae6lkudb1rc8zsh} = {1'b0
                           , txrvwlqb8aeb5k6eo4p0tb2
                           , m1vcvvn1ntgzmmwe1bse
                           , ixpwz6oo67i61vepd74
                           , zxvzk3_vgha5csgrrci6
                           };

  assign {yq4gyp3pb7p,eihugo5lxty1ao1uxvhn68jh} = {1'b0
                           , igk23ds0cu4_sziqf
                           , q7emifz3jwxt_jv0_w
                           , da2pgeraioxt6edc
                           , gve831mbnld8ehisxrlrzk
                           };

  assign {ct3ez8g,ph3072ol08mqn_adsird67uf1} = {1'b0
                           , jkzbkg87eqm75wurn5snetjvg
                           , qc2wdr75ushg0r17szgvi9
                           , rf5x6hqfa2yhnqvhegzhfkh
                           , lfd_p_beayl64b7h_g1h06dxs7
                           };

  assign {kjfys9rmr7,qzru8eufkdrjwbh5j3iayridl0j} = {1'b0
                           , rsvzuajc8qp4__n0807
                           , l1hbm4iglo7pz0pdg_ayjs
                           , u2fwd1l2_bdiuiftn
                           , d3ope9_k74q0c5awum24
                           };

  assign {o09x3joq73tu
                           , q8mbpl9ben1u54xn_d
                           , f20ikomgiyzoonhphcz
                           , t7hb1k3tkjzooetwf
                           , gra9m8aonyccam2vtm6
                           } = {1'b0,hjab85nvos0ly5k7d5qc0a3n};

  wire ct75ug06hab3z6y9_m = no3in967u5raf7fs9kl[kmj83muj1f9gt];
  wire k6we617nhpxx8v2uk = ct75ug06hab3z6y9_m;

  wire t317bq_xu7d4mqzeg668 = no3in967u5raf7fs9kl[iqktc22qa2x4xf0zy];
  wire kyi9z2trwg8bx7tq2 = t317bq_xu7d4mqzeg668;

  wire im9c8rgr5s9xufp0iv = no3in967u5raf7fs9kl[vu69rf8t84hai];
  wire b_017b1lvxz4dy4d2ygiv = im9c8rgr5s9xufp0iv;


  wire ymoolxn883auk6omt = no3in967u5raf7fs9kl[h4xfhp090mye];
  wire oofsawkm35y3hfigea2u = ymoolxn883auk6omt;

  
  
  
  
  
  
  
  
  


  wire yr_a1y9a_rx_;
  wire [tgongp9jmy57cyf-1:0] d5vywzwdg84jz7ffdy3;

  assign {yr_a1y9a_rx_, d5vywzwdg84jz7ffdy3} = 
      {                    1'b0
                           , kyi9z2trwg8bx7tq2
                           , b_017b1lvxz4dy4d2ygiv
                           , k6we617nhpxx8v2uk
                           , oofsawkm35y3hfigea2u
      };

  ux607_gnrl_icb_splt # (
  .ALLOW_DIFF (0),
  .ALLOW_0CYCL_RSP (1),
                       
                       
  .FIFO_OUTS_NUM   (8),
  .FIFO_CUT_READY  (1),
  .SPLT_NUM   (tgongp9jmy57cyf),
  .SPLT_PTR_W (tgongp9jmy57cyf),
  .SPLT_PTR_1HOT (1),
  .VLD_MSK_PAYLOAD(1), 
  .USR_W      (s3xvyho),
  .AW         (32),
  .DW         (32) 
  ) jjv9u5yznto7e30(
  .i_icb_splt_indic       (d5vywzwdg84jz7ffdy3),        

  .splt_active            (),

  .i_icb_cmd_valid        (c6kkvm_h8s0mvx4ftuhp )     ,
  .i_icb_cmd_ready        (hrbp69rjgu_d2z82pu )     ,
  .i_icb_cmd_read         (schp22no0ojsdix6_p )      ,
  .i_icb_cmd_addr         (w_pgye9mqq713nhkax )      ,
  .i_icb_cmd_wdata        (v7wulnc5uiem1r_nope )     ,
  .i_icb_cmd_wmask        (ecvhc6gcpfteg133dys6)      ,
  .i_icb_cmd_burst        (mroyh40g9dv1yei_fz)     ,
  .i_icb_cmd_beat         (vf1q5jg437v0wixmm )     ,
  .i_icb_cmd_excl         (yr0c7ctrmhb_movc )     ,
  .i_icb_cmd_lock         (zt4adl9qxxedlvknaqi58 )     ,
  .i_icb_cmd_size         (ho91hs321kw4nilurz89 )     ,
  .i_icb_cmd_usr          (no3in967u5raf7fs9kl  )     ,
 
  .i_icb_rsp_valid        (xln1wnk65jj86mqgmi )     ,
  .i_icb_rsp_ready        (m9qvkyy1wrqn4dhpgl_jq )     ,
  .i_icb_rsp_err          (q30nvrqaexwf_wontxwn)        ,
  .i_icb_rsp_excl_ok      (hd9f4_dsbj2z8sjxpcuemku)    ,
  .i_icb_rsp_rdata        (m9pi4njc3tc3c0qjgurmsa )     ,
  .i_icb_rsp_usr          ( )     ,
                               
  .o_bus_icb_cmd_ready    (fo2e9fa1xtekqy_rau1jvp ) ,
  .o_bus_icb_cmd_valid    (fgaj26ic3vlyw4_j9cd2e9iw5e5 ) ,
  .o_bus_icb_cmd_read     (oo66a5i9yj7eu97xzyjljzo4m )  ,
  .o_bus_icb_cmd_addr     (yn3_ae3lzkj5xi4qm4r12 )  ,
  .o_bus_icb_cmd_wdata    (t0xc_soqbh3onidnjvuak5 ) ,
  .o_bus_icb_cmd_wmask    (hb58z51gm9p0robvubcqsio45n7)  ,
  .o_bus_icb_cmd_burst    (k6_7qe0217bxabwti931g5pf),
  .o_bus_icb_cmd_beat     (mqpao8z9f30uq2rzuys2zt ),
  .o_bus_icb_cmd_excl     (ubwy6_856dlynocswg3b0h3 ),
  .o_bus_icb_cmd_lock     (j016rws5wewra_ent6uzmgq8 ),
  .o_bus_icb_cmd_size     (ujjmevva2mtja2eiajfdu ),
  .o_bus_icb_cmd_usr      (ous1ovavtg25yc9cmar2  ),
  
  .o_bus_icb_rsp_valid    (zw0jju5nmyaae6lkudb1rc8zsh ) ,
  .o_bus_icb_rsp_ready    (hjab85nvos0ly5k7d5qc0a3n ) ,
  .o_bus_icb_rsp_err      (eihugo5lxty1ao1uxvhn68jh)    ,
  .o_bus_icb_rsp_excl_ok  (ph3072ol08mqn_adsird67uf1),
  .o_bus_icb_rsp_rdata    (qzru8eufkdrjwbh5j3iayridl0j ) ,
  .o_bus_icb_rsp_usr      ({tgongp9jmy57cyf*s3xvyho{1'b0}}) ,
                             
  .clk                    (gf33atgy  )                     ,
  .rst_n                  (ru_wi)
  );

  wire d5fptzj7eskpoasxbduz;
  wire s16c0l3pa7ub_oo_2jmrxr77;


  assign bebngvg8sove = g1jacxqkf1oj5l4jvp9a7qacc3 | zmzpuim70lsljt2ccu2c1 
                     | d5fptzj7eskpoasxbduz | s16c0l3pa7ub_oo_2jmrxr77
                     ;

  


  wire                         v1dkb0e2nhwi3g_j34xpdv8c_;
  wire                         r00zov76zpty2mri16x4;
  wire [32-1:0]   skeknqq48f5ld2vnziie; 
  wire                         eea954idskf_wqod3j5h; 
  wire [32-1:0]        sohljey9h_v3mp19sf75mhqpk;
  wire [4-1:0]     lm47iysydszdfaxg5m4_cvm_;
  wire [1:0]                   z9x463flxmgc7yh4khxe0e;
  wire                         wppo0loytrfty8mll2kz;
  wire                         b5ue_g94ax9ldwgpwy95gov3a; 
  wire                         tusx8jw5mkhn9x3hma54; 
  wire                         bshrogt1nai6olo5ohc313tp; 
  
  wire                         jt307hz8c8pbufs1ujddcw2qu;
  wire                         na917ddgwn7f6oal6zmxa;
  wire                         juc2a8pw404przuh0hjf2u  ;
  
  wire [32-1:0]        vq2w4x14h6t5y82wj2vye_8;

  gg8y0ynhq316osuxxk11w2j04po # (
    .hejad2_b4dywimoxw5 (0),
    .evi4vkasjp742kf4 (1),
    .ys68i6_dw7b2m2   (4),
    .nm_fj    (32),
    .onr7l    (32), 
    .xrvos0msri0(2),
    .b8vod12(2),
      
      
      
    .w1ztl72rp0snpfsmgyhg (1),

    .q8s6zigflsp6aqc4dx (0),
    .m4i6t98hqvrs_enkod (0),
    .s3xvyho (3)
  )ohc1dnqsrxmp57f7rbcarm_(
    .aqamddt_moiuy           (1'b1), 
    .rlwva_uzdseg           (nprvxoyk8ecm174bi8), 

    .zmzpuim70lsljt2ccu2c1      (d5fptzj7eskpoasxbduz), 

    .v9ov1b3vn5k4ctkb        (pz0q76ea_yiq3saws0z),
    .ub9pjiu4juf6nuqoq2w6        (af1vxcl5oex51d4gyi),
    .ogvavqa7ta836s         (nnrcvgi4rjznrrjwsmfil ),
    .aw0a19a967dn7n0x25w         (ls7uc9xf_3_8qydto9c ),
    .sc169gxpr38lpe8        (xlr_1ussy71yinbg7iq),
    .hg1g2yh6yktfe_btdst7        (tcx5fhw92rxev45vp_eu),
    .h6hn_gz20krea1         (fogsi4b5xwfjpe40xo96 ),
    .l089k6vccrfphrtw         (1'b0 ),
    .leieaos4fnc5s_81kr         (fca60sudk287naxrfp ),
    .j4d0rl87t28yrb94i        (3'b0),
    .k994rox28a17feu         (2'b0),
    .qku53_e41ce0r6rtb          ({sje1v6_k812gs7c8vi4xhl,ybuoa7610v5vhluwnr6,p1z2bh3236unk7cfygp3}),
                     
    .dy9ll1o6t6ytby71hf4        (fgp78l66kwouy_i3u),   
    .ow4hbh48f0mt6le4o        (b7hycfm6whjnvn1zfcash6),   
    .uzwj715coelxmfqs          (plc0t8yx2zh5r1guqv  ),     
    .sihcnyg6z96riwnnw_np      (                 ), 
    .dek0xt7q6guk2vf6        (ysrx86ke5yal46xmk),
    .efi4ga746crcrx          (),
    
    .me2s8h5yw65ail5        (v1dkb0e2nhwi3g_j34xpdv8c_),
    .dtyl4o87hqhm03wj57        (r00zov76zpty2mri16x4),
    .xiyx61_yd314uojrls         (eea954idskf_wqod3j5h ),
    .k68zoq6vpu0olvs99f         (skeknqq48f5ld2vnziie ),
    .m63rlc2ixlaphiq        (sohljey9h_v3mp19sf75mhqpk),
    .drdtbfa60cpn5ihc        (lm47iysydszdfaxg5m4_cvm_),
    .da5mm7z1qer9hx385ck         (wppo0loytrfty8mll2kz ),
    .tg7q7ezs0lgu3bv36l4         (                    ),
    .hycxa49k327vm1ncjh         (z9x463flxmgc7yh4khxe0e ),
    .rnrkzgtukyiil52jqbp7        (                    ),
    .wta_51f6oa6zy5t         (                    ),
    .vzw7nivk4j2idd          ({b5ue_g94ax9ldwgpwy95gov3a,tusx8jw5mkhn9x3hma54,bshrogt1nai6olo5ohc313tp}),
                         
    .mg6xxata423v5aaikz4v        (jt307hz8c8pbufs1ujddcw2qu),
    .yuew3x5jdkrr87g        (na917ddgwn7f6oal6zmxa),
    .nkx3bwv604xt1          (juc2a8pw404przuh0hjf2u  ),
    .db9kwedxc8ekbwcenl8s9      (1'b0                ),
    .lbvrc0jeu6t70bw        (vq2w4x14h6t5y82wj2vye_8),
    .wxjl9xtjejiyjn1          (3'h0                ),

    .gf33atgy                    (gf33atgy  ),
    .ru_wi                  (ru_wi)
  );

  wire [3:0] p_91br3q3b7mx9zqeweih;

  assign p_91br3q3b7mx9zqeweih[0] = 1'b1;
  assign p_91br3q3b7mx9zqeweih[1] = tusx8jw5mkhn9x3hma54 | b5ue_g94ax9ldwgpwy95gov3a; 
  assign p_91br3q3b7mx9zqeweih[2] = 1'b0; 
  assign p_91br3q3b7mx9zqeweih[3] = 1'b0;


 ux607_gnrl_icb2ahbl
  #(
      .SUPPORT_LOCK     (0),
      .AW(32),
      .DW(32) 
    ) q6oby79npl2tnmlo9fb(
    .icb2ahbl_pend_active(s16c0l3pa7ub_oo_2jmrxr77),
    .bus_clk_en        (nprvxoyk8ecm174bi8), 
    .icb_cmd_valid     (v1dkb0e2nhwi3g_j34xpdv8c_),  
    .icb_cmd_ready     (r00zov76zpty2mri16x4),  
    .icb_cmd_read      (eea954idskf_wqod3j5h ), 
    .icb_cmd_addr      (skeknqq48f5ld2vnziie ), 
    .icb_cmd_wdata     (sohljey9h_v3mp19sf75mhqpk),  
    .icb_cmd_wmask     (lm47iysydszdfaxg5m4_cvm_), 
    .icb_cmd_size      (z9x463flxmgc7yh4khxe0e ),
    .icb_cmd_lock      (wppo0loytrfty8mll2kz),
    .icb_cmd_excl      (1'b0),
    .icb_cmd_burst     (3'b0),
    .icb_cmd_hseq      (1'b0),
    .icb_cmd_hprot     (p_91br3q3b7mx9zqeweih), 
    .icb_cmd_attri     (2'b0), 
    .icb_cmd_dmode     (bshrogt1nai6olo5ohc313tp), 
                       
    .icb_rsp_valid     (jt307hz8c8pbufs1ujddcw2qu),  
    
    .icb_rsp_err       (juc2a8pw404przuh0hjf2u  ),
    .icb_rsp_excl_ok   (                    ),
    .icb_rsp_rdata     (vq2w4x14h6t5y82wj2vye_8),  
                      
    .ahbl_htrans       (lueem7uei21mn66  ),  
    .ahbl_hwrite       (vgodhub5af4gihqv5eef  ),  
    .ahbl_haddr        (lueqjwqinfpts52   ),  
    .ahbl_hsize        (lv9moee8_5_8dsy5   ),  
    .ahbl_hlock        (                 ), 
    .ahbl_hexcl        (                 ), 
    .ahbl_hburst       (                 ),  
    .ahbl_hwdata       (ck0wbvgghs6n9j4  ),  
    .ahbl_hprot        (uecfgtalcganlj42vmq   ),
    .ahbl_hattri       (                 ),
    .ahbl_master       (                 ),
    .ahbl_hrdata       (msxgfr_x73l96858p1s  ),  
    .ahbl_hresp        (tze074ath5y6h2m41   ),  
    .ahbl_hresp_exok   (1'b0             ),  
    .ahbl_hready       (o752t3g6xbcxc6if88wi  ),  
       
    .clk               (gf33atgy),
    .rst_n             (ru_wi)
  );



endmodule




















module u52cit50_7l (
  
  input                          cv0k9k_ijjnnylw1s7b_0d,

  input                          swpk4h0gei3t_34xogbqncbo4,
  output                         u9qmfl3rwx0dhr92z875vx7q,
  input  [32-1:0]   unu_x_i6jmr33nz0yitzk, 
  input                          bei3qhdtd0euq2emblogsu_x, 
  input  [64-1:0]        bf0_ynb648lqi7s93eieo0ln,
  input  [8-1:0]     wf8o7p9_qfthhoxs747wyeuwkky,
  input  [2:0]                   ygro7xue7x7rtdafkj3o4q4,
  input  [1:0]                   drrly3q0ocg8d4pwh3m9o77,
  input                          g654a6a9cesbee7xs6_uu9lu5,
  input                          x7fex0jf9da6a5v1c28upl72t,
  input  [1:0]                   ege0_1ufqm8i68zo4il6cwe46d,
  input                          ngyxf4n1cpcgks_s2zmgfb260, 
  
  input                          c7m50uaw8lmp_iv4ci38q2, 
  
  input                          m04a1mtbabwezldp1crh4rg6z, 
  input                          hwjq1ubtaei44lpk609fm2hb8, 
  
  input                          e28p_fu1k484ncul0p85ko,
  
  
  
  input                          a0_d_zdz9h9fgk46e8arf,

  input                          twr9y24wxhs3qj2z9f2hzpaig6,
  output                         w8b46r9cof57xvd5zo1u4zh8,
  input  [32-1:0]   wn1l4cmih7rwce1rb7wk3f9wy, 
  input                          cgnzbuo_1yz6v42seb25duv, 
  input  [64-1:0]        zopev7f487spn9mwvuowqo,
  input  [8-1:0]     p32jk0lb8g31kqlpvmllo75qim,
  input  [2:0]                   g973rcaou05i456suvk_89dm,
  input  [1:0]                   wflv6rhfdwyxttak111v1l,
  input                          ggsmt4nzx8pwlowehinqvk60f,
  input                          xu8494ii8ectqb91224uuer,
  input  [1:0]                   r6rk128ijo839ougen9stbe,
  input                          xo6ciibewn8p8xey97jcsqi5, 
  
  input                          evz1w_girwszyfnlcg4mwvtjo, 
  
  input                          ju5f9fb1erjep_bv8gpfn6, 
  input                          hadi1_f3quoaotjv5758x8kksot2, 
  
  input                          bdi4gjlb0po4ejcztowoqil7,
  
  
  
  
  
  output                         bvg_3t_ujbpur7b_h7f63jse,
  input                          m5l6wu3uz_jfqasz8e3tsvrm,
  output                         g9so28ythfl0q7xnk66p1  ,
  output                         e66wluxk71p2ldu3a1qk994bq,
  output [64-1:0]        ig2roj0y08x8_ntp3knz9rd, 
  
  output                         m7tq_t57mr5bovbb9ghffl4k,
  input                          gpcgdcri3e6_fxrw8wwtysoqqr,
  output                         a6s4kxg1ibr6mntc85jik  ,
  output                         hizzalmpwr8cqkxqi80wvbt65x,

  input                          xmbe_e4vm6ofjbn7lq,
  output                         nv5a7f_68p9ebw,

 
 
 
 
 
 
 
 
 
 
 
 
 
 
 
 
 
 
 
 
 
 
 
 
 
 
 
 
 
 
 
 
 
  input                          rsgiw0g_vwk7sxen_4zrphe7, 
  output                         ghredfib76bt_a9caiytel4,
  input    [32-1:0] neuurwim9m_f3o_6nal7q7ft, 
  input                          lpf8x_t3lmkkdri3nbex80,
  input  [64-1:0]        si54q2nl6njfvmi6thon6_0,
  input  [8-1:0]     ppe31c4mhmxn9qqmpibp3ohumo2h,
  input    [2:0]                 smpikn1zm93setxcwgrzoiybl8,
  input    [1:0]                 a6jqkrqyut1oz9lpndklbhv,
  input                          dp41iy8ngtqmissjqvvy10ihu,
  input                          aum4efqs_h1yct3n53gypfa,
  input  [1:0]                   j_iw8afyzfudhp5xe0v8v231,
  input                          rpje1avuaivhahlv82bint, 
  input                          i0bh8gwxh68vtael53ff2y_ir5x, 
  
  input                          e41m_8qgi_o4t4e2_v4c6pxn5g4, 
  
  input                          gzq7xf16ajsco5h0qj7civq, 
  input                          rkkjbx03o1tifh3uilzkztfkb, 

  output                         bygw_825g7_dt283loevm5zym41e, 
  input                          ir3fzbymkf93yhmjzi8gfgeq0,
  output                         c0st8ve3a3f8xhdx147o8, 
  output                         wglnz1ixornvjx16dv6bvtdx6zpf,
  output   [64-1:0]      h4r65p765_t877awntcuf03d6d3,
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  output              		 wex3zbl1x6s4be1en,   
  output [1:0]        		 pszbl2iobld50k,   
  output              		 vfuu2l_7oof31qn0_a,   
  output [32    -1:0] bvy9o58rgxtbjz_xph,    
  output [2:0]        		 gcpthp2sfxb3cxo,
  output [2:0]        		 xzjdk5deciqs4l3my_l,
  output [3:0]        		 peug05ptx4vv93u4xc, 
  output [64    -1:0]    dlg9f36umgj9xdv0wa,   
  input  [64    -1:0]    yienty7ycnc25au,   
  input  [1:0]        		 rxlx2eq69oye0ba3,    
  input               		 j2amhrzbhku8dzd,  
  
  input                         wh6iy6zpdqsnv2y,
  output                        bd6yatp5cqq,
  output [4-1:0]         fl1qsvyu,
  output [32-1:0]  b9889wezsu,
  output [7:0]                  an__mxugc4,
  output [2:0]                  poj6g8vw9e,
  output [1:0]                  dafaivw3ze9g3hi,
  output [1:0]                  q2c0d6fxz_1bw,
  output [3:0]                  wblesminvapwua,
  output [2:0]                  v3cim36gj8g,
  output [3:0]                  ss22f8fuy2uhr,
  output [3:0]                  hoaoalj5pcdnpnm0,
  output [1-1:0]           rh8f1e3jgg3xi,
  
  input                         roral7fym4h3_,
  output                        b_gwvq35iq0_yvk,
  output [4-1:0]         lqm2hm0cjm5zt,
  output [32-1:0]  f3n3tpjs44e0_,
  output [7:0]                  dmc59hxf352z,
  output [2:0]                  a63l3og_8qak5jy,
  output [1:0]                  m0wp58qmji79,
  output [1:0]                  c8qmnfk1vqai,
  output [3:0]                  pbov8g9yizcwr,
  output [2:0]                  t8qjehupeajtzjr,
  output [3:0]                  hhp1rh0x0jn,
  output [3:0]                  w9yptl69xj6p,
  output [1-1:0]           yvcpy_gyehs4lji, 

  input                         kted7ph0krq,
  output                        a93i3d2hji,
  output [4-1:0]         of5p5cb8p4,
  output [64-1:0]       g1bi1xzuv64,
  output [8-1:0]    gj6p5b5ik3r9p,
  output                        m1fmaas4oww6,
  
  output                         hjstsi51gm,
  input                          onpqhy0s69,
  input [4-1:0]           aw7xjbi,
  input [64-1:0]         z0cc2y_uzoh_,
  input [1:0]                    y8tc_vywu82ugn,
  input                          o2h9d51o6m6,
  
  output                         nneek3ep5xykwl,
  input                          g8khua4l0y77zjp,
  input [4-1:0]           wmlp1a2b,
  input [1:0]                    weop50xb_avne,

  input                         su81e8dxdzng9d,
  input  gf33atgy,
  input  ru_wi
);

  
  localparam ale66u8k_50s8h4vdf4 = 0;
  localparam y61y499cunmtec  = 1;
  localparam a69a9ho1_kmpwc58n  = 2;
  localparam qn77zdua2lv05_ = 3;
  
  localparam gmv4r4dwujuot8a    = 4;
  localparam au8wnhbd2ozhfnnm  = 5;
  localparam s3xvyho = 6;
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  

  

  wire                         e4stso6tqp24vtt1tcak;
  wire                         m4in9wvkmutt_2mbpp4_j99;
  wire [32-1:0]   o3wrqwdzrt6so3spi3; 
  wire                         k08z5yu3rp_h5e7rub45wc; 
  wire [64-1:0]        orp433bgabdl57ym9zy;
  wire [64/8-1:0]      y1xjrtn3dgtxt18owoy6v;
  wire [2:0]                   lei05x1tdavgybso3xx;
  wire [1:0]                   anbmutawonwkdzdf7_;
  wire                         q2dp4mqsyq2hik08puc;
  wire                         zwgh_mf5sjip_yjbqbipo;
  wire [1:0]                   fg1yivrpsa618j_m0;
  wire                         kuqzfsk5p_zkwifcllye;
  wire                         osrdp3voxz5litcbd8mn;
  wire                         nccwb2tis04r3aaizdeh  ;
  wire                         wpdacu5ezxy4u9wxvnkratj6k;
  wire [64-1:0]        dqmy5amgqz8fuc8tocs;
  wire [s3xvyho-1:0]             rwkyo3nts0vnx64nmsov;

  wire [32-1:0] zys87dxafg7t5ll4o9 = 32'h0c000000;


  wire [32-1:0] rqbq0wq0_ojyw61v5 = 32'h02000000;

  
  wire                         nyz4paq9wjmwnvec_qfcu;
  wire                         fbhep995w4u17d22q277bo;
  wire [32-1:0]   g7c1mz7x6l1995sleo; 
  wire                         hl9yr8xou4foidqcxfa; 
  wire [64-1:0]        t74jedrkg_qn6tot6j;
  wire [8-1:0]     b8e707vj9boum2d0qvae2n;
  wire [2:0]                   ypyo2840fc9aou90j2mx_;
  wire [1:0]                   iicq5het5eg6ak_ss;
  wire                         zi9qv11end4ryfgzuudiby;
  wire                         u8op2__c0tfzcw0wy43d;
  wire [1:0]                   gk94omg1l9x7y_izfw08jm;
  wire                         s4f71jz9bb1u107gz7; 
  
  wire                         gy89y1sbfrskgq__rqn; 
  
  wire                         pn9ov6za1__92hofye8; 
  
  
  wire                         ug517q63iw46be392gixq23;
  wire                         y8sm4fg11fr3ofeiid4xu1;
  wire                         r43gs1mgsg15cyz3l8p    ;
  wire                         w93szs_2dzfr7cnyka2rn;
  wire [64-1:0]        us04poxovcha0t_8fnbu0f;
  
  wire                         dwy5k580q1beoesve73yleo;
  wire                         s8u4qdadsx27mgb3xyq_4gh;
  wire [32-1:0]   fc96xquw9u2s7bydi8; 
  wire                         e7e3qpjdc6ab5meyi; 
  wire [64-1:0]        dtd2nggzt96e9ofyj9;
  wire [8-1:0]     qircfy9ww3hwj431j7v;
  wire [2:0]                   xx4qeaaoc58v87c960x;
  wire [1:0]                   ixjgz15ffv3w7d9i_8;
  wire                         u62c8lyumd35ivwu4n1k7i;
  wire                         uk6jdldtxhgkfyesn5tg;
  wire [1:0]                   bd4zr8b8s4gbw7d4p3;
  wire                         a59e56gv92_za48pm1w5; 
  
  wire                         vopck74q7d_oa2f1_jf; 
  
  wire                         k2stspij_wbwj8w6pw9h; 
  
  
  wire                         mvefezow68teycp0scqosi2;
  wire                         pb1hr6cca086eg6ao3t355;
  wire                         s0l9azs15v8bj3te613_    ;
  wire                         z9a5c9cf7kiixfyz_audoq56t;
  wire [64-1:0]        utxgj9zpk_s0tosddo6aip;
  
  wire                         ecsybkzlr_tnfzkkl;
  wire                         vcecy3v4xf_qy94tzdc;
  wire [32-1:0]   eabhzanwqrvthj_rlml; 
  wire                         u4t71ko0a3pvyy0j; 
  wire [64-1:0]        y0bk8_hafbzuvphkr;
  wire [8-1:0]     p9vqll_zaxph64g51hyw;
  wire [2:0]                   cjseq5umppte3cp8f;
  wire [1:0]                   ic4lkkbrpx9ea5vfrx;
  wire                         v8u8mxxrl5epcmhaug;
  wire                         uk61v1wkskblgqzefy;
  wire [1:0]                   nxftdyjsy7jzy0k5omiy;
  wire                         jc9gu663aewk43nzkv; 
  
  wire                         jjcuvzmq_lk95jsjatz; 
  
  wire                         hdfk21faqtz079pv4; 
  
  
  wire                         qs8qyiyu8croiog92x;
  wire                         jp5kqk2q92p1i5px;
  wire                         b14z66mbuek5er6vr07    ;
  wire                         e8im2g49fb_d7x6c_5v70r;
  wire [64-1:0]        hdzpd7sew2sb4vuz;

  wire                         zd39vt7ja0cfzbczae98ls;




  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
 
  
  
  
  
  
  

  
  
  
  
  

  
  
  

  
  
  
  
  
  
  
  
  
  


  
  
  
  
  
  
  
  
  
  
  

  
  
  


  
  

  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
 
  
  
  
  
  
  
  
  
  
  

  
  
  
  
  
  
  
  
  
  
  
  
  
  


  
  localparam j5h4y56363kzi = 1;
  
  
  

  
  
  
  localparam pnbq1ed8o6an3aj = 0;
  
  localparam ubq4gj1kd8vql_2k2 = 1 + j5h4y56363kzi + pnbq1ed8o6an3aj;
  localparam v7uxeap96r379eztgx_ = (ubq4gj1kd8vql_2k2+1<=2)?1:(ubq4gj1kd8vql_2k2+1<=4)?2:(ubq4gj1kd8vql_2k2+1<=8)?3:(ubq4gj1kd8vql_2k2+1<=16)?4:(ubq4gj1kd8vql_2k2+1<=32)?5:(ubq4gj1kd8vql_2k2+1<=64)?6:(ubq4gj1kd8vql_2k2+1<=128)?7:(ubq4gj1kd8vql_2k2+1<=256)?8:(ubq4gj1kd8vql_2k2+1<=512)?9:(ubq4gj1kd8vql_2k2+1<=1024)?10:(ubq4gj1kd8vql_2k2+1<=2048)?11:(ubq4gj1kd8vql_2k2+1<=4096)?12:-1;

  localparam rqisc5uit8b_e8gzd75qx0 = 2;
  localparam n3j88a5l2ie9azx26n1g4q = 1;
  
  
  
  localparam l2u1zkau57eoz02g = 1;
  localparam cg9ef_pk_3zg7yjh_y = 1;

  
      localparam jskm09jea_69dp8a10afb = l2u1zkau57eoz02g;
  
  
  

      localparam tgongp9jmy57cyf   = jskm09jea_69dp8a10afb + 1;
      localparam qt1g9k6wsu_o7dpwq_   = cg9ef_pk_3zg7yjh_y + 1;


  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  

  wire                         b0o3_z1qhzguxuvx03v93gz;
  wire                         tslw7f9ona4tph8dm0nt;
  wire [32-1:0]   y2wr5gyopdnthewqrxe7; 
  wire                         zlz5s0ait6hwykg4b; 
  wire [64-1:0]        v2se1vid1uml27uvf2t4yli;
  wire [8-1:0]     g8ttk2wz9kvwdwkzp5kwp;
  wire [2:0]                   h4a4okoossdfjraixe2sl;
  wire [1:0]                   tnppka2a6z82_mietistn;
  wire                         tsjfjoan2dw95g05__g5q;
  wire                         hy9p1vxnb29wsf43qczd;
  wire [1:0]                   zefzgdtbg9u39vfb3;
  wire [ s3xvyho-1:0]            pds36p2k5301dpc_spd;
  wire                         hnnr5of3orcsqxyfb86ma;
  
  wire                         jl91z78pj9nm0rbl3t7www6;
  
  wire                         wjtoelq31c7h13gu_yhskwl;
  wire                         x_6hf7jugp8hwgu0j10t1;
  
  wire                         t6f_omqkgrkzy903;
  
  wire                         obdyu6w0wqx4b3g8t;
  
  wire                         yk58l7ldat5ahcp4j1i;
  wire                         e8h0j_anz7mzuobmbwzv8g;
  wire                         uebzayybqiyy1cicc  ;
  wire                         afb8snj62vkl7pacmyj3;
  wire [64-1:0]        zuv8v13fabr90783u1lc0;

  wire                         vzikn9_n0lvrdaomdo5ys;
  wire                         n1_vj412ga534kpmgnc7;
  wire [32-1:0]   ksjpl34uepyev0_db5ejr; 
  wire                         xzlaan0xyx3f5eo20zoo; 
  wire [64-1:0]        ww86vetlr_66ts64yhf00;
  wire [8-1:0]     w76w2dx5nq4zgy_xsa5;
  wire [2:0]                   l4eydle02q0gt8sp79xmpj;
  wire [1:0]                   u5iq9uuj_lmerh15q8z;
  wire                         emsvw7kp7xfm9g5s5y;
  wire                         w99a9y3nh8ju8d3ns6jr;
  wire [1:0]                   t7rgyydfts3enyenh;
  wire [ s3xvyho-1:0]            tmf4vv1fos8e5drcx985;
  wire                         iwmw44ethjx3dsud0egh;
  
  wire                         l2hjyz8uo5ft9i_3d_;
  
  wire                         ji71tydckvigh3o__p24_m;
  wire                         cugxuq_z5o_cojyelhop2;
  
  wire                         ypof75b4bl9g4e_an;
  
  
  wire                         sg96uazxf6dpizg7vad;
  wire                         qe9rerwzfqnxm49kvj69u;
  wire                         ba1jgqojkjt_p5wrx1x  ;
  wire                         jgvpcfglnc5lptyi2ca5hkmuv;
  wire [64-1:0]        xw434vczefnnjhys6_ = 64'b0;

  
  wire [s3xvyho-1:0] aefo8_8uzbuokhbce01o_f3gv;
  
  assign aefo8_8uzbuokhbce01o_f3gv[ale66u8k_50s8h4vdf4 ] = 1'b0;
  assign aefo8_8uzbuokhbce01o_f3gv[y61y499cunmtec ] = rkkjbx03o1tifh3uilzkztfkb;
  assign aefo8_8uzbuokhbce01o_f3gv[a69a9ho1_kmpwc58n ] = i0bh8gwxh68vtael53ff2y_ir5x;
  
  assign aefo8_8uzbuokhbce01o_f3gv[qn77zdua2lv05_ ] = e41m_8qgi_o4t4e2_v4c6pxn5g4;
  
  
  assign aefo8_8uzbuokhbce01o_f3gv[gmv4r4dwujuot8a   ] = ~gzq7xf16ajsco5h0qj7civq;
  assign aefo8_8uzbuokhbce01o_f3gv[au8wnhbd2ozhfnnm    ] = rpje1avuaivhahlv82bint; 
  
  
 
 
 
 
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  

  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  

  wire [s3xvyho-1:0] w_vsry_9dxmzxi82l4ixe;
  
  assign w_vsry_9dxmzxi82l4ixe[ale66u8k_50s8h4vdf4 ] = hwjq1ubtaei44lpk609fm2hb8;
  assign w_vsry_9dxmzxi82l4ixe[y61y499cunmtec ] = m04a1mtbabwezldp1crh4rg6z;
  assign w_vsry_9dxmzxi82l4ixe[a69a9ho1_kmpwc58n ] = ngyxf4n1cpcgks_s2zmgfb260;
  
  assign w_vsry_9dxmzxi82l4ixe[qn77zdua2lv05_ ] = c7m50uaw8lmp_iv4ci38q2;
  
  
  assign w_vsry_9dxmzxi82l4ixe[gmv4r4dwujuot8a   ] = 1'b0;
  assign w_vsry_9dxmzxi82l4ixe[au8wnhbd2ozhfnnm    ] = e28p_fu1k484ncul0p85ko;
 
 
 
 
 
 
  
  
  
  
  
  
  
  
  
  

  wire [s3xvyho-1:0] q2tk1oc68a_omyt1frcii1n;
  
  assign q2tk1oc68a_omyt1frcii1n[ale66u8k_50s8h4vdf4 ] = hadi1_f3quoaotjv5758x8kksot2;
  assign q2tk1oc68a_omyt1frcii1n[y61y499cunmtec ] = ju5f9fb1erjep_bv8gpfn6;
  assign q2tk1oc68a_omyt1frcii1n[a69a9ho1_kmpwc58n ] = xo6ciibewn8p8xey97jcsqi5;
  
  assign q2tk1oc68a_omyt1frcii1n[qn77zdua2lv05_ ] = evz1w_girwszyfnlcg4mwvtjo;
  
  
  assign q2tk1oc68a_omyt1frcii1n[gmv4r4dwujuot8a   ] = 1'b0;
  assign q2tk1oc68a_omyt1frcii1n[au8wnhbd2ozhfnnm    ] = bdi4gjlb0po4ejcztowoqil7;
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  wire [s3xvyho-1:0] qxad9kpc6i78vg0de9d6b;
 
  wire [s3xvyho-1:0] rfrshotpkdzarifve08g5n;
  

  wire ouat_m1vwjc0l5igzo2z4g;
  wire gyja61p9t197hw65hvyi63g;
  wire [32-1:0] v10jhardhhvft6w6t3u;
  wire mrrzsfopopzgqr_nro5;
  wire [64-1:0] pp5egelk49dgurfb3w;
  wire [8-1:0] n9sl3nl16qlprh9ocn6trcs;
  wire [2:0] g3iy6vml027o3gv9wt;
  wire [1:0] z0y5vk22vnz94pcxx;
  wire l1368lp6updfhsbebtzpc;
  wire rvqfn2hxjfeh8egdvsc;
  wire [1:0] c55olxxsckol_k4eb9fyu;
  wire [s3xvyho-1:0] jmo524gyok0abs1u1;


  wire n0wp_tjsit08gjo9ggcxe_a;
  wire ebnc6trwg85shv8_iz8qpa2;
  wire n93c2nog4f68lktvd0;
  wire uezhv2clc8f9woh7dc5ss1;
  wire [64-1:0] j2p0ug10na1wztrfj39;
  wire [s3xvyho-1:0] guqjz9gxv28q8f719;

  wire [ubq4gj1kd8vql_2k2*1-1:0] k1_j5ubhqqpfrl3p0bi186va9;
  wire [ubq4gj1kd8vql_2k2*1-1:0] w0hjg2xow0ymilw7bcxpm2l;
  wire [ubq4gj1kd8vql_2k2*32-1:0] xzpsiztjmn62eb967x1xkc6;
  wire [ubq4gj1kd8vql_2k2*1-1:0] a_dm6kd_qbw2cv84wtboltif01;
  wire [ubq4gj1kd8vql_2k2*64-1:0] ae00o9ay050qc5d5zxf18282b92;
  wire [ubq4gj1kd8vql_2k2*8-1:0] puxr8jzij0m30qcwmdz2sufl51;
  wire [ubq4gj1kd8vql_2k2*3-1:0] sxjmcdip1m7ighns0k5aue59fj;
  wire [ubq4gj1kd8vql_2k2*2-1:0] noyjdh392j1x0s9g1b_lk;
  wire [ubq4gj1kd8vql_2k2*1-1:0] s6vj39lt1yt7f1ytk3pr3;
  wire [ubq4gj1kd8vql_2k2*1-1:0] wspjbjcpf459zy17qhyz8jmqy7;
  wire [ubq4gj1kd8vql_2k2*2-1:0] y7jg1o7n3jl52fxr0isdv8;
  wire [ubq4gj1kd8vql_2k2*s3xvyho-1:0] w8o2oxw46tp1zf4rujrx4zyxw;

  wire [ubq4gj1kd8vql_2k2*1-1:0] qkiytqsa_fo9x5ls7yb_x1k2;
  wire [ubq4gj1kd8vql_2k2*1-1:0] idw2i93am7m9wy_5hzipgymj5k3;
  wire [ubq4gj1kd8vql_2k2*1-1:0] wzmdtyq65i82w_tt0juwqle;
  wire [ubq4gj1kd8vql_2k2*1-1:0] kz10yoaxkacgm38dwv37tl2ixfv;
  wire [ubq4gj1kd8vql_2k2*64-1:0] fyvkbec2dn4rlcslyiyttfrx;
  wire [ubq4gj1kd8vql_2k2*s3xvyho-1:0] od5a1yudx9bmyqpwleexh4h9;

  
  assign k1_j5ubhqqpfrl3p0bi186va9 =
      
                           {
                             
                            
                            rsgiw0g_vwk7sxen_4zrphe7,
                            
                            
                            
                            
                             swpk4h0gei3t_34xogbqncbo4
                           } ;

  
  
  

  
  wire[ubq4gj1kd8vql_2k2-1:0] ccxw7l8izxzjj14ozqkgvvyd6 =
                           {
                           
                           
                           
                           
                           
                           
                           
                           
                           
                            
                            
                            
                            
                            
                            
                            
                            rsgiw0g_vwk7sxen_4zrphe7,
                            
                            
                            
                            
                               cv0k9k_ijjnnylw1s7b_0d
                           } ;

  assign xzpsiztjmn62eb967x1xkc6 =
                           {
                             
                            
                             neuurwim9m_f3o_6nal7q7ft,
                            
                            
                            
                            
                             unu_x_i6jmr33nz0yitzk
                           } ;

  assign a_dm6kd_qbw2cv84wtboltif01 =
                           {
                             
                            
                             lpf8x_t3lmkkdri3nbex80,
                            
                            
                            
                            
                             bei3qhdtd0euq2emblogsu_x
                           } ;

  assign ae00o9ay050qc5d5zxf18282b92 =
                           {
                             
                            
                             si54q2nl6njfvmi6thon6_0,
                            
                            
                            
                            
                             bf0_ynb648lqi7s93eieo0ln
                           } ;

  assign puxr8jzij0m30qcwmdz2sufl51 =
                           {
                             
                            
                             ppe31c4mhmxn9qqmpibp3ohumo2h,
                            
                            
                            
                            
                             wf8o7p9_qfthhoxs747wyeuwkky
                           } ;
                         
  assign sxjmcdip1m7ighns0k5aue59fj =
                           {
                             
                            
                             smpikn1zm93setxcwgrzoiybl8,
                            
                            
                            
                            
                             ygro7xue7x7rtdafkj3o4q4
                           } ;
                         
  assign noyjdh392j1x0s9g1b_lk =
                           {
                             
                            
                             a6jqkrqyut1oz9lpndklbhv,
                            
                            
                            
                            
                             drrly3q0ocg8d4pwh3m9o77
                           } ;
                         
  assign s6vj39lt1yt7f1ytk3pr3 =
                           {
                             
                            
                             1'b0,
                            
                            
                            
                            
                             g654a6a9cesbee7xs6_uu9lu5
                           } ;

  assign wspjbjcpf459zy17qhyz8jmqy7 =
                           {
                             
                            
                             aum4efqs_h1yct3n53gypfa,
                            
                            
                            
                            
                             x7fex0jf9da6a5v1c28upl72t
                           } ;
                           
  assign y7jg1o7n3jl52fxr0isdv8 =
                           {
                             
                            
                             j_iw8afyzfudhp5xe0v8v231,
                            
                            
                            
                            
                             ege0_1ufqm8i68zo4il6cwe46d
                           } ;

 assign w8o2oxw46tp1zf4rujrx4zyxw =
                           {
                             
                            
                             aefo8_8uzbuokhbce01o_f3gv,
                            
                            
                            
                            
                             w_vsry_9dxmzxi82l4ixe 
                           } ;

  assign                   {
                             
                            
                             ghredfib76bt_a9caiytel4,
                            
                            
                            
                            
                             u9qmfl3rwx0dhr92z875vx7q
                           } = w0hjg2xow0ymilw7bcxpm2l;

  
  assign                   {
                             
                            
                             bygw_825g7_dt283loevm5zym41e,
                            
                            
                            
                            
                             bvg_3t_ujbpur7b_h7f63jse
                           } = qkiytqsa_fo9x5ls7yb_x1k2;

  assign                   {
                             
                            
                             c0st8ve3a3f8xhdx147o8,
                            
                            
                            
                            
                             g9so28ythfl0q7xnk66p1
                           } = wzmdtyq65i82w_tt0juwqle;
  
  
  
  
  assign                   {
                             
                            
                             wglnz1ixornvjx16dv6bvtdx6zpf,
                            
                            
                            
                            
                             e66wluxk71p2ldu3a1qk994bq
                           } = kz10yoaxkacgm38dwv37tl2ixfv;
                           
  assign                   {
                             
                            
                             h4r65p765_t877awntcuf03d6d3,
                            
                            
                            
                            
                             ig2roj0y08x8_ntp3knz9rd
                           } = fyvkbec2dn4rlcslyiyttfrx;

  assign                   {
                             
                            
                             rfrshotpkdzarifve08g5n,
                            
                            
                            
                            
                             qxad9kpc6i78vg0de9d6b 
                           } = od5a1yudx9bmyqpwleexh4h9;


  assign idw2i93am7m9wy_5hzipgymj5k3 = {
                             
                            
                             ir3fzbymkf93yhmjzi8gfgeq0,
                            
                            
                            
                            
                             m5l6wu3uz_jfqasz8e3tsvrm
                           };

  wire l0_5x2ohgu6m77k54mg;

  ux607_gnrl_icb_arbt # (
   
  .ALLOW_BURST (1),

  .ARBT_SCHEME (3),
  .FIFO_CUT_READY  (0),
  .ALLOW_0CYCL_RSP (0),
                       
  .FIFO_OUTS_NUM   (8),
  .ARBT_NUM   (ubq4gj1kd8vql_2k2),
  .ARBT_PTR_W (v7uxeap96r379eztgx_),
  .USR_W      (s3xvyho),
  .AW         (32),
  .DW         (64) 
  ) dafi4naq0de2reg2jk(
  .arbt_active            (l0_5x2ohgu6m77k54mg),
  .o_icb_cmd_valid        (ouat_m1vwjc0l5igzo2z4g )     ,
  .o_icb_cmd_ready        (gyja61p9t197hw65hvyi63g )     ,
  .o_icb_cmd_read         (mrrzsfopopzgqr_nro5 )      ,
  .o_icb_cmd_addr         (v10jhardhhvft6w6t3u )      ,
  .o_icb_cmd_wdata        (pp5egelk49dgurfb3w )     ,
  .o_icb_cmd_wmask        (n9sl3nl16qlprh9ocn6trcs)      ,
  .o_icb_cmd_burst        (g3iy6vml027o3gv9wt)     ,
  .o_icb_cmd_beat         (z0y5vk22vnz94pcxx )     ,
  .o_icb_cmd_excl         (rvqfn2hxjfeh8egdvsc )     ,
  .o_icb_cmd_lock         (l1368lp6updfhsbebtzpc )     ,
  .o_icb_cmd_size         (c55olxxsckol_k4eb9fyu )     ,
  .o_icb_cmd_usr          (jmo524gyok0abs1u1  )     ,
                                
  .o_icb_rsp_valid        (n0wp_tjsit08gjo9ggcxe_a )     ,
  .o_icb_rsp_ready        (ebnc6trwg85shv8_iz8qpa2 )     ,
  .o_icb_rsp_err          (n93c2nog4f68lktvd0)        ,
  .o_icb_rsp_excl_ok      (uezhv2clc8f9woh7dc5ss1)    ,
  .o_icb_rsp_rdata        (j2p0ug10na1wztrfj39 )     ,
  .o_icb_rsp_usr          (guqjz9gxv28q8f719)     ,
                               
  .i_bus_icb_cmd_sel_vec  (ccxw7l8izxzjj14ozqkgvvyd6) ,

  .i_bus_icb_cmd_ready    (w0hjg2xow0ymilw7bcxpm2l ) ,
  .i_bus_icb_cmd_valid    (k1_j5ubhqqpfrl3p0bi186va9 ) ,
  .i_bus_icb_cmd_read     (a_dm6kd_qbw2cv84wtboltif01 )  ,
  .i_bus_icb_cmd_addr     (xzpsiztjmn62eb967x1xkc6 )  ,
  .i_bus_icb_cmd_wdata    (ae00o9ay050qc5d5zxf18282b92 ) ,
  .i_bus_icb_cmd_wmask    (puxr8jzij0m30qcwmdz2sufl51)  ,
  .i_bus_icb_cmd_burst    (sxjmcdip1m7ighns0k5aue59fj),
  .i_bus_icb_cmd_beat     (noyjdh392j1x0s9g1b_lk ),
  .i_bus_icb_cmd_excl     (wspjbjcpf459zy17qhyz8jmqy7 ),
  .i_bus_icb_cmd_lock     (s6vj39lt1yt7f1ytk3pr3 ),
  .i_bus_icb_cmd_size     (y7jg1o7n3jl52fxr0isdv8 ),
  .i_bus_icb_cmd_usr      (w8o2oxw46tp1zf4rujrx4zyxw ),
                                
  .i_bus_icb_rsp_valid    (qkiytqsa_fo9x5ls7yb_x1k2 ) ,
  .i_bus_icb_rsp_ready    (idw2i93am7m9wy_5hzipgymj5k3 ) ,
  .i_bus_icb_rsp_err      (wzmdtyq65i82w_tt0juwqle)    ,
  .i_bus_icb_rsp_excl_ok  (kz10yoaxkacgm38dwv37tl2ixfv),
  .i_bus_icb_rsp_rdata    (fyvkbec2dn4rlcslyiyttfrx ) ,
  .i_bus_icb_rsp_usr      (od5a1yudx9bmyqpwleexh4h9) ,
                             
  .clk                    (gf33atgy  )                     ,
  .rst_n                  (ru_wi)
  );


  
  wire zprirz0krv_a3820iy7an = jmo524gyok0abs1u1[ale66u8k_50s8h4vdf4];
  wire t06t7flkpby01affnv56x64 = jmo524gyok0abs1u1[y61y499cunmtec];
  wire k8aii0cb2ywh7xvp5ud9 = jmo524gyok0abs1u1[a69a9ho1_kmpwc58n];
  
  wire vyaut44yc_lmxpxuhm = jmo524gyok0abs1u1[qn77zdua2lv05_];
  
  
  wire sedka9v4vmgj3jq44 = jmo524gyok0abs1u1[gmv4r4dwujuot8a];
  
  
  
  
  
  
  
  
  
  

  
  
  
  wire [s3xvyho-1:0] ip2id1q9t3n0hwai0_;



  
  
  
  
  
  
  
  
  assign pn9ov6za1__92hofye8 = ip2id1q9t3n0hwai0_[y61y499cunmtec];
  assign s4f71jz9bb1u107gz7 = ip2id1q9t3n0hwai0_[a69a9ho1_kmpwc58n];
  
  assign gy89y1sbfrskgq__rqn = ip2id1q9t3n0hwai0_[qn77zdua2lv05_];
  

  wire [tgongp9jmy57cyf*1-1:0] fgaj26ic3vlyw4_j9cd2e9iw5e5;
  wire [tgongp9jmy57cyf*1-1:0] fo2e9fa1xtekqy_rau1jvp;
  wire [tgongp9jmy57cyf*32-1:0] yn3_ae3lzkj5xi4qm4r12;
  wire [tgongp9jmy57cyf*1-1:0] oo66a5i9yj7eu97xzyjljzo4m;
  wire [tgongp9jmy57cyf*64-1:0] t0xc_soqbh3onidnjvuak5;
  wire [tgongp9jmy57cyf*8-1:0] hb58z51gm9p0robvubcqsio45n7;
  wire [tgongp9jmy57cyf*3-1:0] k6_7qe0217bxabwti931g5pf;
  wire [tgongp9jmy57cyf*2-1:0] mqpao8z9f30uq2rzuys2zt;
  wire [tgongp9jmy57cyf*1-1:0] j016rws5wewra_ent6uzmgq8;
  wire [tgongp9jmy57cyf*1-1:0] ubwy6_856dlynocswg3b0h3;
  wire [tgongp9jmy57cyf*2-1:0] ujjmevva2mtja2eiajfdu;
  wire [tgongp9jmy57cyf*s3xvyho-1:0] ous1ovavtg25yc9cmar2;

  wire [tgongp9jmy57cyf*1-1:0] zw0jju5nmyaae6lkudb1rc8zsh;
  wire [tgongp9jmy57cyf*1-1:0] hjab85nvos0ly5k7d5qc0a3n;
  wire [tgongp9jmy57cyf*1-1:0] eihugo5lxty1ao1uxvhn68jh;
  wire [tgongp9jmy57cyf*1-1:0] ph3072ol08mqn_adsird67uf1;
  wire [tgongp9jmy57cyf*64-1:0] qzru8eufkdrjwbh5j3iayridl0j;
  wire [tgongp9jmy57cyf*s3xvyho-1:0] zfrr8h198j86wso3hnmq6h7_; 

  
  assign {
  
  
  
                             nyz4paq9wjmwnvec_qfcu,
                             b0o3_z1qhzguxuvx03v93gz
                           } = fgaj26ic3vlyw4_j9cd2e9iw5e5;


  assign {
  
  
  
                             g7c1mz7x6l1995sleo,
                             y2wr5gyopdnthewqrxe7
                           } = yn3_ae3lzkj5xi4qm4r12;

  assign {
  
  
  
                             hl9yr8xou4foidqcxfa,
                             zlz5s0ait6hwykg4b
                           } = oo66a5i9yj7eu97xzyjljzo4m;

  assign {
  
  
  
                             t74jedrkg_qn6tot6j,
                             v2se1vid1uml27uvf2t4yli
                           } = t0xc_soqbh3onidnjvuak5;

  assign {
  
  
  
                             b8e707vj9boum2d0qvae2n,
                             g8ttk2wz9kvwdwkzp5kwp
                           } = hb58z51gm9p0robvubcqsio45n7;
                         
  assign {
  
  
  
                             ypyo2840fc9aou90j2mx_,
                             h4a4okoossdfjraixe2sl
                           } = k6_7qe0217bxabwti931g5pf;
                         
  assign {
  
  
  
                             iicq5het5eg6ak_ss,
                             tnppka2a6z82_mietistn
                           } = mqpao8z9f30uq2rzuys2zt;
                         
  assign {
  
  
  
                             zi9qv11end4ryfgzuudiby,
                             tsjfjoan2dw95g05__g5q
                           } = j016rws5wewra_ent6uzmgq8;

  assign {
  
  
  
                             u8op2__c0tfzcw0wy43d,
                             hy9p1vxnb29wsf43qczd
                           } = ubwy6_856dlynocswg3b0h3;
                           
  assign {
  
  
  
                             gk94omg1l9x7y_izfw08jm,
                             zefzgdtbg9u39vfb3
                           } = ujjmevva2mtja2eiajfdu;

  assign {
  
  
  
                             ip2id1q9t3n0hwai0_,
                             pds36p2k5301dpc_spd
                           } = ous1ovavtg25yc9cmar2;

  assign fo2e9fa1xtekqy_rau1jvp = {
  
  
  
                             fbhep995w4u17d22q277bo,
                             tslw7f9ona4tph8dm0nt
                           };

  
  assign zw0jju5nmyaae6lkudb1rc8zsh = {
  
  
  
                             ug517q63iw46be392gixq23,
                             yk58l7ldat5ahcp4j1i
                           };

  assign eihugo5lxty1ao1uxvhn68jh = {
  
  
  
                             r43gs1mgsg15cyz3l8p,
                             uebzayybqiyy1cicc
                           };

  assign ph3072ol08mqn_adsird67uf1 = {
  
  
  
                             w93szs_2dzfr7cnyka2rn,
                             afb8snj62vkl7pacmyj3
                           };

  assign qzru8eufkdrjwbh5j3iayridl0j = {
  
  
  
                             us04poxovcha0t_8fnbu0f,
                             zuv8v13fabr90783u1lc0
                           };

  assign zfrr8h198j86wso3hnmq6h7_ = {
  
  
  
                             {s3xvyho{1'b0}},
                             {s3xvyho{1'b0}}
                           };


  assign {
  
  
  
                             y8sm4fg11fr3ofeiid4xu1,
                             e8h0j_anz7mzuobmbwzv8g
                           } = hjab85nvos0ly5k7d5qc0a3n;

                           
  
  
  
  
  
  
  


  wire [32-1:0] r480zryu00zrqkrbk = 32'h00000000;
  
  
  
  wire v2xw59pj55k_pw75 = t06t7flkpby01affnv56x64 & (v10jhardhhvft6w6t3u[32-1:12] ==  r480zryu00zrqkrbk[32-1:12]);
  
  wire t4sgvg01791v9_wp720d = v2xw59pj55k_pw75 
                      
                      
                      
                      ;





  wire e8c99awftgwnivv0elc7 = 
                             (~t4sgvg01791v9_wp720d)
                      
                      
                      
                             ;

  wire [tgongp9jmy57cyf-1:0] t_xxjammw198wpina78e6g = 
      {
  
  
  
                             t4sgvg01791v9_wp720d,
                             e8c99awftgwnivv0elc7
      };

  ux607_gnrl_icb_splt # (
  
  .USE_ALL_READY(1),
  .ALLOW_DIFF (0),
  
  
  
  
  
  
  
  .VLD_MSK_PAYLOAD(0), 
  .ALLOW_0CYCL_RSP (0),
  
  
  .FIFO_OUTS_NUM   (8),
  
  
  
  
  .FIFO_CUT_READY  (0),
  
  .SPLT_NUM   (tgongp9jmy57cyf),
  .SPLT_PTR_W (tgongp9jmy57cyf),
  .SPLT_PTR_1HOT (1),
  .USR_W      (s3xvyho),
  .AW         (32),
  .DW         (64) 
  ) flgxi_8bmhbfrf1n2(
  .splt_active (),
  .i_icb_splt_indic       (t_xxjammw198wpina78e6g),        
  .i_icb_cmd_valid        (ouat_m1vwjc0l5igzo2z4g )     ,
  .i_icb_cmd_ready        (gyja61p9t197hw65hvyi63g )     ,
  .i_icb_cmd_read         (mrrzsfopopzgqr_nro5 )      ,
  .i_icb_cmd_addr         (v10jhardhhvft6w6t3u )      ,
  .i_icb_cmd_wdata        (pp5egelk49dgurfb3w )     ,
  .i_icb_cmd_wmask        (n9sl3nl16qlprh9ocn6trcs)      ,
  .i_icb_cmd_burst        (g3iy6vml027o3gv9wt)     ,
  .i_icb_cmd_beat         (z0y5vk22vnz94pcxx )     ,
  .i_icb_cmd_excl         (rvqfn2hxjfeh8egdvsc )     ,
  .i_icb_cmd_lock         (l1368lp6updfhsbebtzpc )     ,
  .i_icb_cmd_size         (c55olxxsckol_k4eb9fyu )     ,
  .i_icb_cmd_usr          (jmo524gyok0abs1u1  )     ,
 
  .i_icb_rsp_valid        (n0wp_tjsit08gjo9ggcxe_a )     ,
  .i_icb_rsp_ready        (ebnc6trwg85shv8_iz8qpa2 )     ,
  .i_icb_rsp_err          (n93c2nog4f68lktvd0)        ,
  .i_icb_rsp_excl_ok      (uezhv2clc8f9woh7dc5ss1)    ,
  .i_icb_rsp_rdata        (j2p0ug10na1wztrfj39 )     ,
  .i_icb_rsp_usr          (guqjz9gxv28q8f719)     ,
                               
  .o_bus_icb_cmd_ready    (fo2e9fa1xtekqy_rau1jvp ) ,
  .o_bus_icb_cmd_valid    (fgaj26ic3vlyw4_j9cd2e9iw5e5 ) ,
  .o_bus_icb_cmd_read     (oo66a5i9yj7eu97xzyjljzo4m )  ,
  .o_bus_icb_cmd_addr     (yn3_ae3lzkj5xi4qm4r12 )  ,
  .o_bus_icb_cmd_wdata    (t0xc_soqbh3onidnjvuak5 ) ,
  .o_bus_icb_cmd_wmask    (hb58z51gm9p0robvubcqsio45n7)  ,
  .o_bus_icb_cmd_burst    (k6_7qe0217bxabwti931g5pf),
  .o_bus_icb_cmd_beat     (mqpao8z9f30uq2rzuys2zt ),
  .o_bus_icb_cmd_excl     (ubwy6_856dlynocswg3b0h3 ),
  .o_bus_icb_cmd_lock     (j016rws5wewra_ent6uzmgq8 ),
  .o_bus_icb_cmd_size     (ujjmevva2mtja2eiajfdu ),
  .o_bus_icb_cmd_usr      (ous1ovavtg25yc9cmar2  ),
  
  .o_bus_icb_rsp_valid    (zw0jju5nmyaae6lkudb1rc8zsh ) ,
  .o_bus_icb_rsp_ready    (hjab85nvos0ly5k7d5qc0a3n ) ,
  .o_bus_icb_rsp_err      (eihugo5lxty1ao1uxvhn68jh)    ,
  .o_bus_icb_rsp_excl_ok  (ph3072ol08mqn_adsird67uf1),
  .o_bus_icb_rsp_rdata    (qzru8eufkdrjwbh5j3iayridl0j ) ,
  .o_bus_icb_rsp_usr      (zfrr8h198j86wso3hnmq6h7_) ,
                             
  .clk                    (gf33atgy  )                     ,
  .rst_n                  (ru_wi)
  );


  
  
  
  
  

  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  



  
  
  
  

  

  
  
  localparam v5m7unadv1nc4wqny = 2;
  
  wire [s3xvyho-1:0] c3xdv4h_4n95dk5x4;
  assign k2stspij_wbwj8w6pw9h = c3xdv4h_4n95dk5x4[y61y499cunmtec];
  assign a59e56gv92_za48pm1w5 = c3xdv4h_4n95dk5x4[a69a9ho1_kmpwc58n];
  
  assign vopck74q7d_oa2f1_jf = c3xdv4h_4n95dk5x4[qn77zdua2lv05_];
  

  wire [v5m7unadv1nc4wqny*1-1:0] fodcwy7kpfhsennlosy5vb3_v;
  wire [v5m7unadv1nc4wqny*1-1:0] g2yv27q_cbuwrdhyiwfpj;
  wire [v5m7unadv1nc4wqny*32-1:0] k36qftc1r5_2mw27344lonql;
  wire [v5m7unadv1nc4wqny*1-1:0] cqyc7kxwmqhl7do24px3;
  wire [v5m7unadv1nc4wqny*64-1:0] bl0xd5sad3vnmuk4xgop;
  wire [v5m7unadv1nc4wqny*8-1:0] ykwdl0lq8792mi0finz7oq;
  wire [v5m7unadv1nc4wqny*3-1:0] nu7lefdidh393nc1wou1y5;
  wire [v5m7unadv1nc4wqny*2-1:0] be9bjun1mzamdtodhfky;
  wire [v5m7unadv1nc4wqny*1-1:0] wi5zpggdjffdiphzm34;
  wire [v5m7unadv1nc4wqny*1-1:0] v_v8h1cow63gd5cineu7434;
  wire [v5m7unadv1nc4wqny*2-1:0] ityvzq_en9f5jbpyugb;
  wire [v5m7unadv1nc4wqny*s3xvyho-1:0] kllozwf7xxbetjwcty3a8ye;

  wire [qt1g9k6wsu_o7dpwq_*1-1:0] etlg6dk8qszft1po6bq_;
  wire [qt1g9k6wsu_o7dpwq_*1-1:0] i5a5h7dk65k6fx7q6_611at;
  wire [qt1g9k6wsu_o7dpwq_*1-1:0] cx3qhbal52m95qbo18c;
  wire [qt1g9k6wsu_o7dpwq_*1-1:0] cpqbmjj4innq8d21sspw80tbq;
  wire [qt1g9k6wsu_o7dpwq_*64-1:0] l5yrezudfgeh36o6jucmbgt;

  
  assign {
                             dwy5k580q1beoesve73yleo,
                             vzikn9_n0lvrdaomdo5ys
                           } = fodcwy7kpfhsennlosy5vb3_v;


  assign {
                             fc96xquw9u2s7bydi8,
                             ksjpl34uepyev0_db5ejr
                           } = k36qftc1r5_2mw27344lonql;

  assign {
                             e7e3qpjdc6ab5meyi,
                             xzlaan0xyx3f5eo20zoo
                           } = cqyc7kxwmqhl7do24px3;

  assign {
                             dtd2nggzt96e9ofyj9,
                             ww86vetlr_66ts64yhf00
                           } = bl0xd5sad3vnmuk4xgop;

  assign {
                             qircfy9ww3hwj431j7v,
                             w76w2dx5nq4zgy_xsa5
                           } = ykwdl0lq8792mi0finz7oq;
                         
  assign {
                             xx4qeaaoc58v87c960x,
                             l4eydle02q0gt8sp79xmpj
                           } = nu7lefdidh393nc1wou1y5;
                         
  assign {
                             ixjgz15ffv3w7d9i_8,
                             u5iq9uuj_lmerh15q8z
                           } = be9bjun1mzamdtodhfky;
                         
  assign {
                             u62c8lyumd35ivwu4n1k7i,
                             emsvw7kp7xfm9g5s5y
                           } = wi5zpggdjffdiphzm34;

  assign {
                             uk6jdldtxhgkfyesn5tg,
                             w99a9y3nh8ju8d3ns6jr
                           } = v_v8h1cow63gd5cineu7434;
                           
  assign {
                             bd4zr8b8s4gbw7d4p3,
                             t7rgyydfts3enyenh
                           } = ityvzq_en9f5jbpyugb;

  assign {
                             c3xdv4h_4n95dk5x4,
                             tmf4vv1fos8e5drcx985
                           } = kllozwf7xxbetjwcty3a8ye;

  assign g2yv27q_cbuwrdhyiwfpj = {
                             s8u4qdadsx27mgb3xyq_4gh,
                             n1_vj412ga534kpmgnc7
                           };

  
  assign etlg6dk8qszft1po6bq_ = {
                             mvefezow68teycp0scqosi2,
                             sg96uazxf6dpizg7vad
                           };

  assign cx3qhbal52m95qbo18c = {
                             s0l9azs15v8bj3te613_,
                             ba1jgqojkjt_p5wrx1x
                           };

  assign cpqbmjj4innq8d21sspw80tbq = {
                             z9a5c9cf7kiixfyz_audoq56t,
                             jgvpcfglnc5lptyi2ca5hkmuv
                           };

  assign l5yrezudfgeh36o6jucmbgt = {
                             utxgj9zpk_s0tosddo6aip,
                             xw434vczefnnjhys6_
                           };

  assign {
                             pb1hr6cca086eg6ao3t355,
                             qe9rerwzfqnxm49kvj69u
                           } = i5a5h7dk65k6fx7q6_611at;

  wire sin_eazp8x5b_8cxd22bl93 = ju5f9fb1erjep_bv8gpfn6 & (wn1l4cmih7rwce1rb7wk3f9wy[32-1:12] ==  r480zryu00zrqkrbk[32-1:12]);
  
  wire wf2z41kvx7gjdz8q1uxcrzd7bo = sin_eazp8x5b_8cxd22bl93;





  wire j58o4k6lwo8u6lm0avs8x59z = ~wf2z41kvx7gjdz8q1uxcrzd7bo;

  wire [qt1g9k6wsu_o7dpwq_-1:0] v9txrz0bgz_nu63bsr71y5s7in1r = 
      {
                             wf2z41kvx7gjdz8q1uxcrzd7bo,
                             j58o4k6lwo8u6lm0avs8x59z
      };

  wire l7jatybdl1tykzogmyfp36xo2x6wt;

  ux607_gnrl_icb_splt # (
  
  .USE_ALL_READY(1),
  .ALLOW_DIFF (0),
  
  
  
  
  
  
  
  .VLD_MSK_PAYLOAD(0), 
  .ALLOW_0CYCL_RSP (0),
  
  
  .FIFO_OUTS_NUM   (8),
  
  
  
  
  .FIFO_CUT_READY  (0),
  
  .SPLT_NUM   (qt1g9k6wsu_o7dpwq_),
  .SPLT_PTR_W (qt1g9k6wsu_o7dpwq_),
  .SPLT_PTR_1HOT (1),
  .USR_W      (s3xvyho),
  .AW         (32),
  .DW         (64) 
  ) dls1otq6euzvehbo8qpj_s8kwxwj(
  .splt_active            (l7jatybdl1tykzogmyfp36xo2x6wt),
  .i_icb_splt_indic       (v9txrz0bgz_nu63bsr71y5s7in1r),        

  .i_icb_cmd_valid        (twr9y24wxhs3qj2z9f2hzpaig6 )     ,
  .i_icb_cmd_ready        (w8b46r9cof57xvd5zo1u4zh8 )     ,
  .i_icb_cmd_read         (cgnzbuo_1yz6v42seb25duv )      ,
  .i_icb_cmd_addr         (wn1l4cmih7rwce1rb7wk3f9wy )      ,
  .i_icb_cmd_wdata        (zopev7f487spn9mwvuowqo )     ,
  .i_icb_cmd_wmask        (p32jk0lb8g31kqlpvmllo75qim)      ,
  .i_icb_cmd_burst        (g973rcaou05i456suvk_89dm)     ,
  .i_icb_cmd_beat         (wflv6rhfdwyxttak111v1l )     ,
  .i_icb_cmd_excl         (xu8494ii8ectqb91224uuer )     ,
  .i_icb_cmd_lock         (ggsmt4nzx8pwlowehinqvk60f )     ,
  .i_icb_cmd_size         (r6rk128ijo839ougen9stbe )     ,
  .i_icb_cmd_usr          (q2tk1oc68a_omyt1frcii1n  )     ,
 
  .i_icb_rsp_valid        (m7tq_t57mr5bovbb9ghffl4k )     ,
  .i_icb_rsp_ready        (gpcgdcri3e6_fxrw8wwtysoqqr )     ,
  .i_icb_rsp_err          (a6s4kxg1ibr6mntc85jik)        ,
  .i_icb_rsp_excl_ok      (hizzalmpwr8cqkxqi80wvbt65x)    ,
  .i_icb_rsp_rdata        ( )     ,
  .i_icb_rsp_usr          ( )     ,
                               
  .o_bus_icb_cmd_ready    (g2yv27q_cbuwrdhyiwfpj ) ,
  .o_bus_icb_cmd_valid    (fodcwy7kpfhsennlosy5vb3_v ) ,
  .o_bus_icb_cmd_read     (cqyc7kxwmqhl7do24px3 )  ,
  .o_bus_icb_cmd_addr     (k36qftc1r5_2mw27344lonql )  ,
  .o_bus_icb_cmd_wdata    (bl0xd5sad3vnmuk4xgop ) ,
  .o_bus_icb_cmd_wmask    (ykwdl0lq8792mi0finz7oq)  ,
  .o_bus_icb_cmd_burst    (nu7lefdidh393nc1wou1y5),
  .o_bus_icb_cmd_beat     (be9bjun1mzamdtodhfky ),
  .o_bus_icb_cmd_excl     (v_v8h1cow63gd5cineu7434 ),
  .o_bus_icb_cmd_lock     (wi5zpggdjffdiphzm34 ),
  .o_bus_icb_cmd_size     (ityvzq_en9f5jbpyugb ),
  .o_bus_icb_cmd_usr      (kllozwf7xxbetjwcty3a8ye  ),
  
  .o_bus_icb_rsp_valid    (etlg6dk8qszft1po6bq_ ) ,
  .o_bus_icb_rsp_ready    (i5a5h7dk65k6fx7q6_611at ) ,
  .o_bus_icb_rsp_err      (cx3qhbal52m95qbo18c)    ,
  .o_bus_icb_rsp_excl_ok  (cpqbmjj4innq8d21sspw80tbq),
  .o_bus_icb_rsp_rdata    (l5yrezudfgeh36o6jucmbgt ) ,
  .o_bus_icb_rsp_usr      ({qt1g9k6wsu_o7dpwq_*s3xvyho{1'b0}}) ,
                             
  .clk                    (gf33atgy  )                     ,
  .rst_n                  (ru_wi)
  );
  
  assign cugxuq_z5o_cojyelhop2 = tmf4vv1fos8e5drcx985[ale66u8k_50s8h4vdf4];
  assign iwmw44ethjx3dsud0egh = tmf4vv1fos8e5drcx985[a69a9ho1_kmpwc58n];
  
  assign l2hjyz8uo5ft9i_3d_ = tmf4vv1fos8e5drcx985[qn77zdua2lv05_];
  
  assign ji71tydckvigh3o__p24_m = tmf4vv1fos8e5drcx985[y61y499cunmtec];
  
  
  assign ypof75b4bl9g4e_an    = tmf4vv1fos8e5drcx985[au8wnhbd2ozhfnnm];
  

  o0kamfqxkze9obdxf3 #(
           .nm_fj (32),
           .onr7l (64),
           .h1b (8),
           .o7hawonznex2 (1),
           .n9z24gbmpt_t(8),
           .cibz (4),
           .s3xvyho (1)
) wreg2xp98wrhw8idnrf1(
           .roral7fym4h3_ (roral7fym4h3_),
           .b_gwvq35iq0_yvk (b_gwvq35iq0_yvk),
           .lqm2hm0cjm5zt (lqm2hm0cjm5zt),
           .f3n3tpjs44e0_ (f3n3tpjs44e0_),
           .dmc59hxf352z (dmc59hxf352z),
           .a63l3og_8qak5jy (a63l3og_8qak5jy),
           .m0wp58qmji79 (m0wp58qmji79),
           .c8qmnfk1vqai (c8qmnfk1vqai),
           .pbov8g9yizcwr (pbov8g9yizcwr),
           .t8qjehupeajtzjr (t8qjehupeajtzjr),
           .hhp1rh0x0jn (hhp1rh0x0jn),
           .w9yptl69xj6p (w9yptl69xj6p),
           .yvcpy_gyehs4lji (yvcpy_gyehs4lji), 
           .kted7ph0krq (kted7ph0krq),
           .a93i3d2hji (a93i3d2hji),
           .of5p5cb8p4 (of5p5cb8p4),
           .g1bi1xzuv64 (g1bi1xzuv64),
           .gj6p5b5ik3r9p (gj6p5b5ik3r9p),
           .m1fmaas4oww6 (m1fmaas4oww6),
           .nneek3ep5xykwl (nneek3ep5xykwl),
           .g8khua4l0y77zjp (g8khua4l0y77zjp),
           .wmlp1a2b (wmlp1a2b),
           .weop50xb_avne (weop50xb_avne),
           .su81e8dxdzng9d (su81e8dxdzng9d),
           .vzikn9_n0lvrdaomdo5ys (vzikn9_n0lvrdaomdo5ys),
           .n1_vj412ga534kpmgnc7 (n1_vj412ga534kpmgnc7),
           .ksjpl34uepyev0_db5ejr (ksjpl34uepyev0_db5ejr),
           .xzlaan0xyx3f5eo20zoo (xzlaan0xyx3f5eo20zoo), 
           .ww86vetlr_66ts64yhf00 (ww86vetlr_66ts64yhf00),
           .w76w2dx5nq4zgy_xsa5 (w76w2dx5nq4zgy_xsa5),
           .l4eydle02q0gt8sp79xmpj (l4eydle02q0gt8sp79xmpj),
           .u5iq9uuj_lmerh15q8z (u5iq9uuj_lmerh15q8z),
           .emsvw7kp7xfm9g5s5y (emsvw7kp7xfm9g5s5y),
           .w99a9y3nh8ju8d3ns6jr (w99a9y3nh8ju8d3ns6jr),
           .t7rgyydfts3enyenh (t7rgyydfts3enyenh),
           .iwmw44ethjx3dsud0egh (iwmw44ethjx3dsud0egh),
  
           .l2hjyz8uo5ft9i_3d_ (l2hjyz8uo5ft9i_3d_),
  
           .ji71tydckvigh3o__p24_m (ji71tydckvigh3o__p24_m),
           .cugxuq_z5o_cojyelhop2 (cugxuq_z5o_cojyelhop2),
  
           .ypof75b4bl9g4e_an (ypof75b4bl9g4e_an),
  
           .sg96uazxf6dpizg7vad (sg96uazxf6dpizg7vad),
           .qe9rerwzfqnxm49kvj69u (qe9rerwzfqnxm49kvj69u),
           .ba1jgqojkjt_p5wrx1x (ba1jgqojkjt_p5wrx1x),
           .jgvpcfglnc5lptyi2ca5hkmuv (jgvpcfglnc5lptyi2ca5hkmuv),
           .gf33atgy (gf33atgy),
           .ru_wi (ru_wi)
  );



  assign x_6hf7jugp8hwgu0j10t1 = pds36p2k5301dpc_spd[ale66u8k_50s8h4vdf4];
  assign hnnr5of3orcsqxyfb86ma = pds36p2k5301dpc_spd[a69a9ho1_kmpwc58n];
  
  assign jl91z78pj9nm0rbl3t7www6 = pds36p2k5301dpc_spd[qn77zdua2lv05_];
  
  assign wjtoelq31c7h13gu_yhskwl = pds36p2k5301dpc_spd[y61y499cunmtec];
  assign obdyu6w0wqx4b3g8t   = pds36p2k5301dpc_spd[gmv4r4dwujuot8a];
  
  
  assign t6f_omqkgrkzy903    = pds36p2k5301dpc_spd[au8wnhbd2ozhfnnm];
  

  w17x4i82vejgdgfxy6 # (
           .nm_fj (32),
           .onr7l (64),
           .h1b (8),
           .o7hawonznex2 (1),
           .cibz (4),
           .s3xvyho (1)
  ) zxmowh35i7snmkma47l(
           .wh6iy6zpdqsnv2y (wh6iy6zpdqsnv2y),
           .bd6yatp5cqq (bd6yatp5cqq),
           .fl1qsvyu (fl1qsvyu),
           .b9889wezsu (b9889wezsu),
           .an__mxugc4 (an__mxugc4),
           .poj6g8vw9e (poj6g8vw9e),
           .dafaivw3ze9g3hi (dafaivw3ze9g3hi),
           .q2c0d6fxz_1bw (q2c0d6fxz_1bw),
           .wblesminvapwua (wblesminvapwua),
           .v3cim36gj8g (v3cim36gj8g),
           .ss22f8fuy2uhr (ss22f8fuy2uhr),
           .hoaoalj5pcdnpnm0 (hoaoalj5pcdnpnm0),
           .rh8f1e3jgg3xi (rh8f1e3jgg3xi),
           .hjstsi51gm (hjstsi51gm),
           .onpqhy0s69 (onpqhy0s69),
           .aw7xjbi (aw7xjbi),
           .z0cc2y_uzoh_ (z0cc2y_uzoh_),
           .y8tc_vywu82ugn (y8tc_vywu82ugn),
           .o2h9d51o6m6 (o2h9d51o6m6),
           .su81e8dxdzng9d (su81e8dxdzng9d),
           .b0o3_z1qhzguxuvx03v93gz (b0o3_z1qhzguxuvx03v93gz),
           .tslw7f9ona4tph8dm0nt (tslw7f9ona4tph8dm0nt),
           .y2wr5gyopdnthewqrxe7 (y2wr5gyopdnthewqrxe7), 
           .zlz5s0ait6hwykg4b (zlz5s0ait6hwykg4b), 
           .v2se1vid1uml27uvf2t4yli (v2se1vid1uml27uvf2t4yli),
           .g8ttk2wz9kvwdwkzp5kwp (g8ttk2wz9kvwdwkzp5kwp),
           .h4a4okoossdfjraixe2sl (h4a4okoossdfjraixe2sl),
           .tnppka2a6z82_mietistn (tnppka2a6z82_mietistn),
           .tsjfjoan2dw95g05__g5q (tsjfjoan2dw95g05__g5q),
           .hy9p1vxnb29wsf43qczd (hy9p1vxnb29wsf43qczd),
           .zefzgdtbg9u39vfb3 (zefzgdtbg9u39vfb3),
           .hnnr5of3orcsqxyfb86ma (hnnr5of3orcsqxyfb86ma),
  
           .jl91z78pj9nm0rbl3t7www6 (jl91z78pj9nm0rbl3t7www6),
  
           .wjtoelq31c7h13gu_yhskwl (wjtoelq31c7h13gu_yhskwl),
           .x_6hf7jugp8hwgu0j10t1 (x_6hf7jugp8hwgu0j10t1),
  
           .t6f_omqkgrkzy903 (t6f_omqkgrkzy903),
  
           .obdyu6w0wqx4b3g8t (obdyu6w0wqx4b3g8t),
  
           .yk58l7ldat5ahcp4j1i (yk58l7ldat5ahcp4j1i),
           .e8h0j_anz7mzuobmbwzv8g (e8h0j_anz7mzuobmbwzv8g),
           .uebzayybqiyy1cicc   (uebzayybqiyy1cicc  ),
           .afb8snj62vkl7pacmyj3 (afb8snj62vkl7pacmyj3),
           .zuv8v13fabr90783u1lc0 (zuv8v13fabr90783u1lc0),

           .gf33atgy (gf33atgy),
           .ru_wi (ru_wi)
  );



  localparam k028vzf3ra7ssohjrbrh = 2;

  wire [rqisc5uit8b_e8gzd75qx0*1-1:0] l5tsab0sqo0n_d6ievr89wvmov9;
  wire [rqisc5uit8b_e8gzd75qx0*1-1:0] d3wf7rqyp28k808_4yv2amqx8;
  wire [rqisc5uit8b_e8gzd75qx0*32-1:0] fz_9jjmrwbl0x0jq3w84ctqg;
  wire [rqisc5uit8b_e8gzd75qx0*1-1:0] ltveuvdp6nss7h1qrdxlo_4t5unaq;
  wire [rqisc5uit8b_e8gzd75qx0*64-1:0] jxzssxptuxnifssmw57euftkk;
  wire [rqisc5uit8b_e8gzd75qx0*8-1:0] vo0co_zh4gjy1gqlsdset7qlfvham;
  wire [rqisc5uit8b_e8gzd75qx0*3-1:0] huf3f8zo1ujvtytk_hlqbgrcd3rej;
  wire [rqisc5uit8b_e8gzd75qx0*2-1:0] ods0tis9x5o8n44srbyjk_9y;
  wire [rqisc5uit8b_e8gzd75qx0*1-1:0] l456ch0bikniun5fije181vc;
  wire [rqisc5uit8b_e8gzd75qx0*1-1:0] mos8c7gufts5jnylgq0osbefd5br;
  wire [rqisc5uit8b_e8gzd75qx0*2-1:0] v7mdx55sudzukvuitqbprtfi46g;
  wire [rqisc5uit8b_e8gzd75qx0*s3xvyho-1:0] pt66m5chwm0kco8rilh685td89c;

  wire [rqisc5uit8b_e8gzd75qx0*1-1:0] e64l534duvjvnh5mxnhe_re0k;
  wire [rqisc5uit8b_e8gzd75qx0*1-1:0] vjlqqk6gu_7cb0swk5uw_wane50q;
  wire [rqisc5uit8b_e8gzd75qx0*1-1:0] j24k7uyfmdr4t08h73d612374swq;
  wire [rqisc5uit8b_e8gzd75qx0*1-1:0] ai5c6dtwzv4u_jfexv40c5vb9uj;
  wire [rqisc5uit8b_e8gzd75qx0*64-1:0] ojevdg64xndfmxteurf43mdtln;

  wire [1-1:0] jt8c9rjwkn8lcqqhng9_0rkwzm;
  wire [1-1:0] z97xlmd_06lshqp4qpvdjjk9;
  wire [32-1:0] ys9svkgs7ehid3g6v2nmh_ewvzhj;
  wire [1-1:0] mdj3azutscdsl_jw_6rdo8w2;
  wire [64-1:0] me9_l0p1q9qgf3ksjd8gq5o6jiwlz;
  wire [8-1:0] h4q40ks30q_za7zfiq_dz2woq;
  wire [3-1:0] q2xi1lc6v9ihg5hmkmuxzhwn2;
  wire [2-1:0] p833vj11pxzwjlafweeowfh0c3u;
  wire [1-1:0] l54mdbe69nlx2rmysv1m3r48r;
  wire [1-1:0] n_ikxrtrrqgzmailkj5ebe0ky8;
  wire [2-1:0] zi9k2d9ah3o0g79me87i6_w;
  wire [s3xvyho-1:0] fu2buyqapzdehjfqjdg6nkx;

  wire [1-1:0] nau9wwz7sajptf6pn7jcib_8of;
  wire [1-1:0] gh3kwcfv8zoqnorfvfqk8akktqan;
  wire [1-1:0] q75njoov56n858zcf65rbo87qnr;
  wire [1-1:0] r7mnoinehf9ok5bazlrk7r8x3cgwby;
  wire [64-1:0] nt9i8ly88u0w48tbbfculm_akruf;

  wire                        twj6lwlfjeszrahzsibq59;

  wire [s3xvyho-1:0] o9vfhezgtb2rfa3fn;
  assign hdfk21faqtz079pv4 = o9vfhezgtb2rfa3fn[y61y499cunmtec];
  assign jc9gu663aewk43nzkv = o9vfhezgtb2rfa3fn[a69a9ho1_kmpwc58n];
  
  assign jjcuvzmq_lk95jsjatz = o9vfhezgtb2rfa3fn[qn77zdua2lv05_];
  


  
  
  
  
  
  
  wire b7a3c8f0ucgrh1pe44;
  wire anzgxl3b1fzrx156hfmje;
  
  
  
  
  
  
  
  
  
  
  
  assign b7a3c8f0ucgrh1pe44 = ~dwy5k580q1beoesve73yleo;
  assign anzgxl3b1fzrx156hfmje =  dwy5k580q1beoesve73yleo;
  
  
  

  
  assign l5tsab0sqo0n_d6ievr89wvmov9 =
      
                           {
                             nyz4paq9wjmwnvec_qfcu,
                             dwy5k580q1beoesve73yleo
                           } ;

  wire[rqisc5uit8b_e8gzd75qx0-1:0] y7bjqwl6wgs3ob8uzdu98lsgf308_n2 =
                           {
                               b7a3c8f0ucgrh1pe44 
                             , anzgxl3b1fzrx156hfmje
                           } ;

  assign fz_9jjmrwbl0x0jq3w84ctqg =
                           {
                             g7c1mz7x6l1995sleo,
                             fc96xquw9u2s7bydi8
                           } ;

  assign ltveuvdp6nss7h1qrdxlo_4t5unaq =
                           {
                             hl9yr8xou4foidqcxfa,
                             e7e3qpjdc6ab5meyi
                           } ;

  assign jxzssxptuxnifssmw57euftkk =
                           {
                             t74jedrkg_qn6tot6j,
                             dtd2nggzt96e9ofyj9
                           } ;

  assign vo0co_zh4gjy1gqlsdset7qlfvham =
                           {
                             b8e707vj9boum2d0qvae2n,
                             qircfy9ww3hwj431j7v
                           } ;
                         
  assign huf3f8zo1ujvtytk_hlqbgrcd3rej =
                           {
                             ypyo2840fc9aou90j2mx_,
                             xx4qeaaoc58v87c960x
                           } ;
                         
  assign ods0tis9x5o8n44srbyjk_9y =
                           {
                             iicq5het5eg6ak_ss,
                             ixjgz15ffv3w7d9i_8
                           } ;
                         
  assign l456ch0bikniun5fije181vc =
                           {
                             1'b0,
                             1'b0 
                           } ;

  assign mos8c7gufts5jnylgq0osbefd5br =
                           {
                             u8op2__c0tfzcw0wy43d,
                             uk6jdldtxhgkfyesn5tg
                           } ;
                           
  assign v7mdx55sudzukvuitqbprtfi46g =
                           {
                             gk94omg1l9x7y_izfw08jm,
                             bd4zr8b8s4gbw7d4p3
                           } ;

 assign pt66m5chwm0kco8rilh685td89c =
                           {
                             ip2id1q9t3n0hwai0_,
                             c3xdv4h_4n95dk5x4 
                           } ;

  assign                   {
                             fbhep995w4u17d22q277bo,
                             s8u4qdadsx27mgb3xyq_4gh
                           } = d3wf7rqyp28k808_4yv2amqx8;

  
  assign                   {
                             ug517q63iw46be392gixq23,
                             mvefezow68teycp0scqosi2
                           } = e64l534duvjvnh5mxnhe_re0k;

  assign                   {
                             r43gs1mgsg15cyz3l8p,
                             s0l9azs15v8bj3te613_
                           } = j24k7uyfmdr4t08h73d612374swq;

  assign                   {
                             w93szs_2dzfr7cnyka2rn,
                             z9a5c9cf7kiixfyz_audoq56t
                           } = ai5c6dtwzv4u_jfexv40c5vb9uj;
                           
  assign                   {
                             us04poxovcha0t_8fnbu0f,
                             utxgj9zpk_s0tosddo6aip
                           } = ojevdg64xndfmxteurf43mdtln;

  assign vjlqqk6gu_7cb0swk5uw_wane50q = {
                             y8sm4fg11fr3ofeiid4xu1,
                             pb1hr6cca086eg6ao3t355
                           };


  ux607_gnrl_icb_arbt # (
   
  .ALLOW_BURST (1),

  .ARBT_SCHEME (3),
  
  .FIFO_CUT_READY  (0),
  .ALLOW_0CYCL_RSP (0),
                       
  .FIFO_OUTS_NUM   (8),
  .ARBT_NUM   (rqisc5uit8b_e8gzd75qx0),
  .ARBT_PTR_W (n3j88a5l2ie9azx26n1g4q),
  .USR_W      (s3xvyho),
  .AW         (32),
  .DW         (64) 
  ) bwxarlys2b6g88zf(
  .arbt_active            (zd39vt7ja0cfzbczae98ls),
  .o_icb_cmd_valid        (jt8c9rjwkn8lcqqhng9_0rkwzm )     ,
  .o_icb_cmd_ready        (z97xlmd_06lshqp4qpvdjjk9 )     ,
  .o_icb_cmd_read         (mdj3azutscdsl_jw_6rdo8w2 )      ,
  .o_icb_cmd_addr         (ys9svkgs7ehid3g6v2nmh_ewvzhj )      ,
  .o_icb_cmd_wdata        (me9_l0p1q9qgf3ksjd8gq5o6jiwlz )     ,
  .o_icb_cmd_wmask        (h4q40ks30q_za7zfiq_dz2woq)      ,
  .o_icb_cmd_burst        (q2xi1lc6v9ihg5hmkmuxzhwn2)     ,
  .o_icb_cmd_beat         (p833vj11pxzwjlafweeowfh0c3u )     ,
  .o_icb_cmd_excl         (n_ikxrtrrqgzmailkj5ebe0ky8 )     ,
  .o_icb_cmd_lock         (l54mdbe69nlx2rmysv1m3r48r )     ,
  .o_icb_cmd_size         (zi9k2d9ah3o0g79me87i6_w )     ,
  .o_icb_cmd_usr          (fu2buyqapzdehjfqjdg6nkx  )     ,
                                      
  .o_icb_rsp_valid        (nau9wwz7sajptf6pn7jcib_8of )     ,
  .o_icb_rsp_ready        (gh3kwcfv8zoqnorfvfqk8akktqan )     ,
  .o_icb_rsp_err          (q75njoov56n858zcf65rbo87qnr)        ,
  .o_icb_rsp_excl_ok      (r7mnoinehf9ok5bazlrk7r8x3cgwby)    ,
  .o_icb_rsp_rdata        (nt9i8ly88u0w48tbbfculm_akruf )     ,
  .o_icb_rsp_usr          ({s3xvyho{1'b0}}   )     ,
                               
  .i_bus_icb_cmd_sel_vec  (y7bjqwl6wgs3ob8uzdu98lsgf308_n2) ,

  .i_bus_icb_cmd_ready    (d3wf7rqyp28k808_4yv2amqx8 ) ,
  .i_bus_icb_cmd_valid    (l5tsab0sqo0n_d6ievr89wvmov9 ) ,
  .i_bus_icb_cmd_read     (ltveuvdp6nss7h1qrdxlo_4t5unaq )  ,
  .i_bus_icb_cmd_addr     (fz_9jjmrwbl0x0jq3w84ctqg )  ,
  .i_bus_icb_cmd_wdata    (jxzssxptuxnifssmw57euftkk ) ,
  .i_bus_icb_cmd_wmask    (vo0co_zh4gjy1gqlsdset7qlfvham)  ,
  .i_bus_icb_cmd_burst    (huf3f8zo1ujvtytk_hlqbgrcd3rej),
  .i_bus_icb_cmd_beat     (ods0tis9x5o8n44srbyjk_9y ),
  .i_bus_icb_cmd_excl     (mos8c7gufts5jnylgq0osbefd5br ),
  .i_bus_icb_cmd_lock     (l456ch0bikniun5fije181vc ),
  .i_bus_icb_cmd_size     (v7mdx55sudzukvuitqbprtfi46g ),
  .i_bus_icb_cmd_usr      (pt66m5chwm0kco8rilh685td89c ),
                         
  .i_bus_icb_rsp_valid    (e64l534duvjvnh5mxnhe_re0k ) ,
  .i_bus_icb_rsp_ready    (vjlqqk6gu_7cb0swk5uw_wane50q ) ,
  .i_bus_icb_rsp_err      (j24k7uyfmdr4t08h73d612374swq)    ,
  .i_bus_icb_rsp_excl_ok  (ai5c6dtwzv4u_jfexv40c5vb9uj),
  .i_bus_icb_rsp_rdata    (ojevdg64xndfmxteurf43mdtln ) ,
  .i_bus_icb_rsp_usr      () ,
                             
  .clk                    (gf33atgy  )                     ,
  .rst_n                  (ru_wi)
  );

  ux607_gnrl_icb_buffer # (
    .OUTS_CNT_W   (4),
    .AW    (32),
    .DW    (64), 

    .CMD_MSKO(0),

    .CMD_DP(2),
    .RSP_DP(2),
      
      
      
    .RSP_ALWAYS_READY (1),
      
      
      
    .CMD_CUT_READY (1),
    .RSP_CUT_READY (1),
    .USR_W (s3xvyho)
  )v7pkxitoqbhkeuctz76pf(
    .bus_clk_en             (1'b1),

    .icb_buffer_active      (twj6lwlfjeszrahzsibq59),
    .i_icb_cmd_valid        (jt8c9rjwkn8lcqqhng9_0rkwzm),
    .i_icb_cmd_ready        (z97xlmd_06lshqp4qpvdjjk9),
    .i_icb_cmd_read         (mdj3azutscdsl_jw_6rdo8w2 ),
    .i_icb_cmd_addr         (ys9svkgs7ehid3g6v2nmh_ewvzhj ),
    .i_icb_cmd_wdata        (me9_l0p1q9qgf3ksjd8gq5o6jiwlz),
    .i_icb_cmd_wmask        (h4q40ks30q_za7zfiq_dz2woq),
    .i_icb_cmd_lock         (l54mdbe69nlx2rmysv1m3r48r ),
    .i_icb_cmd_excl         (n_ikxrtrrqgzmailkj5ebe0ky8 ),
    .i_icb_cmd_size         (zi9k2d9ah3o0g79me87i6_w ),
    .i_icb_cmd_burst        (q2xi1lc6v9ihg5hmkmuxzhwn2),
    .i_icb_cmd_beat         (p833vj11pxzwjlafweeowfh0c3u ),
    .i_icb_cmd_usr          (fu2buyqapzdehjfqjdg6nkx  ),
                     
    .i_icb_rsp_valid        (nau9wwz7sajptf6pn7jcib_8of),
    .i_icb_rsp_ready        (gh3kwcfv8zoqnorfvfqk8akktqan),
    .i_icb_rsp_err          (q75njoov56n858zcf65rbo87qnr  ),
    .i_icb_rsp_excl_ok      (r7mnoinehf9ok5bazlrk7r8x3cgwby),
    .i_icb_rsp_rdata        (nt9i8ly88u0w48tbbfculm_akruf),
    .i_icb_rsp_usr          (),
    
    .o_icb_cmd_valid        (e4stso6tqp24vtt1tcak),
    .o_icb_cmd_ready        (m4in9wvkmutt_2mbpp4_j99),
    .o_icb_cmd_read         (k08z5yu3rp_h5e7rub45wc ),
    .o_icb_cmd_addr         (o3wrqwdzrt6so3spi3 ),
    .o_icb_cmd_wdata        (orp433bgabdl57ym9zy),
    .o_icb_cmd_wmask        (y1xjrtn3dgtxt18owoy6v),
    .o_icb_cmd_lock         (q2dp4mqsyq2hik08puc ),
    .o_icb_cmd_excl         (zwgh_mf5sjip_yjbqbipo ),
    .o_icb_cmd_size         (fg1yivrpsa618j_m0 ),
    .o_icb_cmd_burst        (lei05x1tdavgybso3xx),
    .o_icb_cmd_beat         (anbmutawonwkdzdf7_ ),
    .o_icb_cmd_usr          (rwkyo3nts0vnx64nmsov),
                         
    .o_icb_rsp_valid        (kuqzfsk5p_zkwifcllye),
    .o_icb_rsp_ready        (osrdp3voxz5litcbd8mn),
    .o_icb_rsp_err          (nccwb2tis04r3aaizdeh  ),
    .o_icb_rsp_excl_ok      (wpdacu5ezxy4u9wxvnkratj6k),
    .o_icb_rsp_rdata        (dqmy5amgqz8fuc8tocs),
    .o_icb_rsp_usr          ({s3xvyho{1'b0}}  ),

    .clk                    (gf33atgy  ),
    .rst_n                  (ru_wi)
  );

 ux607_gnrl_icb2ahbl
  #(
      .SUPPORT_LOCK     (0),
      .AW(32),
      .MON_DATA_WIDTH(3),
      .DW(64) 
    ) jrk8__gbwyk5p(
    .icb2ahbl_pend_active(),
    .bus_clk_en        (1'b1),
    .icb_cmd_valid     (ecsybkzlr_tnfzkkl),  
    .icb_cmd_ready     (vcecy3v4xf_qy94tzdc),  
    .icb_cmd_read      (u4t71ko0a3pvyy0j ), 
    .icb_cmd_addr      (eabhzanwqrvthj_rlml ), 
    .icb_cmd_wdata     (y0bk8_hafbzuvphkr),  
    .icb_cmd_wmask     (8'b0), 
    .icb_cmd_size      (nxftdyjsy7jzy0k5omiy ),
    .icb_cmd_lock      (1'b0 ),
    .icb_cmd_excl      (1'b0 ),
    .icb_cmd_burst     (3'b0),  
    .icb_cmd_hseq      (1'b0 ), 
    .icb_cmd_hprot     (4'b0), 
    .icb_cmd_attri     (2'b0), 
    .icb_cmd_dmode     (1'b0), 
                       
    .icb_rsp_valid     (qs8qyiyu8croiog92x),  
    
    .icb_rsp_err       (b14z66mbuek5er6vr07    ),
    .icb_rsp_excl_ok   (e8im2g49fb_d7x6c_5v70r),
    .icb_rsp_rdata     (hdzpd7sew2sb4vuz),  
                      
    .ahbl_htrans       (pszbl2iobld50k  ),  
    .ahbl_hwrite       (vfuu2l_7oof31qn0_a  ),  
    .ahbl_haddr        (bvy9o58rgxtbjz_xph   ),  
    .ahbl_hsize        (gcpthp2sfxb3cxo   ),  
    .ahbl_hlock        (), 
    .ahbl_hexcl        (), 
    .ahbl_hburst       (xzjdk5deciqs4l3my_l),  
    .ahbl_hwdata       (dlg9f36umgj9xdv0wa  ),  
    .ahbl_hprot        (peug05ptx4vv93u4xc),
    .ahbl_hattri       (),
    .ahbl_master       (),
    .ahbl_hrdata       (yienty7ycnc25au  ),  
    .ahbl_hresp        (rxlx2eq69oye0ba3   ),  
    .ahbl_hresp_exok   (1'b0   ),  
    .ahbl_hready       (j2amhrzbhku8dzd  ),  
       
    .clk               (gf33atgy),
    .rst_n             (ru_wi)
  );

  
  wire oedsjse0mgifw4;
  wire xrmzcyhiwrtffg2 = ecsybkzlr_tnfzkkl & vcecy3v4xf_qy94tzdc;
  wire jmjp6v54e5w5 = qs8qyiyu8croiog92x & jp5kqk2q92p1i5px;
     
  wire h8xkmf95fhew = xrmzcyhiwrtffg2 | jmjp6v54e5w5;
  wire l8leuuwqvb147 = xrmzcyhiwrtffg2 | (~jmjp6v54e5w5);
     
  ux607_gnrl_dfflr #(1) ujp_o3_9pbnnlfl8 (h8xkmf95fhew, l8leuuwqvb147, oedsjse0mgifw4, gf33atgy, ru_wi);

  assign wex3zbl1x6s4be1en = ecsybkzlr_tnfzkkl | oedsjse0mgifw4;


  assign nv5a7f_68p9ebw = 
                      l0_5x2ohgu6m77k54mg |
                      l7jatybdl1tykzogmyfp36xo2x6wt |
                      
                      
                      swpk4h0gei3t_34xogbqncbo4 |
                      rsgiw0g_vwk7sxen_4zrphe7 | 
                    
                    
                    
                      twr9y24wxhs3qj2z9f2hzpaig6 |
                      zd39vt7ja0cfzbczae98ls |
                      twj6lwlfjeszrahzsibq59 | 
                      wex3zbl1x6s4be1en |
                      1'b0;

  
  
     assign ecsybkzlr_tnfzkkl   = e4stso6tqp24vtt1tcak;
     assign m4in9wvkmutt_2mbpp4_j99   = vcecy3v4xf_qy94tzdc;
     assign eabhzanwqrvthj_rlml    = o3wrqwdzrt6so3spi3 ; 
     assign u4t71ko0a3pvyy0j    = k08z5yu3rp_h5e7rub45wc ; 
     assign cjseq5umppte3cp8f   = lei05x1tdavgybso3xx;
     assign ic4lkkbrpx9ea5vfrx    = anbmutawonwkdzdf7_ ;
     assign y0bk8_hafbzuvphkr   = orp433bgabdl57ym9zy;
     assign p9vqll_zaxph64g51hyw   = y1xjrtn3dgtxt18owoy6v;
     assign v8u8mxxrl5epcmhaug    = q2dp4mqsyq2hik08puc ;
     assign uk61v1wkskblgqzefy    = zwgh_mf5sjip_yjbqbipo ;
     assign nxftdyjsy7jzy0k5omiy    = fg1yivrpsa618j_m0 ;
     assign o9vfhezgtb2rfa3fn     = rwkyo3nts0vnx64nmsov  ;

     assign kuqzfsk5p_zkwifcllye   = qs8qyiyu8croiog92x  ;
     assign jp5kqk2q92p1i5px   = osrdp3voxz5litcbd8mn  ;
     assign nccwb2tis04r3aaizdeh     = b14z66mbuek5er6vr07    ;
     assign wpdacu5ezxy4u9wxvnkratj6k = e8im2g49fb_d7x6c_5v70r;
     assign dqmy5amgqz8fuc8tocs   = hdzpd7sew2sb4vuz;

endmodule



















module fp3ou97fzh9for8cue9y6 #(
    parameter iu_89 = 1,
    parameter m_rz39tx6bnugdx = 5
)(
    input  gf33atgy,
    input  ru_wi,
    input  dbcjt09pmjkdprn,
    input  [1:0] gsy4z_7std_ruja54_37j,
    input  jjt5ro1ekg7v7uhoesn8f,
    input  [m_rz39tx6bnugdx-1:0] kg87hyc2ic61h2q6wd7j5sb,
    input  e8cte26q6yj870i027qa9r62,
    input  fz_isl8q3blzlbl2zzf,
    input  [31:0] u4r4b_6kp09q767q,
    output k4xratl2pp6xdh98,
    output [7:0] oyzrjkmgclshj
);

wire dgrt7jaaqbkmr;
wire jxx7cnp3_0sh11li0b;
ux607_gnrl_dffr #(1) v_n23_acr8pmljtt7k(dbcjt09pmjkdprn,dgrt7jaaqbkmr,gf33atgy,ru_wi);

wire l8jr4q_z1fsrcuv_r6s = dbcjt09pmjkdprn & (~dgrt7jaaqbkmr);
wire b_1jcordsdhwqke6ra9= (~dbcjt09pmjkdprn) & dgrt7jaaqbkmr;

wire wcw_oy9ki2pngt = e8cte26q6yj870i027qa9r62 & fz_isl8q3blzlbl2zzf;  

wire e91yshw3o6bm821q = (~oyzrjkmgclshj[0]) & (gsy4z_7std_ruja54_37j[0]) & (gsy4z_7std_ruja54_37j[1] ? b_1jcordsdhwqke6ra9 :
                                                                l8jr4q_z1fsrcuv_r6s);
wire b60s8pkxd278437s = jjt5ro1ekg7v7uhoesn8f & (gsy4z_7std_ruja54_37j[0]) & (kg87hyc2ic61h2q6wd7j5sb == iu_89[m_rz39tx6bnugdx-1:0]);
wire y955ssw8d8eq36g9gzyotci;

assign jxx7cnp3_0sh11li0b = wcw_oy9ki2pngt ? u4r4b_6kp09q767q[0] :
                       e91yshw3o6bm821q ? 1'b1 : 
                       b60s8pkxd278437s ? 1'b0 : 
                       y955ssw8d8eq36g9gzyotci;
                                      

wire otf3fj4j68p0341e3z = wcw_oy9ki2pngt | e91yshw3o6bm821q | b60s8pkxd278437s;
ux607_gnrl_dfflr #(1) mn5zo5tj711wu_h_xqz7k(otf3fj4j68p0341e3z, jxx7cnp3_0sh11li0b, y955ssw8d8eq36g9gzyotci, gf33atgy, ru_wi);

assign oyzrjkmgclshj = gsy4z_7std_ruja54_37j[0] ? {7'b0,y955ssw8d8eq36g9gzyotci} : {7'b0,dgrt7jaaqbkmr};





wire g4olr45r_y646l5p1ktc0t = (~gsy4z_7std_ruja54_37j[0]);
wire js0kp8sisse2zl1iw67egjh = gsy4z_7std_ruja54_37j[0] &  (~gsy4z_7std_ruja54_37j[1]);
wire t2jm3oogurogf42rtyuc598sbks = gsy4z_7std_ruja54_37j[0] &  gsy4z_7std_ruja54_37j[1];
assign k4xratl2pp6xdh98 = (dbcjt09pmjkdprn & (g4olr45r_y646l5p1ktc0t |  js0kp8sisse2zl1iw67egjh)) 
                    | ((~dbcjt09pmjkdprn) & t2jm3oogurogf42rtyuc598sbks)
                    ;

endmodule



















module d2x3825_dhbv0h # (
    parameter vb1dh27fsxbyysw = 32,
    parameter t5twosugmt3qlv = 5
)(
    input   dk2xhkj77a,
    input   gf33atgy,
    input   zh6e0v0mmz,
    input   ru_wi,
    
    input                           a3v1iy5k0,
    input                           cjwv,

    input [vb1dh27fsxbyysw-20:0]       fcjh1nct4r,

    input                           th06du2c8e2_b7k,
    output                          irjoi8wvo25u209f_5,
    input  [16-1:0]                 zvk11dhgg2s67mkq,
    input  [4-1:0]                  lhibcc3xwm6cy,
    input                           zxe59xihintdqfy9d,
    input  [31:0]                   u4r4b_6kp09q767q,

    output                          klkflmsyyf5w7ar,
    input                           wy36iirxspfw56864,
    output [31:0]                   h7f6k_ims_9p3,
    output                          lkjqs6kiuyj,

    input                           dz0zrf512290tvcy4q,
    input                           gfy3zost37aq8qmr,
    input                           dn8riluj40uunvq5,
    input                           dxi_ue3gf5zqqqxwgq2a,
    input                           aw82i964do,
    input                           fbzs0o4ysyuzeg_qdj,
    input                           me1n4pvwxa7n3u8l05,
    input                           qaidts35dk5jcji0n,
    input                           y8_gkxsfle,
    input                           fzdb65fcrotwcaccus_cwo,
    input [7:0]                     tcy_87vt9vet39knuw,
    output                          fc_4ns_w1nh4h02z_dgg,
    output                          jqsukc5b5drcc1e78,
    output                          gnn46rd7vvofruqij,

    output                          y12wg4mlovhn13,
    output                          kfrxhvr3mwznw,
    output [9:0]                    b4lwcgm6l21pi,
    output                          zwcbp7zqfei5xz,
    input [7:0]                     f_i1959b4xizzq9jea,
    output [7:0]                    hjrk_rwjkqj3zk_b, 
    output                          znzjygllppv1s0a8cqub3c
);

 
    localparam lhc8m69xvstkozu5iz8i4 = (vb1dh27fsxbyysw<=2)?1:(vb1dh27fsxbyysw<=4)?2:(vb1dh27fsxbyysw<=8)?3:(vb1dh27fsxbyysw<=16)?4:(vb1dh27fsxbyysw<=32)?5:(vb1dh27fsxbyysw<=64)?6:(vb1dh27fsxbyysw<=128)?7:(vb1dh27fsxbyysw<=256)?8:(vb1dh27fsxbyysw<=512)?9:(vb1dh27fsxbyysw<=1024)?10:(vb1dh27fsxbyysw<=2048)?11:(vb1dh27fsxbyysw<=4096)?12:-1;
    localparam ujp_32rzn = 1; 

    wire h5maomnmovgqtb7 = th06du2c8e2_b7k & irjoi8wvo25u209f_5;
    wire fz_isl8q3blzlbl2zzf = h5maomnmovgqtb7 & (~zxe59xihintdqfy9d);
    wire dh1lon9y8avka453f7vc = h5maomnmovgqtb7 & zxe59xihintdqfy9d;

    wire                                e6e9h0kbbxy00yvvbp0bywk;
    wire                                dc0ovps7up6g7sxmwjd4;
    wire                                sgyw532glkiyqyuycg_ymn;
    wire                                hzql4_1_2nrk6cp7kzhr9mz0;

    wire [vb1dh27fsxbyysw-1:0]             e8cte26q6yj870i027qa9r62;
    wire [vb1dh27fsxbyysw-1:0]             w0nv2a98k9wdk7ddkoo6wuf5;
    wire [vb1dh27fsxbyysw-1:0]             bloeijx3qz0wz5u_avwjaa2we;
    wire [vb1dh27fsxbyysw-1:0]             u0xuahg9aulem6ytjre5dm;

    wire [vb1dh27fsxbyysw-1:0]             f63dz5dw05rfd8s39jwx1s_5;
    wire [vb1dh27fsxbyysw-1:0]             enu9bknh9ueizhtexpv7ggo9qoggsu;

    wire                                mzp5pkv6xl9_nmhw;
    wire                                c5a84c6g_dbse_yvi61emns; 
    wire                                ij34sjy812rgbeddhqm0ts; 
    wire [vb1dh27fsxbyysw-1:0]             dcs94jjnvo_oqe_;
    wire [vb1dh27fsxbyysw-1:0]             q9dddg5qvq6azwmv5;
    wire [vb1dh27fsxbyysw-1:0]             sc9i3oongjhvjssm8b;

    wire [7:0]                          bqe4lf3omz8wflk3ncm1d;
    wire [7:0]                          ij93945qy0t4clwq0b;
    wire [7:0]                          a7wgjswsdhh5p;
    wire [7:0]                          wvmr61jza7zhd5o0u[0:vb1dh27fsxbyysw-1];
    wire [7:0]                          mglzjmd3n4ynn8[0:vb1dh27fsxbyysw-1];
    wire [7:0]                          mysay5szii2i_ucs[0:vb1dh27fsxbyysw-1];
    wire [31:0]                         lva2sw2f_nq_1u5780; 
    wire [31:0]                         l05bm7_xtgbitxwsk_3; 
    wire [31:0]                         w5t0kiz2tj15hher468m_ngc; 
    wire [31:0]                         hkmb5i4b7onky8b45mmb4l6y; 
    reg [31:0]                          isd23fnq13pcssxpxiacb;


    wire [7:0]                          ufx6dsiuus18;
    wire [3:0]                          oi2196y9j6yk8xp9 = ufx6dsiuus18[4:1];

    wire [7:0]                          bpkwqkepwyytmwn1;
    wire [7:0]                          uauce93oo4hzcipngfgg;
    wire [vb1dh27fsxbyysw-1:0]             k4xratl2pp6xdh98;
    wire [7:0]                          oyzrjkmgclshj[0:vb1dh27fsxbyysw-1];
    wire [7:0]                          qhzxh33vz7eo6[0:vb1dh27fsxbyysw-1];
    wire [7:0]                          q_8115sz8oh72wnv9[0:vb1dh27fsxbyysw-1];
    wire [vb1dh27fsxbyysw-1:0]             tbf0wzltxdlu9ouilvocb_f62;
    wire [vb1dh27fsxbyysw-1:0]             l6hr3z_7lt62kdb3uv;
    wire                                x3g5a2s4f40otq82g[0:vb1dh27fsxbyysw-1];
    wire [7:0]                          z1gysizgxf7x[0:vb1dh27fsxbyysw-1];
    
    wire [t5twosugmt3qlv+1:0]           cs8o9yf70cpsaptxwa8fw[0:1024-1];
    wire [lhc8m69xvstkozu5iz8i4-1:0]        ewuevraupdwly6mk[0:1024-1];
    wire                                b_mg90m6kvte2my[0:1024-1];
    wire [t5twosugmt3qlv+1:0]           cnuw69qo3fzpi_gvoks[0:512-1];
    wire [lhc8m69xvstkozu5iz8i4-1:0]        x4nde8np28iox7ld6[0:512-1];
    wire                                t7uaatnytij2rxbx_[0:512-1];
    wire [t5twosugmt3qlv+1:0]           wd4tl3kzyo2makk8hmub8ur[0:256-1];
    wire [lhc8m69xvstkozu5iz8i4-1:0]        nllx21_afqb0n56[0:256-1];
    wire                                l0nweuwdfw2kjx[0:256-1];
    wire [t5twosugmt3qlv+1:0]           jtcj0dxaxhjlurc5gfl[0:128-1];
    wire [lhc8m69xvstkozu5iz8i4-1:0]        nzjykoo5f5inx[0:128-1];
    wire                                kn80b7morgbmwi[0:128-1];
    wire  [t5twosugmt3qlv+1:0]          r0ki6qe51tzyh2whxc766ogx6c[0:128-1];
    wire [lhc8m69xvstkozu5iz8i4-1:0]        t7l574slosih7kbpu[0:128-1];
    wire                                dg6zafx148yz8sw3ov[0:128-1];
    wire [t5twosugmt3qlv+1:0]           trj7s2bz3q4vf16py7m[0:64-1];
    wire [lhc8m69xvstkozu5iz8i4-1:0]        f3qfh_jevfed_upqy[0:64-1];
    wire                                q0v1rll39lnx73p7js[0:64-1];
    wire [t5twosugmt3qlv+1:0]           z0hjl1wjq8ei6ieztp1[0:32-1];
    wire [lhc8m69xvstkozu5iz8i4-1:0]        bpp6p7vkmuxq1c[0:32-1];
    wire                                jws7hk88tt3f6b_[0:32-1];
    wire [t5twosugmt3qlv+1:0]           dyox403g0x8m3vk4lq87[0:16-1];
    wire [lhc8m69xvstkozu5iz8i4-1:0]        ojjpx95auel9lv41[0:16-1];
    wire                                vvd1xnft8xsx8fw[0:16-1];
    wire [t5twosugmt3qlv+1:0]           bz51c1m6i9n84p57z04m0cy3[0:8-1];
    wire [lhc8m69xvstkozu5iz8i4-1:0]        z_pjmahhwfs8e3[0:8-1];
    wire                                lhdbc5jp0xhoqkdj_[0:8-1];
    wire [t5twosugmt3qlv+1:0]           vur8dsqh1pl4d0iudz1[0:4-1];
    wire [lhc8m69xvstkozu5iz8i4-1:0]        ru9cuys4dsjqxj[0:4-1];
    wire                                zwxt7psyirz17nv1e[0:4-1];
    wire [t5twosugmt3qlv+1:0]           ji8ld5zj652vb27pp41lxhz[0:2-1];
    wire                                c9knky648tss4r;
    wire                                a1e5qxqwk2vqmi;
    wire [lhc8m69xvstkozu5iz8i4-1:0]        l6hajgyuwup3[0:2-1];
    wire                                rv7mscu1x_nst6unwe[0:2-1];
    wire [t5twosugmt3qlv-1:0]           k6ix738ho6z5n9pf0q; 
    wire [lhc8m69xvstkozu5iz8i4-1:0]        u9168cqr58mcf9o;
    wire                                a3d9_sxxv10x0p2;
    wire                                n1370wxcl1g3pcsc;
    wire [t5twosugmt3qlv-1:0]           unkiitefecxvlolongpdq; 
    wire [lhc8m69xvstkozu5iz8i4-1:0]        mq5j0llnmwskb;
    wire                                v156ejbtigxm;
    wire                                w4u7t2qr86wlre1q_;
    wire [511:0]                        cr3t0k86r4d8agx2ywuo4l;
    wire [255:0]                        fw36sqgo5cj10nugct0k9t9;
    wire [127:0]                        kwwl1u77947opcopu3xorlnuu0y;
    wire [63:0]                         jko9nd77j6nd59psqzrsoyyq23u;
    wire [31:0]                         lkroaab1847a6v6zxyn76uocu1i;
    wire [15:0]                         mge86onnzy09u1ih2r7t8430km;
    wire [7:0]                          rzbzrc0zp54_wj9vzzuoc_0no;
    wire [3:0]                          q6s2jwog3wprf35nkflne621qc;
    wire [1:0]                          la26c47o9w9ovgihtnrdv_s0y;
    wire                                meoguzh3c2qpc_l2pvh5a;
    wire [vb1dh27fsxbyysw-1:0]             fln04o4c2bbbxzho;
    wire                                jjt5ro1ekg7v7uhoesn8f;
    wire [lhc8m69xvstkozu5iz8i4-1:0]        kg87hyc2ic61h2q6wd7j5sb;
    genvar i;
    integer nzd5e;

    wire utcba393zjysral1 = fbzs0o4ysyuzeg_qdj | qaidts35dk5jcji0n;
    
    
    
    
    
    
    assign e6e9h0kbbxy00yvvbp0bywk  = (zvk11dhgg2s67mkq[15:2] == 14'h0);
    assign dc0ovps7up6g7sxmwjd4 = (zvk11dhgg2s67mkq[15:2] == 14'h1);
    assign sgyw532glkiyqyuycg_ymn  = (zvk11dhgg2s67mkq[15:2] == 14'h2);
    
    assign hzql4_1_2nrk6cp7kzhr9mz0  = (zvk11dhgg2s67mkq[15:2] == 14'h802);  

    wire[vb1dh27fsxbyysw-1:0] dbcjt09pmjkdprn;
    assign dbcjt09pmjkdprn[2:0] = 3'b0;
    assign dbcjt09pmjkdprn[3] = a3v1iy5k0; 
    assign dbcjt09pmjkdprn[6:4] = 3'b0;
    assign dbcjt09pmjkdprn[7] = cjwv;
    assign dbcjt09pmjkdprn[10:8] = 3'b0;
    assign dbcjt09pmjkdprn[15:12] = 4'b0;
    assign dbcjt09pmjkdprn[17] = 1'b0;
    assign dbcjt09pmjkdprn[11] = 1'b0;
    assign dbcjt09pmjkdprn[16] = 1'b0;
    assign dbcjt09pmjkdprn[18] = 1'b0;

    generate
    for(i=19; i<vb1dh27fsxbyysw; i=i+1) begin:ftap9xdiknn9iuoyruluvpv3l2pdcq61
                assign dbcjt09pmjkdprn[i] = fcjh1nct4r[i-19];
    end
    endgenerate


    generate
    
    for(i=0; i<vb1dh27fsxbyysw; i=i+1) begin: eul321mfnywpyqngjmh 
        
        assign f63dz5dw05rfd8s39jwx1s_5[i]   = ({18'h0,zvk11dhgg2s67mkq[15:2]} == (($unsigned(i)*4 + 32'h1000)>>2));
        
        
        
        assign enu9bknh9ueizhtexpv7ggo9qoggsu[i] = ({18'h0,zvk11dhgg2s67mkq[15:2]} == (($unsigned(i)*4 + 32'h3000)>>2)) & (utcba393zjysral1 | ((~l6hr3z_7lt62kdb3uv[i])));
        assign e8cte26q6yj870i027qa9r62[i]    =  (f63dz5dw05rfd8s39jwx1s_5[i] | enu9bknh9ueizhtexpv7ggo9qoggsu[i]) & lhibcc3xwm6cy[0];
        assign w0nv2a98k9wdk7ddkoo6wuf5[i]    =  (f63dz5dw05rfd8s39jwx1s_5[i] | enu9bknh9ueizhtexpv7ggo9qoggsu[i]) & lhibcc3xwm6cy[1];
        assign bloeijx3qz0wz5u_avwjaa2we[i]  =  (f63dz5dw05rfd8s39jwx1s_5[i] | enu9bknh9ueizhtexpv7ggo9qoggsu[i]) & lhibcc3xwm6cy[2];
        assign u0xuahg9aulem6ytjre5dm[i]  =  (f63dz5dw05rfd8s39jwx1s_5[i] | enu9bknh9ueizhtexpv7ggo9qoggsu[i]) & lhibcc3xwm6cy[3];
    end
    
    endgenerate


    assign mzp5pkv6xl9_nmhw = fz_isl8q3blzlbl2zzf & e6e9h0kbbxy00yvvbp0bywk & lhibcc3xwm6cy[0];
    assign a7wgjswsdhh5p = {3'b0,u4r4b_6kp09q767q[4:1],1'b1}; 
    ux607_gnrl_dfflr #(7) s0yzi5h3iyop_l(mzp5pkv6xl9_nmhw,a7wgjswsdhh5p[7:1],ufx6dsiuus18[7:1],gf33atgy,ru_wi);
    assign ufx6dsiuus18[0] = 1'b1;

    assign c5a84c6g_dbse_yvi61emns = fz_isl8q3blzlbl2zzf & sgyw532glkiyqyuycg_ymn & lhibcc3xwm6cy[3];
    assign bqe4lf3omz8wflk3ncm1d =  u4r4b_6kp09q767q[31:24];
    ux607_gnrl_dfflr #(8) mv10p4p7dx9_keahj8ax7mmot(c5a84c6g_dbse_yvi61emns,bqe4lf3omz8wflk3ncm1d,bpkwqkepwyytmwn1,gf33atgy,ru_wi);  
    wire [7:0] wcwi_da3mgcgstv7e6b0 = bpkwqkepwyytmwn1;
               
    assign ij34sjy812rgbeddhqm0ts = fz_isl8q3blzlbl2zzf & (sgyw532glkiyqyuycg_ymn | hzql4_1_2nrk6cp7kzhr9mz0) & lhibcc3xwm6cy[1];
    assign ij93945qy0t4clwq0b =  u4r4b_6kp09q767q[15:8];
    ux607_gnrl_dfflr #(8) vohk2f_4rv1gjjyh5x09gt(ij34sjy812rgbeddhqm0ts,ij93945qy0t4clwq0b,uauce93oo4hzcipngfgg,gf33atgy,ru_wi);  
    wire s36z1abpqp = ~(aw82i964do | y8_gkxsfle);
    wire [7:0] qcihcwu9x3x_2vn2dezwl = uauce93oo4hzcipngfgg;
        
    generate
    
    for(i=0; i<vb1dh27fsxbyysw; i=i+1) begin:psex47sw5j7s0cfohh_7dw_o
    if((i < 19) & (i!=3) & (i!=7) 
    ) begin:d8v9pr2euv8ktix_wnxz_ovdi
        assign oyzrjkmgclshj[i] = 8'b0;
        assign k4xratl2pp6xdh98[i] = 1'b0;
    end
    else if(i<19) begin:f3dhh90e8oj77qbaw60rv98mq
        fp3ou97fzh9for8cue9y6 #(
            .iu_89(i),
            .m_rz39tx6bnugdx(lhc8m69xvstkozu5iz8i4)
        ) uc0h3cfrcrfvr5nq4gintqtxrtbkf6sdug(
            .gf33atgy                 (gf33atgy),
            .ru_wi               (ru_wi),
            .dbcjt09pmjkdprn          (dbcjt09pmjkdprn[i]),
            .gsy4z_7std_ruja54_37j  (q_8115sz8oh72wnv9[i][2:1]),
            .jjt5ro1ekg7v7uhoesn8f (jjt5ro1ekg7v7uhoesn8f),  
            .kg87hyc2ic61h2q6wd7j5sb (kg87hyc2ic61h2q6wd7j5sb),
            .e8cte26q6yj870i027qa9r62 (e8cte26q6yj870i027qa9r62[i]),
            .fz_isl8q3blzlbl2zzf    (fz_isl8q3blzlbl2zzf),
            .u4r4b_6kp09q767q       (u4r4b_6kp09q767q),
            .k4xratl2pp6xdh98     (k4xratl2pp6xdh98[i]),
            .oyzrjkmgclshj         (oyzrjkmgclshj[i])
        );
    end
    else begin:l1rp2twfmqca15qgknq3fx77dl
        fp3ou97fzh9for8cue9y6 #(
            .iu_89(i),
            .m_rz39tx6bnugdx(lhc8m69xvstkozu5iz8i4)
        ) vk964470w2_wymc03a42ttvi3coi4ztf8c(
            .gf33atgy                 (gf33atgy),
            .ru_wi               (ru_wi),
            .dbcjt09pmjkdprn          (dbcjt09pmjkdprn[i]),
            .gsy4z_7std_ruja54_37j  (q_8115sz8oh72wnv9[i][2:1]),
            .jjt5ro1ekg7v7uhoesn8f (jjt5ro1ekg7v7uhoesn8f),  
            .kg87hyc2ic61h2q6wd7j5sb (kg87hyc2ic61h2q6wd7j5sb),
            .e8cte26q6yj870i027qa9r62 (e8cte26q6yj870i027qa9r62[i]),
            .fz_isl8q3blzlbl2zzf    (fz_isl8q3blzlbl2zzf),
            .u4r4b_6kp09q767q       (u4r4b_6kp09q767q),
            .k4xratl2pp6xdh98     (k4xratl2pp6xdh98[i]),
            .oyzrjkmgclshj         (oyzrjkmgclshj[i])
        );

    end

    if((i < 19) & (i!=3) & (i!=7)
                ) begin:r2ufmfs32hlmsx33ckhm1n
            assign mglzjmd3n4ynn8[i] = {{(t5twosugmt3qlv){1'b0}},{(8-t5twosugmt3qlv){1'b1}}}; 
            assign mysay5szii2i_ucs[i] = {2'b11,6'b0};
            assign wvmr61jza7zhd5o0u[i] = 8'b0;
            assign tbf0wzltxdlu9ouilvocb_f62[i] = 1'b0;
    end
    else begin:i6hr1xzre4rv8fnpv7lx5ko5to8
        assign wvmr61jza7zhd5o0u[i] = {7'b0,u4r4b_6kp09q767q[8]};
        if(i>=19) begin:n7m6mw92b9joxwz59a0ycc2x
        
        assign tbf0wzltxdlu9ouilvocb_f62[i] = (utcba393zjysral1 | f63dz5dw05rfd8s39jwx1s_5[i]) ? ((u4r4b_6kp09q767q[23:22] == 2'b11) ? 1'b1 : (u4r4b_6kp09q767q[23:22] == 2'b01) ? 1'b0 : q_8115sz8oh72wnv9[i][7]) : q_8115sz8oh72wnv9[i][7];
        assign mysay5szii2i_ucs[i] = {tbf0wzltxdlu9ouilvocb_f62[i],1'b1,3'b0,u4r4b_6kp09q767q[18:16]};
        end
        else begin:bynlgnmz94ftqthutguz9f2kq6fv
        assign tbf0wzltxdlu9ouilvocb_f62[i] = (utcba393zjysral1 | f63dz5dw05rfd8s39jwx1s_5[i]) ? ((u4r4b_6kp09q767q[23:22] == 2'b11) ? 1'b1 : (u4r4b_6kp09q767q[23:22] == 2'b01) ? 1'b0 : q_8115sz8oh72wnv9[i][7]) : q_8115sz8oh72wnv9[i][7];
        assign mysay5szii2i_ucs[i] = {tbf0wzltxdlu9ouilvocb_f62[i],1'b1,3'b0,u4r4b_6kp09q767q[18:16]};
        end
        assign mglzjmd3n4ynn8[i] = {u4r4b_6kp09q767q[31 -: t5twosugmt3qlv], {(8-t5twosugmt3qlv){1'b1}}}; 
    end

        assign q9dddg5qvq6azwmv5[i] = fz_isl8q3blzlbl2zzf & u0xuahg9aulem6ytjre5dm[i];
        assign sc9i3oongjhvjssm8b[i] = fz_isl8q3blzlbl2zzf & bloeijx3qz0wz5u_avwjaa2we[i];
        assign dcs94jjnvo_oqe_[i] = fz_isl8q3blzlbl2zzf & w0nv2a98k9wdk7ddkoo6wuf5[i];
    
        if(t5twosugmt3qlv>=8) begin:h4c20j978b1t5vycxvqf16skwomw9ryubjb5c72hn2
        ux607_gnrl_dfflr #(8) dxdl2mmbom2x6i6kzx(q9dddg5qvq6azwmv5[i],mglzjmd3n4ynn8[i][7:0],z1gysizgxf7x[i][7:0],gf33atgy,ru_wi);  
        end
        else begin:giotpjx1vb_1hbuudzo7v1n3k4ih5tkopot1qbud
        ux607_gnrl_dfflr #(t5twosugmt3qlv) v24hzm8luqmn0vveq0ta443g(q9dddg5qvq6azwmv5[i],mglzjmd3n4ynn8[i][7-:t5twosugmt3qlv],z1gysizgxf7x[i][7-:t5twosugmt3qlv],gf33atgy,ru_wi);  
        assign z1gysizgxf7x[i][7-t5twosugmt3qlv:0] = {(8-t5twosugmt3qlv){1'b1}};
        end
        ux607_gnrl_dfflr #(6) haovvbdr3i1ew6ko5t5kr5f4a(sc9i3oongjhvjssm8b[i],mysay5szii2i_ucs[i][5:0],q_8115sz8oh72wnv9[i][5:0],gf33atgy,ru_wi);  
        ux607_gnrl_dfflrs #(1) b0frn_t_uulfyrj9mybkfjt(sc9i3oongjhvjssm8b[i],mysay5szii2i_ucs[i][7],q_8115sz8oh72wnv9[i][7],gf33atgy,ru_wi);  
        assign q_8115sz8oh72wnv9[i][6] = 1'b1;
        assign l6hr3z_7lt62kdb3uv[i] = q_8115sz8oh72wnv9[i][7];
        ux607_gnrl_dfflr #(8) j4m8oc7fqqts0o3bbk(dcs94jjnvo_oqe_[i],wvmr61jza7zhd5o0u[i],qhzxh33vz7eo6[i],gf33atgy,ru_wi);  
    end
    
    endgenerate





   assign lva2sw2f_nq_1u5780  = {32{e6e9h0kbbxy00yvvbp0bywk}} & {24'b0, 1'b0, 2'b1, oi2196y9j6yk8xp9,1'b1};  
   wire [3:0] sogvxn7eczpk420 = t5twosugmt3qlv[3:0];
   wire [7:0] a0m0antr5oslt = ujp_32rzn[7:0];
   wire [12:0] hr5o7d7xwjcshvl = vb1dh27fsxbyysw[12:0];
   assign l05bm7_xtgbitxwsk_3 = {32{dc0ovps7up6g7sxmwjd4}} & {7'b0,sogvxn7eczpk420,a0m0antr5oslt,hr5o7d7xwjcshvl};
   
   assign w5t0kiz2tj15hher468m_ngc = {32{sgyw532glkiyqyuycg_ymn}} & {bpkwqkepwyytmwn1,8'b0,uauce93oo4hzcipngfgg,8'h0};
   assign hkmb5i4b7onky8b45mmb4l6y = {32{hzql4_1_2nrk6cp7kzhr9mz0}} & {16'b0,uauce93oo4hzcipngfgg,8'h0};
   always @* begin:u8idprjl7175qq_jbsbyq
       isd23fnq13pcssxpxiacb  = 32'b0;
       for(nzd5e=0; nzd5e<vb1dh27fsxbyysw; nzd5e=nzd5e+1) begin: j49wg_eq195lu
            isd23fnq13pcssxpxiacb  =  isd23fnq13pcssxpxiacb  | ({32{(f63dz5dw05rfd8s39jwx1s_5[nzd5e] | enu9bknh9ueizhtexpv7ggo9qoggsu[nzd5e])}} &
                                                  {z1gysizgxf7x[nzd5e],
                                                   
                                                   q_8115sz8oh72wnv9[nzd5e],
                                                   
                                                   
                                                   
                                                   
                                                   
                                                   qhzxh33vz7eo6[nzd5e],
                                                   oyzrjkmgclshj[nzd5e]}
                                                 );
       end
   end







    wire [32-1:0] vf_r9hn9ty7axn         = lva2sw2f_nq_1u5780 
                                    | l05bm7_xtgbitxwsk_3 
                                    | w5t0kiz2tj15hher468m_ngc 
                                    | hkmb5i4b7onky8b45mmb4l6y 
                                    | isd23fnq13pcssxpxiacb;
    





   generate


    for(i=0; i<vb1dh27fsxbyysw; i=i+1) begin:gwtmuqg71vqzj20
        assign x3g5a2s4f40otq82g[i] = q_8115sz8oh72wnv9[i][0];
        assign fln04o4c2bbbxzho[i] = qhzxh33vz7eo6[i][0] & oyzrjkmgclshj[i][0];
        assign cs8o9yf70cpsaptxwa8fw[i] =  {fln04o4c2bbbxzho[i],l6hr3z_7lt62kdb3uv[i],z1gysizgxf7x[i][7 -: t5twosugmt3qlv]}; 
        assign ewuevraupdwly6mk[i] = i[lhc8m69xvstkozu5iz8i4-1:0];
        assign b_mg90m6kvte2my[i] = x3g5a2s4f40otq82g[i];
    end

    
    for(i=vb1dh27fsxbyysw; i<1024; i=i+1) begin:o1o7cansg6fjuqpt2k1qov97bg
        assign cs8o9yf70cpsaptxwa8fw[i] = {(t5twosugmt3qlv+1){1'b0}};
        assign ewuevraupdwly6mk[i] = {lhc8m69xvstkozu5iz8i4{1'b0}};
        assign b_mg90m6kvte2my[i] = 1'b0;
    end


    
    for(i=0; i<512; i=i+1) begin: urf7puwurdc7nugl5b
        assign cr3t0k86r4d8agx2ywuo4l[i] = (cs8o9yf70cpsaptxwa8fw[(2*i) + 1] < cs8o9yf70cpsaptxwa8fw[2*i]);
        assign cnuw69qo3fzpi_gvoks[i] =  cr3t0k86r4d8agx2ywuo4l[i] ? cs8o9yf70cpsaptxwa8fw[2*i]:cs8o9yf70cpsaptxwa8fw[(2*i) + 1];
        assign x4nde8np28iox7ld6[i] =   cr3t0k86r4d8agx2ywuo4l[i] ? ewuevraupdwly6mk[2*i] : ewuevraupdwly6mk[(2*i) + 1];
        assign t7uaatnytij2rxbx_[i] =   cr3t0k86r4d8agx2ywuo4l[i] ? b_mg90m6kvte2my[2*i] : b_mg90m6kvte2my[(2*i) + 1];
    end

    
    for(i=0; i<256; i=i+1) begin: wc3v_g425z367q1mue1
        assign fw36sqgo5cj10nugct0k9t9[i] = (cnuw69qo3fzpi_gvoks[(2*i) + 1] < cnuw69qo3fzpi_gvoks[2*i]);
        assign wd4tl3kzyo2makk8hmub8ur[i] =  fw36sqgo5cj10nugct0k9t9[i] ? cnuw69qo3fzpi_gvoks[2*i]:cnuw69qo3fzpi_gvoks[(2*i) + 1];
        assign nllx21_afqb0n56[i] =   fw36sqgo5cj10nugct0k9t9[i] ? x4nde8np28iox7ld6[2*i] : x4nde8np28iox7ld6[(2*i) + 1];
        assign l0nweuwdfw2kjx[i] =   fw36sqgo5cj10nugct0k9t9[i] ? t7uaatnytij2rxbx_[2*i] : t7uaatnytij2rxbx_[(2*i) + 1];
    end

    
    for(i=0; i<128; i=i+1) begin: mqjkd_lrrz3fh3cwm7668y
        assign kwwl1u77947opcopu3xorlnuu0y[i] = (wd4tl3kzyo2makk8hmub8ur[(2*i) + 1] < wd4tl3kzyo2makk8hmub8ur[2*i]);
        assign jtcj0dxaxhjlurc5gfl[i] =  kwwl1u77947opcopu3xorlnuu0y[i] ? wd4tl3kzyo2makk8hmub8ur[2*i]:wd4tl3kzyo2makk8hmub8ur[(2*i) + 1];
        assign nzjykoo5f5inx[i] =   kwwl1u77947opcopu3xorlnuu0y[i] ? nllx21_afqb0n56[2*i] : nllx21_afqb0n56[(2*i) + 1];
        assign kn80b7morgbmwi[i] =   kwwl1u77947opcopu3xorlnuu0y[i] ? l0nweuwdfw2kjx[2*i] : l0nweuwdfw2kjx[(2*i) + 1];
    end

    for(i=0; i<128; i=i+1) begin: i5g9bwdixwjzeu5gwpeui5vw873sl
        ux607_gnrl_dffr #(t5twosugmt3qlv+2) osm8xku3wk9tvo0bka574hsae7nm(jtcj0dxaxhjlurc5gfl[i], r0ki6qe51tzyh2whxc766ogx6c[i], gf33atgy, ru_wi);
        ux607_gnrl_dffr #(lhc8m69xvstkozu5iz8i4) pxtzz1ympqvv4rq8o(nzjykoo5f5inx[i], t7l574slosih7kbpu[i], gf33atgy, ru_wi); 
        ux607_gnrl_dffr #(1) dkv10jhkal27hpo5caq5wu(kn80b7morgbmwi[i], dg6zafx148yz8sw3ov[i], gf33atgy, ru_wi);
    end

    
    for(i=0; i<64; i=i+1) begin: skn1r4f7vtna16hnlfx
        assign jko9nd77j6nd59psqzrsoyyq23u[i] = (r0ki6qe51tzyh2whxc766ogx6c[(2*i) + 1] < r0ki6qe51tzyh2whxc766ogx6c[2*i]);
        assign trj7s2bz3q4vf16py7m[i] =  jko9nd77j6nd59psqzrsoyyq23u[i] ? r0ki6qe51tzyh2whxc766ogx6c[2*i]:r0ki6qe51tzyh2whxc766ogx6c[(2*i) + 1];
        assign f3qfh_jevfed_upqy[i] =   jko9nd77j6nd59psqzrsoyyq23u[i] ? t7l574slosih7kbpu[2*i] : t7l574slosih7kbpu[(2*i) + 1];
        assign q0v1rll39lnx73p7js[i] =   jko9nd77j6nd59psqzrsoyyq23u[i] ? dg6zafx148yz8sw3ov[2*i] : dg6zafx148yz8sw3ov[(2*i) + 1];
    end


    
    for(i=0; i<32; i=i+1) begin: xcws65db8uymiaoyop6
        assign lkroaab1847a6v6zxyn76uocu1i[i] = (trj7s2bz3q4vf16py7m[(2*i) + 1] < trj7s2bz3q4vf16py7m[2*i]);
        assign z0hjl1wjq8ei6ieztp1[i] =  lkroaab1847a6v6zxyn76uocu1i[i] ? trj7s2bz3q4vf16py7m[2*i]:trj7s2bz3q4vf16py7m[(2*i) + 1];
        assign bpp6p7vkmuxq1c[i] =   lkroaab1847a6v6zxyn76uocu1i[i] ? f3qfh_jevfed_upqy[2*i] : f3qfh_jevfed_upqy[(2*i) + 1];
        assign jws7hk88tt3f6b_[i] =   lkroaab1847a6v6zxyn76uocu1i[i] ? q0v1rll39lnx73p7js[2*i] : q0v1rll39lnx73p7js[(2*i) + 1];
    end

    
    for(i=0; i<16; i=i+1) begin: tg8js04ob2c6l_h3uoe9
        assign mge86onnzy09u1ih2r7t8430km[i] = (z0hjl1wjq8ei6ieztp1[(2*i) + 1] < z0hjl1wjq8ei6ieztp1[2*i]);
        assign dyox403g0x8m3vk4lq87[i] =  mge86onnzy09u1ih2r7t8430km[i] ? z0hjl1wjq8ei6ieztp1[2*i]:z0hjl1wjq8ei6ieztp1[(2*i) + 1];
        assign ojjpx95auel9lv41[i] =   mge86onnzy09u1ih2r7t8430km[i] ? bpp6p7vkmuxq1c[2*i] : bpp6p7vkmuxq1c[(2*i) + 1];
        assign vvd1xnft8xsx8fw[i] =   mge86onnzy09u1ih2r7t8430km[i] ? jws7hk88tt3f6b_[2*i] : jws7hk88tt3f6b_[(2*i) + 1];
    end

    
    for(i=0; i<8; i=i+1) begin: re0wlw7suywy3dyogou
        assign rzbzrc0zp54_wj9vzzuoc_0no[i] = (dyox403g0x8m3vk4lq87[(2*i) + 1] < dyox403g0x8m3vk4lq87[2*i]);
        assign bz51c1m6i9n84p57z04m0cy3[i] =  rzbzrc0zp54_wj9vzzuoc_0no[i] ? dyox403g0x8m3vk4lq87[2*i]:dyox403g0x8m3vk4lq87[(2*i) + 1];
        assign z_pjmahhwfs8e3[i] =   rzbzrc0zp54_wj9vzzuoc_0no[i] ? ojjpx95auel9lv41[2*i] : ojjpx95auel9lv41[(2*i) + 1];
        assign lhdbc5jp0xhoqkdj_[i] =   rzbzrc0zp54_wj9vzzuoc_0no[i] ? vvd1xnft8xsx8fw[2*i] : vvd1xnft8xsx8fw[(2*i) + 1];
    end

    
    for(i=0; i<4; i=i+1) begin: psptlzby4f1z2uux_h
        assign q6s2jwog3wprf35nkflne621qc[i] = (bz51c1m6i9n84p57z04m0cy3[(2*i) + 1] < bz51c1m6i9n84p57z04m0cy3[2*i]);
        assign vur8dsqh1pl4d0iudz1[i] =  q6s2jwog3wprf35nkflne621qc[i] ? bz51c1m6i9n84p57z04m0cy3[2*i]:bz51c1m6i9n84p57z04m0cy3[(2*i) + 1];
        assign ru9cuys4dsjqxj[i] =   q6s2jwog3wprf35nkflne621qc[i] ? z_pjmahhwfs8e3[2*i] : z_pjmahhwfs8e3[(2*i) + 1];
        assign zwxt7psyirz17nv1e[i] =   q6s2jwog3wprf35nkflne621qc[i] ? lhdbc5jp0xhoqkdj_[2*i] : lhdbc5jp0xhoqkdj_[(2*i) + 1];
    end

    
    for(i=0; i<2; i=i+1) begin: ui067tw1gk66engyjixnwg
        assign la26c47o9w9ovgihtnrdv_s0y[i] = (vur8dsqh1pl4d0iudz1[(2*i) + 1] < vur8dsqh1pl4d0iudz1[2*i]);
        assign ji8ld5zj652vb27pp41lxhz[i] =  la26c47o9w9ovgihtnrdv_s0y[i] ? vur8dsqh1pl4d0iudz1[2*i]:vur8dsqh1pl4d0iudz1[(2*i) + 1];
        assign l6hajgyuwup3[i] =   la26c47o9w9ovgihtnrdv_s0y[i] ? ru9cuys4dsjqxj[2*i] : ru9cuys4dsjqxj[(2*i) + 1];
        assign rv7mscu1x_nst6unwe[i] =   la26c47o9w9ovgihtnrdv_s0y[i] ? zwxt7psyirz17nv1e[2*i] : zwxt7psyirz17nv1e[(2*i) + 1];
    end

    endgenerate

    assign meoguzh3c2qpc_l2pvh5a = (ji8ld5zj652vb27pp41lxhz[1] < ji8ld5zj652vb27pp41lxhz[0]);
    assign a3d9_sxxv10x0p2           = meoguzh3c2qpc_l2pvh5a ? ji8ld5zj652vb27pp41lxhz[0][t5twosugmt3qlv+1] :
                                                         ji8ld5zj652vb27pp41lxhz[1][t5twosugmt3qlv+1];
    assign c9knky648tss4r         = meoguzh3c2qpc_l2pvh5a ? ji8ld5zj652vb27pp41lxhz[0][t5twosugmt3qlv] :
                                                         ji8ld5zj652vb27pp41lxhz[1][t5twosugmt3qlv];
    assign k6ix738ho6z5n9pf0q    = {t5twosugmt3qlv{a3d9_sxxv10x0p2}} & (meoguzh3c2qpc_l2pvh5a ? ji8ld5zj652vb27pp41lxhz[0][t5twosugmt3qlv-1:0] : 
                                                                                         ji8ld5zj652vb27pp41lxhz[1][t5twosugmt3qlv-1:0]);
    assign u9168cqr58mcf9o           = {lhc8m69xvstkozu5iz8i4{a3d9_sxxv10x0p2}} & (meoguzh3c2qpc_l2pvh5a ? l6hajgyuwup3[0] :
                                                                       l6hajgyuwup3[1]);
    assign n1370wxcl1g3pcsc          = a3d9_sxxv10x0p2 & (meoguzh3c2qpc_l2pvh5a ? rv7mscu1x_nst6unwe[0] : 
                                                                       rv7mscu1x_nst6unwe[1]);

        ux607_gnrl_dffr #(t5twosugmt3qlv) ejs1o5j1fvikvrf5t4fl(k6ix738ho6z5n9pf0q,unkiitefecxvlolongpdq,gf33atgy,ru_wi);  
        ux607_gnrl_dffr #(lhc8m69xvstkozu5iz8i4) gds432n4omzp(u9168cqr58mcf9o,mq5j0llnmwskb,gf33atgy,ru_wi);  
        ux607_gnrl_dffr #(1) ta1qj9ime4d3x(a3d9_sxxv10x0p2,v156ejbtigxm,gf33atgy,ru_wi);  
        ux607_gnrl_dffr #(1) iq56zi5d6a1t(n1370wxcl1g3pcsc,w4u7t2qr86wlre1q_,gf33atgy,ru_wi);  
        ux607_gnrl_dffr #(1) p4cg94smv6vj2(c9knky648tss4r,a1e5qxqwk2vqmi,gf33atgy,ru_wi);  

    wire [7:0] wrlrjvi6kd5yb;
    wire t3xdb_t72bki0btjk_   = gfy3zost37aq8qmr ? (a1e5qxqwk2vqmi ? (wrlrjvi6kd5yb > f_i1959b4xizzq9jea) : 1'b0) : 1'b1;
    wire pa6pp7c5fx_xe1wd   = gfy3zost37aq8qmr ? (a1e5qxqwk2vqmi ? 1'b0 : (wrlrjvi6kd5yb > tcy_87vt9vet39knuw)) : 1'b1;
    wire [7:0] i25ob9bayn6qsp84sh = {unkiitefecxvlolongpdq,{{(8-t5twosugmt3qlv)}{1'b1}}}; 
    wire [7:0] wtk0ob6j34cx4h76dih = 8'hff >> oi2196y9j6yk8xp9;
    assign wrlrjvi6kd5yb = {8{v156ejbtigxm}} & (wtk0ob6j34cx4h76dih | i25ob9bayn6qsp84sh); 
    assign znzjygllppv1s0a8cqub3c  = v156ejbtigxm & a1e5qxqwk2vqmi  & (wrlrjvi6kd5yb[7:0] > wcwi_da3mgcgstv7e6b0[7:0]);
    assign fc_4ns_w1nh4h02z_dgg = v156ejbtigxm & ~a1e5qxqwk2vqmi & (wrlrjvi6kd5yb[7:0] > qcihcwu9x3x_2vn2dezwl[7:0]);
    wire mfquy8ep091a9agpv48_ombh1 =  ((dz0zrf512290tvcy4q & zwcbp7zqfei5xz) | dxi_ue3gf5zqqqxwgq2a | fzdb65fcrotwcaccus_cwo);
    ux607_gnrl_dffr #(1) ec9t3w75eqvb0tz9_qkg8gbmpm3569x(mfquy8ep091a9agpv48_ombh1, jjt5ro1ekg7v7uhoesn8f, zh6e0v0mmz, ru_wi);
    ux607_gnrl_dfflr #(lhc8m69xvstkozu5iz8i4) vqt5gm74bli39h5r2ssriytwy_9hyhs3(mfquy8ep091a9agpv48_ombh1, mq5j0llnmwskb, kg87hyc2ic61h2q6wd7j5sb, zh6e0v0mmz, ru_wi);



        ux607_gnrl_pipe_stage # (
          .CUT_READY(0),
          .DP(1),
          .DW(32)
        ) cqc6bg2e20t9lh9m3z0ggh (
          .i_vld  (th06du2c8e2_b7k),
          .i_rdy  (irjoi8wvo25u209f_5),
          .i_dat  (vf_r9hn9ty7axn),
          .o_vld  (klkflmsyyf5w7ar),
          .o_rdy  (wy36iirxspfw56864),  
          .o_dat  (h7f6k_ims_9p3),   
        
          .clk  (gf33atgy),
          .rst_n(ru_wi)
        );

    assign lkjqs6kiuyj   = 1'b0;
    wire oxvzs1izpx1rv_0t2_ = 1'b1;
    assign kfrxhvr3mwznw    = a1e5qxqwk2vqmi ? dn8riluj40uunvq5 & (znzjygllppv1s0a8cqub3c & t3xdb_t72bki0btjk_) & oxvzs1izpx1rv_0t2_ :
                                            
                                            (~aw82i964do) & dn8riluj40uunvq5 & (fc_4ns_w1nh4h02z_dgg & pa6pp7c5fx_xe1wd) & oxvzs1izpx1rv_0t2_;
    assign jqsukc5b5drcc1e78  = a1e5qxqwk2vqmi;
    assign gnn46rd7vvofruqij  = ~a1e5qxqwk2vqmi;
    assign hjrk_rwjkqj3zk_b  = wrlrjvi6kd5yb;
    assign zwcbp7zqfei5xz  = w4u7t2qr86wlre1q_;
    assign b4lwcgm6l21pi   = {{(10-lhc8m69xvstkozu5iz8i4){1'b0}},mq5j0llnmwskb};


wire h_qfp9y_34txjy4hsx4y7 = |k4xratl2pp6xdh98; 
wire faqyp35jo48d5m9stfa2oxm = jjt5ro1ekg7v7uhoesn8f;
wire nt0n66a2e33vnm4fvdl = h_qfp9y_34txjy4hsx4y7 | faqyp35jo48d5m9stfa2oxm; 

wire s9sdzfpg_djffkp7;
wire sw0dt4a0crqnk1nadh;
wire f25z101uq1xxwx;
wire z0ztwxvsjsx7u55_u;

assign s9sdzfpg_djffkp7 = (|fln04o4c2bbbxzho) | th06du2c8e2_b7k | klkflmsyyf5w7ar | nt0n66a2e33vnm4fvdl
                    | v156ejbtigxm 
                    ;

ux607_gnrl_dffr #(1) vvcuigf2mszqzb_n2rtm4ymixddeyz_ddrf(s9sdzfpg_djffkp7, sw0dt4a0crqnk1nadh, dk2xhkj77a, ru_wi); 
ux607_gnrl_dffr #(1) tu1woi_yv2n_eolh5koim0zypfgnmf(sw0dt4a0crqnk1nadh, f25z101uq1xxwx, dk2xhkj77a, ru_wi); 
ux607_gnrl_dffr #(1) q2l83er2cfuco1j_jh330kkrguciump(f25z101uq1xxwx, z0ztwxvsjsx7u55_u, dk2xhkj77a, ru_wi); 


    assign y12wg4mlovhn13   = s9sdzfpg_djffkp7 | sw0dt4a0crqnk1nadh | f25z101uq1xxwx | z0ztwxvsjsx7u55_u; 

endmodule




















module w0v8rrkl3p_ar0i2l (

    
  input rb050tnl,
  input a94vd35etec4,
  input el7_p8jit09,
  input [12-1:0] e1go3iu,
  input izhvh9xxvwe2,
  input  [64-1:0] vf5xcr67bqhzlo43_,
  output [64-1:0] l9erxxpnphqd26vg9,
  output u2dvoyt5e7o_03z9z5,
  output s904ol6a25v9zn8,


    
  input  [64-1:0] qeb3z0x5,
  input  ibhfuwrztbm8p4gg,

  input  [3-1:0] i8_5wt0vppx,
  input  osv2437qj_3nuf,



  input  b7g_vsn0zoewh6g1,
  input  [2-1:0] onnv64ydiajl,
  output [2-1:0] r21i4by0bu3ks,

    
  output [64*4-1:0] azll7rq5fab5ou,
  output [64*4-1:0] n6a0r_0zddzrme8,
  input  ns0i7siujgkrghjpqv6,


  output[64-1:0]  hn85hkp2yav,

  output pydatzxqqi,
  output t5trf35s8vy,
  output zbac123pv78sbz3,
  output z4e_m564fxae0kpbjr,

  output zmwq3e9oijvo7d7,
  output q4gqhurcazjpsf4h,

  output hixy2y36a1pn0,
  output ozwene1gdpatk6g,
  output sxvvsxtbhyvt,
  input  rn1o3sl83,

  input  gf33atgy,
  input  ru_wi
  );

 
localparam m0xuxgjqd7dh8v = (4<=2)?1:(4<=4)?2:(4<=8)?3:(4<=16)?4:(4<=32)?5:(4<=64)?6:(4<=128)?7:(4<=256)?8:(4<=512)?9:(4<=1024)?10:(4<=2048)?11:(4<=4096)?12:-1;

wire [64-1:0] dwns7g;
wire [64-1:0] dpc_r;
wire [64-1:0] hm52hlju8jce9ftg;





wire wgglybxiqwjpz3e      = (e1go3iu == 12'h7b0);
wire fouak3vibvtau       = (e1go3iu == 12'h7b1);
wire q0pyqbf15tu4tdzww9 = (e1go3iu == 12'h7b2);



wire [64-1:0] sj2yfdnj4ur_c;
wire efi9tetop_99b9m6qjm2 = (e1go3iu == 12'h7b3);
wire b6itbh9qe_5t_kym71 = pydatzxqqi & efi9tetop_99b9m6qjm2;
wire b5nnug9khey4 = el7_p8jit09 & b6itbh9qe_5t_kym71;

wire c6lbvkska6qd      = pydatzxqqi & wgglybxiqwjpz3e     ;
wire t6furl_ir_       = pydatzxqqi & fouak3vibvtau      ;
wire tjd7oh5_8uvknv6 = pydatzxqqi & q0pyqbf15tu4tdzww9;


assign s904ol6a25v9zn8 = (~pydatzxqqi) & ( 
              wgglybxiqwjpz3e      
            | fouak3vibvtau       
            | q0pyqbf15tu4tdzww9 
            | efi9tetop_99b9m6qjm2 
            );

wire zigaf2rxnzht     = el7_p8jit09 & c6lbvkska6qd    ;
wire ug2z6sy1f      = el7_p8jit09 & t6furl_ir_     ;
wire t8dvdarletf2muh9e = el7_p8jit09 & tjd7oh5_8uvknv6;

wire gunt8gr89tq2  = (e1go3iu == 12'h7a0);
wire b00s0p78drh4z   = (e1go3iu == 12'h7a1);
wire lxcp51g29nqalv   = (e1go3iu == 12'h7a2);
wire tzfj8xp6rkw   = (e1go3iu == 12'h7a3);
wire cjgwj883m1    = (e1go3iu == 12'h7a4);
wire t13mpjnjkl0_uyhwq = (e1go3iu == 12'h7a8);
wire xnt1ut20a4q_x5 = (e1go3iu == 12'h7a3);

wire ajfyzjug7yq2_  =  el7_p8jit09 & gunt8gr89tq2 ;
wire ouuky5aoj_   =  el7_p8jit09 & b00s0p78drh4z  ;
wire q4yijhm2w_lc   =  el7_p8jit09 & lxcp51g29nqalv  ;
wire z6uhklntahxl50   =  el7_p8jit09 & tzfj8xp6rkw  ;
wire rdm1b6tcy9pok    =  el7_p8jit09 & cjgwj883m1   ;
wire osz1c5t4rbjefe =  el7_p8jit09 & t13mpjnjkl0_uyhwq;
wire wypmavpknwip0dg =  el7_p8jit09 & xnt1ut20a4q_x5;

wire nxb2bijaqvnh2w7m9ga  = izhvh9xxvwe2 & gunt8gr89tq2 ;
wire da36aklh2x1yugbf   = izhvh9xxvwe2 & b00s0p78drh4z  ;
wire idm817wr_az479   = izhvh9xxvwe2 & lxcp51g29nqalv  ;

wire [64-1:0] rbz9x0m18nf7d ;
wire [64-1:0] z585kaqlq5f76 ;
wire [64-1:0] b7iuqg01sm8apr ;
wire [64-1:0] olpetlafep   = rbz9x0m18nf7d ;
wire [64-1:0] np4_f1v03ag   = z585kaqlq5f76 ;
wire [64-1:0] vat77cznsta   = 64'b0 ;
   
   
   
wire [64-1:0] u_ni4ncd78b    = {{64-6{1'b0}},4'b1111,2'b0};
wire [64-1:0] qc39qez5cu8  = b7iuqg01sm8apr ;


wire b_a74a2_dk7xhm     = izhvh9xxvwe2 & c6lbvkska6qd    ;
wire ip016fpv80afgj6      = izhvh9xxvwe2 & t6furl_ir_     ;
wire lxb0f8_9_lvkjx2laso1s = izhvh9xxvwe2 & tjd7oh5_8uvknv6;
wire nmfco0vb59lfudihij7 = izhvh9xxvwe2 & b6itbh9qe_5t_kym71;



wire [64-1:0] tanak2a4v784w     = dwns7g    ;
wire [64-1:0] vgtsmf4if4o      = dpc_r     ;
wire [64-1:0] g4u9fas1jthrb0cjye = hm52hlju8jce9ftg;
wire [64-1:0] pl0eyz4550dld = sj2yfdnj4ur_c;


assign {u2dvoyt5e7o_03z9z5, l9erxxpnphqd26vg9} = {1'b0,64'b0} 
               | {wgglybxiqwjpz3e    ,({64{zigaf2rxnzht       }} & tanak2a4v784w    )      }
               | {fouak3vibvtau     ,({64{ug2z6sy1f        }} & vgtsmf4if4o     )      }
               | {q0pyqbf15tu4tdzww9,({64{t8dvdarletf2muh9e   }} & g4u9fas1jthrb0cjye)      }
               | {efi9tetop_99b9m6qjm2,({64{b5nnug9khey4   }} & pl0eyz4550dld)      }
               | {gunt8gr89tq2, ({64{ajfyzjug7yq2_    }} & qc39qez5cu8)       }
               | {b00s0p78drh4z , ({64{ouuky5aoj_     }} & olpetlafep)        }
               | {lxcp51g29nqalv , ({64{q4yijhm2w_lc     }} & np4_f1v03ag)        }
               | {tzfj8xp6rkw , ({64{z6uhklntahxl50     }} & vat77cznsta)        }
               | {cjgwj883m1  , ({64{rdm1b6tcy9pok      }} & u_ni4ncd78b )        }
               | {t13mpjnjkl0_uyhwq  , ({64{osz1c5t4rbjefe}} & {64{1'b0}} )        }
               | {xnt1ut20a4q_x5  , ({64{wypmavpknwip0dg}} & {64{1'b0}} )        }
               ;


assign hn85hkp2yav = dpc_r;



  wire dpc_ena;
  wire [64-1:0] dpc_nxt;
  assign dpc_ena = ip016fpv80afgj6 | ibhfuwrztbm8p4gg;
  assign dpc_nxt[64-1:1] = 
       ibhfuwrztbm8p4gg ? qeb3z0x5[64-1:1] 
                   : vf5xcr67bqhzlo43_[64-1:1];
  assign dpc_nxt[0] = 1'b0; 
  ux607_gnrl_dfflr #(64) q5wvskd7n (dpc_ena, dpc_nxt, dpc_r, gf33atgy, ru_wi);
  

  wire hgn4cf157ngjvbja2 = lxb0f8_9_lvkjx2laso1s;
  wire [64-1:0] w6rc11qukmyn2r3_tr;
  assign w6rc11qukmyn2r3_tr = vf5xcr67bqhzlo43_;
  ux607_gnrl_dfflr #(64) zfzba2zhnlkc51p2l1 (hgn4cf157ngjvbja2, w6rc11qukmyn2r3_tr, hm52hlju8jce9ftg, gf33atgy, ru_wi);
 
  wire vm7j0eia8z0jov = nmfco0vb59lfudihij7;
  wire [64-1:0] d0wpu344ab5mae;
  assign d0wpu344ab5mae = vf5xcr67bqhzlo43_;
  ux607_gnrl_dfflr #(64) azbvumrn8h6_06o (vm7j0eia8z0jov, d0wpu344ab5mae, sj2yfdnj4ur_c, gf33atgy, ru_wi);
 

  wire[64-1:0] dwt4xr7nj [0:4-1];
  wire[64-1:0] qzr9ikzg_vz [0:4-1];
  wire[4-1:0] bt36dhn0q97o3x;
  wire[4-1:0] dgv2oqmmc685v;
  wire[4-1:0] fv66706su4xcaxv;
  wire[4-1:0] rx3dpavi0xj7b4gx;
  wire[4-1:0] ornx_vnpekug3gz;
  wire[4-1:0] il72jv39takrecodwjg[0:4-1];
  wire[4-1:0] l37vb0thqk484l    [0:4-1];
  wire[4-1:0] ox0hspotahshker242;
  wire[4-1:0] f_en44nuq7wxpi6;
  wire[4-1:0] zdauex3dn6kp7jfh;
  wire[4-1:0] lc7l4i7ez6dwylrrke;
  wire[4-1:0] lublr8yrk2iclyv1090;
  wire[4-1:0] qytl9l30d1xwc77h3;
  wire[4-1:0] ekcdji6jnpih8_4dk2tc;
  wire[4-1:0] s4yy9maabthu6i_jf9svf8;
  wire[4-1:0] n24f03wv5exza5j6or0c;
  wire[1-1:0] egctw8sjve74zbjm64f2[0:4-1];
  wire[1-1:0] p389kv4igf_ei2d    [0:4-1];
  wire[4-1:0] dlgms2ikbd24vp0r2;
  wire[59-1:0] lsh9e8uas4hp15ahg1j[0:4-1];
  wire[59-1:0] hev3ez6yazmxe    [0:4-1];
  wire[59-1:0] cn5uuiza89o2dulas69s    [0:4-1];
  wire[4-1:0] vr0xmfp80ka92vtnhtwvnuyf;
  wire[4-1:0] m_44xky76stmh65migajp7t;
  wire[3:0] mfu6jps217vim6x17jhy[0:4-1];


  wire ybn5wo3zvbsf5 = nxb2bijaqvnh2w7m9ga;
  wire [m0xuxgjqd7dh8v-1:0] hpkf4c2rxkqe4p = vf5xcr67bqhzlo43_[m0xuxgjqd7dh8v-1:0];
  ux607_gnrl_dfflr #(m0xuxgjqd7dh8v) soqj1k1jkdlr7341 (ybn5wo3zvbsf5, hpkf4c2rxkqe4p, b7iuqg01sm8apr[m0xuxgjqd7dh8v-1:0], gf33atgy, ru_wi);
  assign b7iuqg01sm8apr[64-1:m0xuxgjqd7dh8v] = {64-1-m0xuxgjqd7dh8v{1'b0}};

  genvar i;

  generate 
  for(i=0; i<4; i=i+1) begin: g790m7g1d8iw 
    assign n6a0r_0zddzrme8 [64*i +: 64] = qzr9ikzg_vz[i];
    assign azll7rq5fab5ou [64*i +: 64] = dwt4xr7nj[i];

    assign fv66706su4xcaxv[i] = (b7iuqg01sm8apr[m0xuxgjqd7dh8v-1:0] == i[m0xuxgjqd7dh8v-1:0]);

    
    
    
    
    assign rx3dpavi0xj7b4gx[i] = (p389kv4igf_ei2d[i] ? pydatzxqqi : 1'b1);
    assign bt36dhn0q97o3x[i] = da36aklh2x1yugbf & fv66706su4xcaxv[i] & rx3dpavi0xj7b4gx[i];
    assign dgv2oqmmc685v[i] = idm817wr_az479 & fv66706su4xcaxv[i] & rx3dpavi0xj7b4gx[i];

    
    ux607_gnrl_dfflr #(64) gvvtvabs3nnfc6z_ (dgv2oqmmc685v[i], vf5xcr67bqhzlo43_, qzr9ikzg_vz[i], gf33atgy, ru_wi);


    
    assign ornx_vnpekug3gz[i] = bt36dhn0q97o3x[i];
                               
    assign il72jv39takrecodwjg[i] = 
                              (vf5xcr67bqhzlo43_[64-1:64-4] == 4'd5) ? 4'd5 :
                              (vf5xcr67bqhzlo43_[64-1:64-4] == 4'd4) ? 4'd4 :
                              (vf5xcr67bqhzlo43_[64-1:64-4] == 4'd3) ? 4'd3 :
                                                                                          4'd2 ;
    ux607_gnrl_dfflr #(2) yyplgejg_5ga55oz0uxrgebse (ornx_vnpekug3gz[i], il72jv39takrecodwjg[i][3:2], l37vb0thqk484l[i][3:2], gf33atgy, ru_wi);
    ux607_gnrl_dfflrs#(1) ogv3oscqy5opmirmxiorf53_  (ornx_vnpekug3gz[i], il72jv39takrecodwjg[i][1]  , l37vb0thqk484l[i][1]  , gf33atgy, ru_wi);
    ux607_gnrl_dfflr #(1) kmp5rp3yt0k03ot72ney7   (ornx_vnpekug3gz[i], il72jv39takrecodwjg[i][0]  , l37vb0thqk484l[i][0]  , gf33atgy, ru_wi);

    assign lublr8yrk2iclyv1090[i] = (il72jv39takrecodwjg[i] == 4'd2);
    assign qytl9l30d1xwc77h3[i] = (il72jv39takrecodwjg[i] == 4'd3);
    assign ekcdji6jnpih8_4dk2tc[i] = (il72jv39takrecodwjg[i] == 4'd4);
    assign s4yy9maabthu6i_jf9svf8[i] = (il72jv39takrecodwjg[i] == 4'd5);

    
    assign ox0hspotahshker242[i] = (l37vb0thqk484l[i] == 4'd2);
    assign f_en44nuq7wxpi6[i] = (l37vb0thqk484l[i] == 4'd3);
    assign zdauex3dn6kp7jfh[i] = (l37vb0thqk484l[i] == 4'd4);
    assign lc7l4i7ez6dwylrrke[i] = (l37vb0thqk484l[i] == 4'd5);

    
    assign n24f03wv5exza5j6or0c[i] = bt36dhn0q97o3x[i] & pydatzxqqi;
    assign egctw8sjve74zbjm64f2[i] = vf5xcr67bqhzlo43_[59];
    ux607_gnrl_dfflr #(1) frig5b7l4n56lewyq5p2 (n24f03wv5exza5j6or0c[i], egctw8sjve74zbjm64f2[i], p389kv4igf_ei2d[i], gf33atgy, ru_wi);

    
    assign dlgms2ikbd24vp0r2[i] = bt36dhn0q97o3x[i];
    assign lsh9e8uas4hp15ahg1j[i] = vf5xcr67bqhzlo43_[64-6:0] & (
            
        ({59{lublr8yrk2iclyv1090[i]}} & {6'd12,{64-29{1'b0}},
                                                             (
                              
                                                                (vf5xcr67bqhzlo43_[17:12] == 6'd1) ? 6'd1 : 6'd0
                                                             ),
                              
                                                             1'b0,
                                                             (
                              
                                                                (vf5xcr67bqhzlo43_[10:7] == 4'd0) ? 4'd0 :
                                                                (vf5xcr67bqhzlo43_[10:7] == 4'd1) ? 4'd1 : 4'd0
                                                                
                                                             ),
                                                               vf5xcr67bqhzlo43_[6],1'b0,vf5xcr67bqhzlo43_[4:0]})
      | ({59{qytl9l30d1xwc77h3[i]}} & {16'b0,1'b1,vf5xcr67bqhzlo43_[9],1'b0,vf5xcr67bqhzlo43_[7:6],
                                                                ((vf5xcr67bqhzlo43_[5:0] == 6'd1) ? 6'd1 : 6'd0)
                                                       })
      | ({59{ekcdji6jnpih8_4dk2tc[i]}} & {17'b0,vf5xcr67bqhzlo43_[9],1'b0,vf5xcr67bqhzlo43_[7:6],
                                                                ((vf5xcr67bqhzlo43_[5:0] == 6'd1) ? 6'd1 : 6'd0)
                                                       })
      | ({59{s4yy9maabthu6i_jf9svf8[i]}} & {17'b0,vf5xcr67bqhzlo43_[9],1'b0,vf5xcr67bqhzlo43_[7:6],
                                                                ((vf5xcr67bqhzlo43_[5:0] == 6'd1) ? 6'd1 : 6'd0)
                                                       })
      );

    ux607_gnrl_dfflr #(17) colo12m11vnwsag00f4fj53a571 (dlgms2ikbd24vp0r2[i], lsh9e8uas4hp15ahg1j[i][26:10], hev3ez6yazmxe[i][26:10], gf33atgy, ru_wi);
    ux607_gnrl_dfflr #(6 ) kssplp2lxotz4r81g2v2fppo  (dlgms2ikbd24vp0r2[i], lsh9e8uas4hp15ahg1j[i][5:0], hev3ez6yazmxe[i][5:0], gf33atgy, ru_wi);
       
    assign  vr0xmfp80ka92vtnhtwvnuyf[i] =  f_en44nuq7wxpi6[i] & ns0i7siujgkrghjpqv6; 
    assign  mfu6jps217vim6x17jhy[i] =  vr0xmfp80ka92vtnhtwvnuyf[i] ? 4'b0 :  lsh9e8uas4hp15ahg1j[i][9:6];
    assign  m_44xky76stmh65migajp7t[i] =  dlgms2ikbd24vp0r2[i] | vr0xmfp80ka92vtnhtwvnuyf[i];
    ux607_gnrl_dfflr #(4 ) tc26_s2x710jwb0syvgu_  (m_44xky76stmh65migajp7t[i], mfu6jps217vim6x17jhy[i], hev3ez6yazmxe[i][9:6], gf33atgy, ru_wi);

    assign hev3ez6yazmxe[i][59-1:27] = {(59-27){1'b0}};
  
    assign cn5uuiza89o2dulas69s[i] = (
            
        ({59{ox0hspotahshker242[i]}} & {6'd12,{64-29{1'b0}},
                                                      (p389kv4igf_ei2d[i] ? hev3ez6yazmxe[i][17:12] : 6'b0),
                                                      hev3ez6yazmxe[i][11:6],1'b0,
                                                      hev3ez6yazmxe[i][4],
                                                      hev3ez6yazmxe[i][3],
                                                      hev3ez6yazmxe[i][2:0] 
                                                      })
      | ({59{f_en44nuq7wxpi6[i]}} & {{64-29{1'b0}},13'b0,1'b1,hev3ez6yazmxe[i][9],1'b0,
                                                       hev3ez6yazmxe[i][7],
                                                       hev3ez6yazmxe[i][6],
                                                      (p389kv4igf_ei2d[i] ? hev3ez6yazmxe[i][5:0] : 6'b0)
                                                      })
      | ({59{zdauex3dn6kp7jfh[i]}} & {{64-29{1'b0}},14'b0,hev3ez6yazmxe[i][9],1'b0,
                                                       hev3ez6yazmxe[i][7],
                                                       hev3ez6yazmxe[i][6],
                                                      (p389kv4igf_ei2d[i] ? hev3ez6yazmxe[i][5:0] : 6'b0)
                                                      })
      | ({59{lc7l4i7ez6dwylrrke[i]}} & {{64-29{1'b0}},14'b0,hev3ez6yazmxe[i][9],1'b0,
                                                       hev3ez6yazmxe[i][7],
                                                       hev3ez6yazmxe[i][6],
                                                      (p389kv4igf_ei2d[i] ? hev3ez6yazmxe[i][5:0] : 6'b0)
                                                      })
      );

    assign dwt4xr7nj[i][64-1:64-4]  = l37vb0thqk484l[i];
    assign dwt4xr7nj[i][59] = p389kv4igf_ei2d[i];
    assign dwt4xr7nj[i][64-6:0]  = cn5uuiza89o2dulas69s[i];

  end
  endgenerate

  wire [m0xuxgjqd7dh8v-1:0] gf912jyw6glbprc = b7iuqg01sm8apr[m0xuxgjqd7dh8v-1:0];

  assign rbz9x0m18nf7d = dwt4xr7nj[gf912jyw6glbprc];
  assign z585kaqlq5f76 = qzr9ikzg_vz[gf912jyw6glbprc];



    
    
    
  wire q9fnwgepl2uk = osv2437qj_3nuf;
  wire [3-1:0] dcause_r;
  wire [3-1:0] zbbv20bxclc7mjl = i8_5wt0vppx;
  ux607_gnrl_dfflr #(3) gkh85m21drzd0fr (q9fnwgepl2uk, zbbv20bxclc7mjl, dcause_r, gf33atgy, ru_wi);
    
      
    
  wire qby5u_h6 = b_a74a2_dk7xhm;
  wire xq5p8ehcqg;
  wire plzc96y6;
  assign xq5p8ehcqg = vf5xcr67bqhzlo43_[2];
  ux607_gnrl_dfflr #(1) t_i310u0fb (qby5u_h6, xq5p8ehcqg, plzc96y6, gf33atgy, ru_wi);


    
  wire tzaz1k4cxwwmr28 = b_a74a2_dk7xhm;
  wire zjhwvj30c7l;
  wire n0a_osbqkff;
  assign zjhwvj30c7l = vf5xcr67bqhzlo43_[4];
  ux607_gnrl_dfflr #(1) sa_cbp3qivatkd (tzaz1k4cxwwmr28, zjhwvj30c7l, n0a_osbqkff, gf33atgy, ru_wi);

    
  wire xavshexsg9 = b7g_vsn0zoewh6g1 | b_a74a2_dk7xhm;
  wire [1:0] x0d87zpapuh;
  wire [1:0] ybqoy9knv;
  assign x0d87zpapuh = b_a74a2_dk7xhm ? vf5xcr67bqhzlo43_[1:0] : onnv64ydiajl;
     
  ux607_gnrl_dfflrs #(2) yssxicr5do96 (xavshexsg9, x0d87zpapuh, ybqoy9knv, gf33atgy, ru_wi);
 

    
    
  wire nyi5c_a7hfs = b_a74a2_dk7xhm;
  wire roue5glh06;
  wire i_pf97_7p3nis;
  assign roue5glh06 = vf5xcr67bqhzlo43_[11];
  ux607_gnrl_dfflr #(1) aerxy166iuqq6bf (nyi5c_a7hfs, roue5glh06, i_pf97_7p3nis, gf33atgy, ru_wi);

    
    
  wire upm54surnxlhe = b_a74a2_dk7xhm;
  wire qkkq5bsx2v2t1qll;
  wire ft2e8rpvq9_;
  assign qkkq5bsx2v2t1qll = vf5xcr67bqhzlo43_[15];
  ux607_gnrl_dfflr #(1) kq1g1yb4j2fvkz (upm54surnxlhe, qkkq5bsx2v2t1qll, ft2e8rpvq9_, gf33atgy, ru_wi);
    
    
  wire uyj4r97taxpf = b_a74a2_dk7xhm;
  wire f1vwaiwj09do;
  wire c8bz9kbbc8;
  assign f1vwaiwj09do = vf5xcr67bqhzlo43_[13];
  ux607_gnrl_dfflr #(1) tqtdaw70fynpaat (uyj4r97taxpf, f1vwaiwj09do, c8bz9kbbc8, gf33atgy, ru_wi);
    
    
  wire r3m1693_gepr = b_a74a2_dk7xhm;
  wire ym009g80rgkalv_4;
  wire khktyrar6;
  assign ym009g80rgkalv_4 = vf5xcr67bqhzlo43_[12];
  ux607_gnrl_dfflr #(1) t4fxgvcy1k3nxx7 (r3m1693_gepr, ym009g80rgkalv_4, khktyrar6, gf33atgy, ru_wi);


    
  wire u_qb3lov3brow_ = b_a74a2_dk7xhm;
  wire gbm_t5wjkexqs3;
  wire f7gcid5pkp5m6kbu;
  assign gbm_t5wjkexqs3 = vf5xcr67bqhzlo43_[10];
  ux607_gnrl_dfflrs #(1) v_g5f1e841di9zx3oy (u_qb3lov3brow_, gbm_t5wjkexqs3, f7gcid5pkp5m6kbu, gf33atgy, ru_wi);
    
    
  wire j2d8mud9bbxku6yb_ = b_a74a2_dk7xhm;
  wire l9vyu9j2kf0m070;
  wire o51zp1lc_f0y;
  assign l9vyu9j2kf0m070 = vf5xcr67bqhzlo43_[9];
  ux607_gnrl_dfflrs #(1) gv2p5yqagu4y17d (j2d8mud9bbxku6yb_, l9vyu9j2kf0m070, o51zp1lc_f0y, gf33atgy, ru_wi);

generate
if (64 > 32) begin : aqsm5ybe48dcv
  assign dwns7g [64-1:32] = {64-32{1'b0}};
end
endgenerate

  assign dwns7g [15]  = ft2e8rpvq9_;
  assign dwns7g [14]  = 1'b0;
  assign dwns7g [13]  = c8bz9kbbc8;
  assign dwns7g [12]  = khktyrar6;

  assign dwns7g [10]    = f7gcid5pkp5m6kbu;
  assign dwns7g [9]     = o51zp1lc_f0y;
  assign dwns7g [8:6]   = dcause_r; 

  assign dwns7g [2]   = plzc96y6;
  assign dwns7g [1:0] = ybqoy9knv;

  assign dwns7g [31:28] = 4'd4;
  assign dwns7g [27:16]  = 12'b0;
  assign dwns7g [11]  = i_pf97_7p3nis;

  assign dwns7g [5]     = 1'b0;
  assign dwns7g [4]   = n0a_osbqkff;

  assign dwns7g [3]   = rn1o3sl83;

  assign ozwene1gdpatk6g = i_pf97_7p3nis;


  assign pydatzxqqi = ~(dcause_r == 3'b0);


  assign t5trf35s8vy = plzc96y6;
  assign zbac123pv78sbz3 = ft2e8rpvq9_;
  assign z4e_m564fxae0kpbjr = c8bz9kbbc8;
  assign hixy2y36a1pn0 = khktyrar6;
  assign r21i4by0bu3ks = ybqoy9knv;

  assign sxvvsxtbhyvt  = n0a_osbqkff ;


  assign zmwq3e9oijvo7d7 = f7gcid5pkp5m6kbu;
  assign q4gqhurcazjpsf4h  = pydatzxqqi & o51zp1lc_f0y;

endmodule





















module pulwy5sk17o3m9m6x (

  input  rb077g2alw88,
  input  kdnujwd70g0p,  
  input  yez0ldac23i95,
  input  gc4b3kdcan6do88ta_,


  input   idi3vfnshcpo,
  output  jzwasdy8fj0howe,
  output  a02zzbowpjn06h,
  input   um8zsjyxn_4p,

  input  v66uy2mvzfhls6,

  input  u_ll4hq1b12s2i1,
  input  w41ourymsjpvm8q1e,
  input  t4bp4v54b9fmhin,
  output truuny5aeeb6afbba,
  output dc8ehbd4k6bl2re764fz,
  input  i3cufk3oe15lxb_x,
  output q9x26ou3eg17z,
  output mzb743s60gk6mhj37sy,
  input  pom74hc61wlcgj8,
  output pik73_qshqijdw,
  output h9xe65iyw9qxvfp6,
  input  ndlpsbtthtn7hv,
  output v6pe_zs7a1rf5a,
  output dz3fwvx3e10_j6bfrgbzu,
  input  dlkg75fv,

  input  u6j3yp5u249c9in70r6h,
  input  pjy0x0i1ftpgz1lr_3dk,

  output io5ukym11gp2utw,
  output agsknykmgwpc,



  
  
    
  input rb050tnl,
  input a94vd35etec4,
  input el7_p8jit09,
  input [12-1:0] e1go3iu,
  input izhvh9xxvwe2,
  input  [64-1:0] vf5xcr67bqhzlo43_,
  output [64-1:0] l9erxxpnphqd26vg9,
  output u2dvoyt5e7o_03z9z5,
  output s904ol6a25v9zn8,

    
  input   [64-1:0] qeb3z0x5,
  input   ibhfuwrztbm8p4gg,

  input   [3-1:0] i8_5wt0vppx,
  input   osv2437qj_3nuf,



  input  b7g_vsn0zoewh6g1,
  input  [2-1:0] onnv64ydiajl,
  output [2-1:0] r21i4by0bu3ks,


  output [64*4-1:0] azll7rq5fab5ou,
  output [64*4-1:0] n6a0r_0zddzrme8,
  input  ns0i7siujgkrghjpqv6,


  output pydatzxqqi,
  output t5trf35s8vy,
  output zbac123pv78sbz3,
  output z4e_m564fxae0kpbjr,
  output zmwq3e9oijvo7d7,
  output q4gqhurcazjpsf4h ,

  output c5ewdqztjw9za,

  output hixy2y36a1pn0,
  output ozwene1gdpatk6g,
  output sxvvsxtbhyvt,
  input  rn1o3sl83,

  output [64-1:0] hn85hkp2yav,


  input              wex3zbl1x6s4be1en,
  input [1:0]        pszbl2iobld50k,   
  input              vfuu2l_7oof31qn0_a,   
  input [32-1:0] bvy9o58rgxtbjz_xph,    
  input [2:0]        gcpthp2sfxb3cxo,
  input [2:0]        xzjdk5deciqs4l3my_l,
  input [3:0]        peug05ptx4vv93u4xc, 
  input [64    -1:0] dlg9f36umgj9xdv0wa,   
  output [64    -1:0] yienty7ycnc25au,   
  output [1:0]        rxlx2eq69oye0ba3,    
  output              j2amhrzbhku8dzd,  

 
output                       fkm9up63o1aeauaqhjb,
input                        to_1lv9wnb3vmu6tvz5rc,
output [32-1:0] ju1kbeplcqy314lfj4, 
output                       r985fbe5k7hgzaq9i, 
output                       bb04gpwotp2s6c7_p1gqkq, 
output                       sqmey185cu3mtixhl, 
output                       rffcsd1o699ytclmx,
output  [64-1:0]     lbr88vbqtg8rht7320frde,
output  [8-1:0]  g7qq38mx3d58n1b15kcia,
output                       demg_fwfkmaeawq30t,
output                       grtb6ypa0px2gi1c,
output  [1:0]                f128d8ws0seoihu1,

input                        m2r7mfmq3afdd1ine,
output                       nhafiywg3hg_52kogwh,
input                        xrqayy6vigrw66z8a  ,
input                        jyy72ywt9nbo10f2jxupacld,
input [64-1:0]       drz92qecqx_qtxwro,
input                        st4f16aums5, 
input                        p05ld2ghmwh, 



  input   j_r1zrxno8j,
  input   kjc1hiyz 
);


  wire debugint;

  assign c5ewdqztjw9za = debugint;



  w0v8rrkl3p_ar0i2l u_ux607_dbg_csr (
    .rb050tnl         (rb050tnl       ),
    .a94vd35etec4       (a94vd35etec4     ),
    .el7_p8jit09       (el7_p8jit09     ),
    .e1go3iu         (e1go3iu       ),
    .izhvh9xxvwe2    (izhvh9xxvwe2  ),
    .vf5xcr67bqhzlo43_    (vf5xcr67bqhzlo43_  ),
    .l9erxxpnphqd26vg9    (l9erxxpnphqd26vg9  ),
    .u2dvoyt5e7o_03z9z5  (u2dvoyt5e7o_03z9z5),
    .s904ol6a25v9zn8    (s904ol6a25v9zn8),

    .qeb3z0x5         (qeb3z0x5        ),
    .ibhfuwrztbm8p4gg     (ibhfuwrztbm8p4gg    ),
    .i8_5wt0vppx      (i8_5wt0vppx     ),
    .osv2437qj_3nuf  (osv2437qj_3nuf ),



    .b7g_vsn0zoewh6g1    (b7g_vsn0zoewh6g1),
    .onnv64ydiajl        (onnv64ydiajl    ),
    .r21i4by0bu3ks       (r21i4by0bu3ks   ),

    .azll7rq5fab5ou      (azll7rq5fab5ou),
    .n6a0r_0zddzrme8      (n6a0r_0zddzrme8),
    .ns0i7siujgkrghjpqv6(ns0i7siujgkrghjpqv6),

    .hixy2y36a1pn0   (hixy2y36a1pn0),
    .ozwene1gdpatk6g      (ozwene1gdpatk6g   ),
    .sxvvsxtbhyvt      (sxvvsxtbhyvt   ),
    .rn1o3sl83       (rn1o3sl83    ),

                                     
    .zmwq3e9oijvo7d7   (zmwq3e9oijvo7d7),
    .q4gqhurcazjpsf4h    (q4gqhurcazjpsf4h ),
    .pydatzxqqi        (pydatzxqqi),
    .t5trf35s8vy      (t5trf35s8vy),
    .zbac123pv78sbz3   (zbac123pv78sbz3),
    .z4e_m564fxae0kpbjr   (z4e_m564fxae0kpbjr),
    .hn85hkp2yav       (hn85hkp2yav),

    .gf33atgy             (j_r1zrxno8j),
    .ru_wi           (kjc1hiyz) 
  );





  wire  go6srylfev;
  wire  tydimrd3y69;
  wire  k9795draeeio5ksrbt = um8zsjyxn_4p & (~pjy0x0i1ftpgz1lr_3dk);

  wire g7wai968_xx8y = jzwasdy8fj0howe & (~k9795draeeio5ksrbt);
  
  wire yb121j9cq = (~k9795draeeio5ksrbt);

  
  ux607_clkgate jc7hbz4i19s8b(
    .clk_in   (idi3vfnshcpo    ),
    .clkgate_bypass(gc4b3kdcan6do88ta_  ),
    .clock_en (g7wai968_xx8y),
    .clk_out  (go6srylfev)
  );

  
  ux607_clkgate fin1qva3k2k4d(
    .clk_in   (idi3vfnshcpo    ),
    .clkgate_bypass(gc4b3kdcan6do88ta_  ),
    .clock_en (yb121j9cq),
    .clk_out  (tydimrd3y69)
  );


  wire na29rv9xyz_vn;
  wire dfnv8e05y_xxox4kof;

  ux607_reset_sync v0cqe_z_nwx1n04h697ap3 (
    .clk      (dlkg75fv),
    .rst_n_a  (kdnujwd70g0p),
    .reset_bypass(yez0ldac23i95),
    .rst_n_sync(dfnv8e05y_xxox4kof) 
  );

  ux607_reset_sync ufowdnwj6d3ociy0_x8betoh (
    .clk      (idi3vfnshcpo),
    .rst_n_a  (kdnujwd70g0p),
    .reset_bypass(yez0ldac23i95),
    .rst_n_sync(na29rv9xyz_vn) 
  );

  wire s69lpiuwzwxu_;
  wire sqvy97shfxgalqcq;
  
  
  wire uapa77w9uuj_t9p = yez0ldac23i95 ? kdnujwd70g0p : s69lpiuwzwxu_;

  ux607_reset_sync fuiavtxj5adoss0hla00p (
    .clk      (idi3vfnshcpo),
    .rst_n_a  (uapa77w9uuj_t9p), 
    .reset_bypass(yez0ldac23i95),
    .rst_n_sync(sqvy97shfxgalqcq) 
  );


  wire o59nl09azxaz;

  b7e3qelmq5qz ir87ykicng (
      .o59nl09azxaz              (o59nl09azxaz),
      .um8zsjyxn_4p             (k9795draeeio5ksrbt),

      .s69lpiuwzwxu_           (s69lpiuwzwxu_    ),
      .sqvy97shfxgalqcq       (sqvy97shfxgalqcq),
      .a02zzbowpjn06h        (a02zzbowpjn06h),
	  .o0pri6gw33y              (debugint        ), 
	  .z5w8jrogg064jr           (pydatzxqqi        ),
	  .u_ll4hq1b12s2i1          (u_ll4hq1b12s2i1    ),
	  .w41ourymsjpvm8q1e      (w41ourymsjpvm8q1e),
	  .t4bp4v54b9fmhin           (t4bp4v54b9fmhin), 
	  .truuny5aeeb6afbba          (truuny5aeeb6afbba),
	  .dc8ehbd4k6bl2re764fz       (dc8ehbd4k6bl2re764fz),
	  .i3cufk3oe15lxb_x           (i3cufk3oe15lxb_x),
	  .q9x26ou3eg17z          (q9x26ou3eg17z), 
	  .mzb743s60gk6mhj37sy       (mzb743s60gk6mhj37sy ), 
	  .pom74hc61wlcgj8           (pom74hc61wlcgj8), 
	  .pik73_qshqijdw          (pik73_qshqijdw),
	  .h9xe65iyw9qxvfp6       (h9xe65iyw9qxvfp6), 
	  .ndlpsbtthtn7hv          (ndlpsbtthtn7hv), 
	  .v6pe_zs7a1rf5a         (v6pe_zs7a1rf5a), 
	  .dz3fwvx3e10_j6bfrgbzu      (dz3fwvx3e10_j6bfrgbzu),
	  .go89gmq               (dlkg75fv), 
	  .hfocw7va5_               (1'b0), 
	  .io5ukym11gp2utw          (io5ukym11gp2utw), 
	  .obvunz7               (tydimrd3y69), 
    .v66uy2mvzfhls6     (v66uy2mvzfhls6),
      .dfnv8e05y_xxox4kof         (dfnv8e05y_xxox4kof),
      .na29rv9xyz_vn         (na29rv9xyz_vn),
      .yez0ldac23i95          (yez0ldac23i95),
	  .agsknykmgwpc          (agsknykmgwpc), 
	  .bmm03who3rv              (idi3vfnshcpo      ), 
	  .wivo                  (go6srylfev           ), 
	  .fkm9up63o1aeauaqhjb     (fkm9up63o1aeauaqhjb ),
	  .to_1lv9wnb3vmu6tvz5rc     (to_1lv9wnb3vmu6tvz5rc ),
	  .ju1kbeplcqy314lfj4      (ju1kbeplcqy314lfj4  ), 
	  .r985fbe5k7hgzaq9i      (r985fbe5k7hgzaq9i  ), 
	  .bb04gpwotp2s6c7_p1gqkq     (bb04gpwotp2s6c7_p1gqkq ), 
	  .sqmey185cu3mtixhl     (sqmey185cu3mtixhl ), 
	  .rffcsd1o699ytclmx     (rffcsd1o699ytclmx ),
	  .lbr88vbqtg8rht7320frde     (lbr88vbqtg8rht7320frde ),
	  .g7qq38mx3d58n1b15kcia     (g7qq38mx3d58n1b15kcia ),
	  .demg_fwfkmaeawq30t      (demg_fwfkmaeawq30t  ),
	  .grtb6ypa0px2gi1c      (grtb6ypa0px2gi1c  ),
	  .f128d8ws0seoihu1      (f128d8ws0seoihu1  ),
	  .m2r7mfmq3afdd1ine     (m2r7mfmq3afdd1ine ),
	  .nhafiywg3hg_52kogwh     (nhafiywg3hg_52kogwh ),
	  .xrqayy6vigrw66z8a       (xrqayy6vigrw66z8a   ),
	  .jyy72ywt9nbo10f2jxupacld   (jyy72ywt9nbo10f2jxupacld),
	  .drz92qecqx_qtxwro     (drz92qecqx_qtxwro ),
	  .st4f16aums5             (st4f16aums5         ), 
	  .p05ld2ghmwh             (p05ld2ghmwh         ), 
	  .tk2pf9erp83             (1'b1              ), 
	  .p9_huoh6oy1jai           (pszbl2iobld50k    ), 
	  .ohod7vxvej8qwj           (vfuu2l_7oof31qn0_a    ), 
	  .evqksuwcgvwotl            (bvy9o58rgxtbjz_xph     ), 
	  .qbiibzbu0j5xu            (gcpthp2sfxb3cxo     ), 
	  .re6g_r1kz98u           (xzjdk5deciqs4l3my_l    ), 
	  .fa9ntbvuu_3cuqr5           (dlg9f36umgj9xdv0wa    ), 
	  .l88j4b6ovz            (peug05ptx4vv93u4xc     ), 
	  .coiuburq3cf           (yienty7ycnc25au    ), 
	  .n2vqwxz4b7yahnp           (j2amhrzbhku8dzd    ), 
	  .v5jhtjwnqklb6oje85        (j2amhrzbhku8dzd    ), 
	  .lzl17_6p6y91nh            (rxlx2eq69oye0ba3     )  

);


  assign jzwasdy8fj0howe = (~u6j3yp5u249c9in70r6h) & (
                                     o59nl09azxaz       |
                                     a02zzbowpjn06h | 
                                     wex3zbl1x6s4be1en  
                                 );




endmodule


module b7e3qelmq5qz (
input                        um8zsjyxn_4p,
output                       o59nl09azxaz,
output                       s69lpiuwzwxu_,
input                        sqvy97shfxgalqcq,
output                       a02zzbowpjn06h,
output                       o0pri6gw33y,
input                        z5w8jrogg064jr,
input                        u_ll4hq1b12s2i1,
input                        w41ourymsjpvm8q1e,
input                        t4bp4v54b9fmhin,
output                       truuny5aeeb6afbba,
output                       dc8ehbd4k6bl2re764fz,
input                        i3cufk3oe15lxb_x,
output                       q9x26ou3eg17z,
output                       mzb743s60gk6mhj37sy,
input                        pom74hc61wlcgj8,
output                       pik73_qshqijdw,
output                       h9xe65iyw9qxvfp6,
input                        ndlpsbtthtn7hv,
output                       v6pe_zs7a1rf5a,
output                       dz3fwvx3e10_j6bfrgbzu,
input                        hfocw7va5_,
output                       io5ukym11gp2utw,
input                        obvunz7,                    
input                        go89gmq,                 
input                        dfnv8e05y_xxox4kof,
input                        na29rv9xyz_vn,
input                        yez0ldac23i95 ,
output                       agsknykmgwpc,
input                        bmm03who3rv,
input                        wivo,
 
output                       fkm9up63o1aeauaqhjb,
input                        to_1lv9wnb3vmu6tvz5rc,
output [32-1:0] ju1kbeplcqy314lfj4, 
output                       r985fbe5k7hgzaq9i, 
output                       bb04gpwotp2s6c7_p1gqkq, 
output                       sqmey185cu3mtixhl, 
output                       rffcsd1o699ytclmx,
output  [64-1:0]     lbr88vbqtg8rht7320frde,
output  [8-1:0]  g7qq38mx3d58n1b15kcia,
output                       demg_fwfkmaeawq30t,
output                       grtb6ypa0px2gi1c,
output  [1:0]                f128d8ws0seoihu1,

input                        m2r7mfmq3afdd1ine,
output                       nhafiywg3hg_52kogwh,
input                        xrqayy6vigrw66z8a  ,
input                        jyy72ywt9nbo10f2jxupacld,
input [64-1:0]       drz92qecqx_qtxwro,
input                        st4f16aums5, 
input                        p05ld2ghmwh, 
input  v66uy2mvzfhls6,
input  [32-1:0] evqksuwcgvwotl,
input                  [2:0] re6g_r1kz98u,
input                  [3:0] l88j4b6ovz,
output      [64-1:0] coiuburq3cf,
input                        n2vqwxz4b7yahnp,
output                       v5jhtjwnqklb6oje85,
output                 [1:0] lzl17_6p6y91nh,
input                        tk2pf9erp83,
input                  [2:0] qbiibzbu0j5xu,
input                  [1:0] p9_huoh6oy1jai,
input       [64-1:0] fa9ntbvuu_3cuqr5,
input                        ohod7vxvej8qwj

);

localparam yv13_lx8u9yhr8p6i	= 8;

localparam smfpyk6 = 1;


wire             [smfpyk6-1:0] eb7x00xzyu84l5;
wire             [smfpyk6-1:0] su_naptw5zy82_smisyx;
wire             [smfpyk6-1:0] aktp_d2l4ho7n9w315xuy;
wire                   [8:0] v0ppt_lszz;
wire                         liu_rgb4nf;
wire                         jfyllx;
wire                         a9c;
wire                  [31:0] yav2e_pam99eaw3okf7;
wire                   [2:0] tfljpdijxf;
wire                   [3:0] c98a8jw632g1;
wire                         m82k9gnjrw;
wire                         gtvu1jhq;
wire                   [2:0] naonfp5kwul39;
wire                   [1:0] lpv3w7_jux0x5;
wire                  [31:0] j8tyg8pg_v_hj12;
wire                         iw4viufqn3;
wire                         hmb;
wire                         qfuuzymrquo;
wire             [smfpyk6-1:0] ns7mo9vqtdv3x;
wire             [smfpyk6-1:0] q1yf3ldhtd59mjj;
wire                  [31:0] eplm38kc000z;
wire                         hj3v8ja2n1snk;
wire                   [1:0] u8hp_cxp52qsad4yus;

assign v0ppt_lszz = yav2e_pam99eaw3okf7[8:0];
assign liu_rgb4nf = u8hp_cxp52qsad4yus[0];
assign	v6pe_zs7a1rf5a	= 1'b0;		
assign	dz3fwvx3e10_j6bfrgbzu	= 1'b0;		
assign	a9c		= pom74hc61wlcgj8;
assign	truuny5aeeb6afbba	= 1'b0;
assign	dc8ehbd4k6bl2re764fz	= 1'b0;
assign	mzb743s60gk6mhj37sy	= qfuuzymrquo;
assign	h9xe65iyw9qxvfp6	= 1'b0;
assign	pik73_qshqijdw	= 1'b0;
assign	jfyllx		= t4bp4v54b9fmhin;
assign	q9x26ou3eg17z	= hmb;
assign su_naptw5zy82_smisyx[0]     = u_ll4hq1b12s2i1;
assign aktp_d2l4ho7n9w315xuy[0] = w41ourymsjpvm8q1e;
assign eb7x00xzyu84l5[0]      = z5w8jrogg064jr;
assign o0pri6gw33y = ns7mo9vqtdv3x[0];
assign io5ukym11gp2utw = q1yf3ldhtd59mjj[0];












gc116p0_4d #(
	.pbftactqbw8     (32 ),
	.vmw6vavuv7md5     (64      ),
	.smfpyk6          (smfpyk6           ),
	.yv13_lx8u9yhr8p6i   (yv13_lx8u9yhr8p6i    ),
	.ph9yy86osx2krs_e_ (9               )
 ) gc116p0_4d (
	.o0pri6gw33y        (ns7mo9vqtdv3x        ), 
	.io5ukym11gp2utw    (q1yf3ldhtd59mjj    ), 
	.o59nl09azxaz        (o59nl09azxaz           ), 
	.nm83rtc_qty        (agsknykmgwpc       ), 

	.dk2xhkj77a         (bmm03who3rv           ), 
	.gf33atgy             (wivo               ), 
	.hfocw7va5_         (sqvy97shfxgalqcq    ), 
    .v66uy2mvzfhls6     (v66uy2mvzfhls6),

	.u_ll4hq1b12s2i1    (su_naptw5zy82_smisyx    ), 
	.z5w8jrogg064jr     (eb7x00xzyu84l5     ), 
	.w41ourymsjpvm8q1e(aktp_d2l4ho7n9w315xuy), 
	.evqksuwcgvwotl      (evqksuwcgvwotl         ), 
	.p9_huoh6oy1jai     (p9_huoh6oy1jai        ), 
	.ohod7vxvej8qwj     (ohod7vxvej8qwj        ), 
	.qbiibzbu0j5xu      (qbiibzbu0j5xu         ), 
	.re6g_r1kz98u     (re6g_r1kz98u        ), 
	.l88j4b6ovz      (l88j4b6ovz         ), 
	.fa9ntbvuu_3cuqr5     (fa9ntbvuu_3cuqr5        ), 
	.tk2pf9erp83       (tk2pf9erp83          ), 
	.n2vqwxz4b7yahnp     (n2vqwxz4b7yahnp        ), 
	.coiuburq3cf     (coiuburq3cf        ), 
	.v5jhtjwnqklb6oje85  (v5jhtjwnqklb6oje85     ), 
	.lzl17_6p6y91nh      (lzl17_6p6y91nh         ), 
	.fkm9up63o1aeauaqhjb (fkm9up63o1aeauaqhjb),
	.to_1lv9wnb3vmu6tvz5rc (to_1lv9wnb3vmu6tvz5rc),
	.ju1kbeplcqy314lfj4  (ju1kbeplcqy314lfj4 ), 
	.r985fbe5k7hgzaq9i  (r985fbe5k7hgzaq9i ), 
	.bb04gpwotp2s6c7_p1gqkq (bb04gpwotp2s6c7_p1gqkq), 
	.sqmey185cu3mtixhl (sqmey185cu3mtixhl), 
	.rffcsd1o699ytclmx (rffcsd1o699ytclmx),
	.lbr88vbqtg8rht7320frde (lbr88vbqtg8rht7320frde),
	.g7qq38mx3d58n1b15kcia (g7qq38mx3d58n1b15kcia),
	.demg_fwfkmaeawq30t  (demg_fwfkmaeawq30t ),
	.grtb6ypa0px2gi1c  (grtb6ypa0px2gi1c ),
	.f128d8ws0seoihu1  (f128d8ws0seoihu1 ),
	.m2r7mfmq3afdd1ine (m2r7mfmq3afdd1ine),
	.nhafiywg3hg_52kogwh (nhafiywg3hg_52kogwh),
	.xrqayy6vigrw66z8a   (xrqayy6vigrw66z8a  ),
	.jyy72ywt9nbo10f2jxupacld(jyy72ywt9nbo10f2jxupacld),
	.drz92qecqx_qtxwro (drz92qecqx_qtxwro),
	.st4f16aums5         (st4f16aums5        ), 
	.p05ld2ghmwh         (p05ld2ghmwh        ), 
	.ehdeq25ha       (v0ppt_lszz          ), 
	.hy7ogyog4pk_4i      (lpv3w7_jux0x5         ),
	.e_pz9vwnoa1r523      (iw4viufqn3         ),
	.o6807ghxyyt       (naonfp5kwul39          ),
	.wjddp1ply5kikfy      (tfljpdijxf         ),
	.x8m46uwduh       (c98a8jw632g1          ),
	.ph7jz_7_o_welqv      (j8tyg8pg_v_hj12         ),
	.jutj9q2kpi        (gtvu1jhq           ),
	.nrxv3rneu2438      (m82k9gnjrw         ),
	.tigza5anv0i48c7      (eplm38kc000z         ),
	.f2r3r2mwmdler   (hj3v8ja2n1snk      ),
	.o4hlkc18armddz       (u8hp_cxp52qsad4yus     ) 
); 

d6pt7ab0 d6pt7ab0 (
    .um8zsjyxn_4p    (um8zsjyxn_4p),
	.sqvy97shfxgalqcq(sqvy97shfxgalqcq),
    .a02zzbowpjn06h(a02zzbowpjn06h),

	.uecloq2rb    (1'b0           ), 
    .dfnv8e05y_xxox4kof(dfnv8e05y_xxox4kof),
    .na29rv9xyz_vn(na29rv9xyz_vn),
    .yez0ldac23i95 (yez0ldac23i95 ),
	.qzy          (go89gmq        ), 
	.a9c          (a9c            ), 
	.jfyllx          (jfyllx            ), 
	.hmb          (hmb            ), 
	.qfuuzymrquo   (qfuuzymrquo     ), 
	.lr4pmtw0e3sm7  (s69lpiuwzwxu_    ), 
	.bmm03who3rv     (bmm03who3rv       ), 
	.obvunz7      (obvunz7        ), 
	.d5gddvhozc     (wivo           ), 
	.gtvu1jhq     (gtvu1jhq       ), 
	.lpv3w7_jux0x5   (lpv3w7_jux0x5     ), 
	.v0ppt_lszz    (yav2e_pam99eaw3okf7), 
	.naonfp5kwul39    (naonfp5kwul39      ), 
	.tfljpdijxf   (tfljpdijxf     ), 
	.c98a8jw632g1    (c98a8jw632g1      ), 
	.j8tyg8pg_v_hj12   (j8tyg8pg_v_hj12     ), 
	.iw4viufqn3   (iw4viufqn3     ), 
	.eplm38kc000z   (eplm38kc000z     ), 
	.m82k9gnjrw   (hj3v8ja2n1snk  ), 
	.hj3v8ja2n1snk(m82k9gnjrw     ), 
	.liu_rgb4nf    (liu_rgb4nf      )  
); 


endmodule


module u_j2imkw7hy7 # (
    parameter vv3o1dwe8bt1m3k  = 32,
    parameter b4ff6gp7ae52l  = 7,
    parameter opmj43kpf6ptzium    = 2,
    parameter y76n53l844691b1v   = 41
  ) (

input                      yg8hetdkahah,
output  [31:0]             w4l6em1v0os9uky,
output                     lb2ioj3kfjgks,
input                      kvdg06d7vo7wv_n,
input   [y76n53l844691b1v-1:0] nmmjpe9w4mnr,
input                      wivo,
input                      zy4t8o4ibj,
input                      oyn5mkpu,
input   [31:0]             y7ftxl,
output                     n1xcixngo_e,
output  [31:0]             rw9vqyx,
output  [1:0]              mhayix,
output                     ad5i86r,
output  [2:0]              tihusk1,
output  [2:0]              abdy0h,
output  [3:0]              awm5ntb_,
output  [31:0]             t6tpgz13_m,
output                     l4pt3
);







localparam   p0t159zwkkyyulx         = 2'b00;
localparam   kapv0q86iup         = 2'b01;
localparam   yp4a2mouig8o9p2_i       = 2'b10;
localparam   jix2wlz5mjjui          = 2'b11;


localparam   mu74phcds4ei3            = 1'b0;
localparam   w6r9rhsqy8sa         = 1'b1;


localparam   ao_qx1lk8t0mh5c          = 2'b00;
localparam   y2w_s42cf6_94         = 2'b01;
localparam   ie_kg74b_wufbrz        = 2'b10;
localparam   yz80u836w74tl          = 2'b11;



wire	p3d97xkgvdmgxtyr6;


wire [y76n53l844691b1v-1:0]	umqf1s212fg;



wire	[1:0]	ucxte_5zd7;



wire 	ueon0c51941rhih3;


wire	s1r5jw3oqi6oylzkyss;
wire	s712q5omiiqjjjk10h;





wire	[b4ff6gp7ae52l-1:0]	er_y8yvk;

assign	p3d97xkgvdmgxtyr6 = oyn5mkpu & kvdg06d7vo7wv_n & ~lb2ioj3kfjgks & ~s1r5jw3oqi6oylzkyss & (mhayix == p0t159zwkkyyulx);
assign	er_y8yvk	     = umqf1s212fg[y76n53l844691b1v-1:(vv3o1dwe8bt1m3k+opmj43kpf6ptzium)];

assign	rw9vqyx        = {{(30-b4ff6gp7ae52l){1'b0}}, er_y8yvk, 2'b0};
assign	ad5i86r       = (umqf1s212fg[opmj43kpf6ptzium-1:0] == ie_kg74b_wufbrz);
assign	n1xcixngo_e    = oyn5mkpu;
assign	tihusk1        = 3'b010;		
assign	abdy0h       = 3'b000;		
assign	awm5ntb_        = 4'b0001;		
assign	t6tpgz13_m       = umqf1s212fg[(vv3o1dwe8bt1m3k+opmj43kpf6ptzium)-1:opmj43kpf6ptzium];
assign	l4pt3         = 1'b1;

assign	ucxte_5zd7 = p3d97xkgvdmgxtyr6 ? yp4a2mouig8o9p2_i : p0t159zwkkyyulx;

ux607_gnrl_dffr #(2) kxn38gfbl3 (ucxte_5zd7 , mhayix, wivo, yg8hetdkahah);













wire	sbtoy62g0fcmt0;

assign	sbtoy62g0fcmt0 = p3d97xkgvdmgxtyr6;

ux607_gnrl_dfflr #(y76n53l844691b1v)    ir9d3sa029k2sbxvy  (sbtoy62g0fcmt0, nmmjpe9w4mnr, umqf1s212fg, wivo, yg8hetdkahah);













wire	hrfypoiq5jcgwox3dc9f;
wire	t3es8qo4cjnyo2p8orh;
wire	q5sql6hopsvr6puo;
wire	xfiijy4o038yi5e_x;

assign	hrfypoiq5jcgwox3dc9f = (mhayix == yp4a2mouig8o9p2_i);
assign	t3es8qo4cjnyo2p8orh = (ueon0c51941rhih3 & oyn5mkpu) | ~kvdg06d7vo7wv_n;
assign	q5sql6hopsvr6puo = hrfypoiq5jcgwox3dc9f | t3es8qo4cjnyo2p8orh;
assign	xfiijy4o038yi5e_x = hrfypoiq5jcgwox3dc9f & ~t3es8qo4cjnyo2p8orh;

ux607_gnrl_dfflr #(1)    t5ie1n0quhg3hqyilz  (q5sql6hopsvr6puo, xfiijy4o038yi5e_x, ueon0c51941rhih3, wivo, yg8hetdkahah);













wire	kk5b5w_v4k0tql0s810yqwk;
assign	kk5b5w_v4k0tql0s810yqwk = s1r5jw3oqi6oylzkyss & ~ad5i86r & (zy4t8o4ibj == mu74phcds4ei3);

ux607_gnrl_dfflr #(32)    m7i1e5sg0z17inz5n5mgeou  (kk5b5w_v4k0tql0s810yqwk, y7ftxl, w4l6em1v0os9uky, wivo, yg8hetdkahah);













wire	qq7p0nantrfgkpx4so;
wire	jou_2cmm19pg1944iq;

assign	s1r5jw3oqi6oylzkyss = ueon0c51941rhih3 & oyn5mkpu;
assign	s712q5omiiqjjjk10h = ~kvdg06d7vo7wv_n;
assign	qq7p0nantrfgkpx4so = s1r5jw3oqi6oylzkyss | s712q5omiiqjjjk10h;
assign	jou_2cmm19pg1944iq = s1r5jw3oqi6oylzkyss & ~s712q5omiiqjjjk10h;

ux607_gnrl_dfflr #(1)    ruo1ok3sywvulyllrebeb  (qq7p0nantrfgkpx4so, jou_2cmm19pg1944iq, lb2ioj3kfjgks, wivo, yg8hetdkahah);















endmodule

module gc116p0_4d # (
  parameter pbftactqbw8     = 32,
  parameter vmw6vavuv7md5     = 32,
  parameter ph9yy86osx2krs_e_ = 9,
  parameter yv13_lx8u9yhr8p6i   = 2,
  parameter smfpyk6          = 1
 ) (
output [smfpyk6-1:0]          o0pri6gw33y,
output [smfpyk6-1:0]          io5ukym11gp2utw,
output                      o59nl09azxaz,
output                      nm83rtc_qty,
input                       dk2xhkj77a,
input                       gf33atgy,
input                       hfocw7va5_,
input  v66uy2mvzfhls6,
input  [smfpyk6-1:0]          u_ll4hq1b12s2i1,
input  [smfpyk6-1:0]          z5w8jrogg064jr,
input  [smfpyk6-1:0]          w41ourymsjpvm8q1e,

input  [pbftactqbw8-1:0]     evqksuwcgvwotl,
input  [1:0]                p9_huoh6oy1jai,
input                       ohod7vxvej8qwj,
input  [2:0]                qbiibzbu0j5xu,
input  [2:0]                re6g_r1kz98u,
input  [3:0]                l88j4b6ovz,
input  [vmw6vavuv7md5-1:0]     fa9ntbvuu_3cuqr5,
input                       tk2pf9erp83,
input                       n2vqwxz4b7yahnp,
output [vmw6vavuv7md5-1:0]     coiuburq3cf,
output                      v5jhtjwnqklb6oje85,
output [1:0]                lzl17_6p6y91nh, 
		  
		  
		  
		  
		  
		  
		  
		  
		  
		  
		  
		  
		  
		  
		  
		  
		  
		  
		  
		  
		  
		  
		  
		  
		  
		  
		  
		  
		  
		  
		  
		  
		  
		  
		  
		  
		  
		  
		  
		  
		  
		  
		  
		  
		  
		  
		  
		  
		  
		  
		  
		  
		  
		  
		  
		  
		  
		  
		  
		  
		  
		  
		  
		  
		  
		  
		  
		  
		  
		  
		  
		  
		  
		  
		  
		  
		  
		  
		  
		  
		  
		  
 
output                         fkm9up63o1aeauaqhjb,
input                          to_1lv9wnb3vmu6tvz5rc,
output [32-1:0]   ju1kbeplcqy314lfj4, 
output                         r985fbe5k7hgzaq9i, 
output                         bb04gpwotp2s6c7_p1gqkq, 
output                         sqmey185cu3mtixhl, 
output                         rffcsd1o699ytclmx,
output  [64-1:0]       lbr88vbqtg8rht7320frde,
output  [8-1:0]    g7qq38mx3d58n1b15kcia,
output                         demg_fwfkmaeawq30t,
output                         grtb6ypa0px2gi1c,
output  [1:0]                  f128d8ws0seoihu1,

input                          m2r7mfmq3afdd1ine,
output                         nhafiywg3hg_52kogwh,
input                          xrqayy6vigrw66z8a  ,
input                          jyy72ywt9nbo10f2jxupacld,
input [64-1:0]         drz92qecqx_qtxwro,
input                          st4f16aums5, 
input                          p05ld2ghmwh, 

input  [ph9yy86osx2krs_e_-1:0] ehdeq25ha,
input  [1:0]                hy7ogyog4pk_4i,
input                       e_pz9vwnoa1r523,
input  [2:0]                o6807ghxyyt,
input  [2:0]                wjddp1ply5kikfy,
input  [3:0]                x8m46uwduh,
input  [31:0]               ph7jz_7_o_welqv,
input                       jutj9q2kpi,
input                       nrxv3rneu2438,
output [31:0]               tigza5anv0i48c7,
output                      f2r3r2mwmdler,
output [1:0]                o4hlkc18armddz
);




parameter uaue4a0q4yu2u48 = 32;
parameter x5jl_73d_gruzgtcqu = 64;







parameter qibbagx75v9uch1w49v2yl5xd1se = "oq2da";
parameter s_hrmp88w3m_7k29y  = "uci2r";

parameter x2wextn4bicpd  = 4;
parameter gw_ey3om395hy = 4;


localparam d8panmbslrc4xeco = 4;       





























































































































localparam phi_3fuvuxlyqs28nm8 = 7'h00;
localparam bt42zx62uwdszqwoqv = 7'h01;
localparam yx886qndzla86sdd_3cv = 7'h02;
localparam dy4oanpu6e5ul1fz7g_ = 7'h03;
localparam odd20qdqw01usps7p = 7'h04;
localparam xw979wmvqaobuhc0xu3vb = 7'h05;
localparam ym_kkhyp5tltm8rtzye = 7'h06;
localparam l3hexpenpx19ve078w = 7'h07;
localparam w63v5w78bfszaqrq = 7'h08;
localparam bdjh2vk2nsr38k7_dngtl = 7'h09;
localparam ht9mdevmmqxwsbsnmoa = 7'h0a;
localparam g09ysbyxrmfbvydajmr6s = 7'h0b;
localparam i8eo0stsft_hj2hrc8 = 7'h0c;
localparam r63v9p0qtxpyxtfgzt6yd = 7'h0d;
localparam ox5a66g9lxe_7vmqmym79 = 7'h0e;
localparam fhpsm86w5w5gn25c9cy = 7'h0f;
localparam ux0b_d7_h0i9zgz5 = 7'h10;
localparam ijaa7ha3lixqhv_6d1pxf = 7'h11;
localparam obz94v8d60oebiebh = 7'h12;
localparam p8wxdxzfp4knovegq65 = 7'h13;
localparam ndu6q4dkyhmrc9g4w_t1 = 7'h14;
localparam gnuq76_e1vji_tt3x = 7'h15;
localparam tahrnunnmc14y7js = 7'h16;
localparam wgmilq0vnwlipd95z9n = 7'h17;

localparam wjwm0mmb8kdtc38hmvxcg7    = 7'h10; 
localparam jcqkgadqjnp1br60kcm7     = 7'h11; 
localparam r9pqyndxl9ydaeube81umk     = 7'h12; 
localparam dakqe9s6bwbckfsw4zlpj     = 7'h13; 
localparam aon_4_u6h74hgk3ispa3if13  = 7'h14; 
localparam aufn2qiboj8l12dufk0p     = 7'h15; 
localparam xpf4_70tcyabeblxkt7aob2y   = 7'h16; 
localparam bcei3m4eneqv0kswce_6      = 7'h17; 
localparam rzuyw47p7ehj1uy43z4w9l63d3 = 7'h18; 
localparam yi9jeqslby_o_kzsjsm3  = 7'h19; 
localparam wu726eflupgjm7hs9uonaad7p  = 7'h1a; 
localparam js76iv7t9nvkn6yv_4661  = 7'h1b; 
localparam fufl25ug_h3jqm3k9o_gkyii  = 7'h1c; 

localparam ggr6ql2zj7x40114w        = 7'h04; 
localparam tcnwfsqopcq2kj        = 7'h05; 
localparam ab_j1frhbffg57rc        = 7'h06; 
localparam jim0ddiqnav_mr        = 7'h07; 

localparam m0jpn5dn80dsf2q        = 7'h08; 
localparam zxe9_q2s5fzxgu_k38        = 7'h09; 
localparam va10rh7n02nkb6        = 7'h0a; 
localparam dmgo2idd7_vdsdnnaq3        = 7'h0b; 
localparam jbtj7er6n1t919tqlx        = 7'h0c; 
localparam qz57tyn0hruiw2xcq        = 7'h0d; 
localparam kfpiwe2xk_8vve0       = 7'h0e; 
localparam esrb21vaoahytvbimz       = 7'h0f; 
localparam u_cztegv7294f0w2ck     = 7'h20; 
localparam ew_k_8affyv8ltn2n9t     = 7'h21; 
localparam c2pgc56ortybp6qk31tah2     = 7'h22; 
localparam vojasz8wlqnrlmd7irtxe     = 7'h23; 
localparam bhmgs3vgnseqkofaq     = 7'h24; 
localparam v1p67sbkplioln574gw     = 7'h25; 
localparam s8hr7m7qhl3pqnt89tus     = 7'h26; 
localparam z6pqul13taj_bw4t8yli     = 7'h27; 
localparam hvhnim02z6srj83lugw     = 7'h28; 
localparam v7um53_ht6a2cwt6ubl2u5     = 7'h29; 
localparam usr_d4ztbwfqnw1ksw    = 7'h2a; 
localparam s8z4ks84p0yw2dqwwu    = 7'h2b; 
localparam fbu4pj38gfgemse5eu    = 7'h2c; 
localparam vf67ei0xuhdiywaae5mejm    = 7'h2d; 
localparam p_0cn2roe14mgc29a_0h    = 7'h2e; 
localparam oo6atcmpor7odv_pblz40y    = 7'h2f; 
localparam zym_cwfh2nuxo_oxcw6bw     = 7'h30; 
localparam klufzp92vwn000j_r     = 7'h34; 
localparam if4yqcjnanofw8tsvk     = 7'h35; 
localparam qnwyvxc9qyjqiu         = 7'h38; 
localparam co7pv8p2kbxe610a1fd6iz   = 7'h39; 
localparam jscy4q366gyq9lj13lo9r_t   = 7'h3a; 
localparam gdv3d9wl61p6agakjyorlu6   = 7'h3b; 
localparam gv3onvtfu_6pjps2fsz57vdz   = 7'h37; 
localparam jebjru_ggwvrtiwo8i      = 7'h3c; 
localparam gzcyq45ld9_ynnk5      = 7'h3d; 
localparam lm2c1fdkx8du93b_9      = 7'h3e; 
localparam g11_czp4uyqfn8ri      = 7'h3f; 
localparam mibasbdgzaznbi2ob     = 7'h40; 

localparam ab7kwrui0s1r8kz79uhlqz7r5mr4   = 8'd0;
localparam kq0d6o4iyx1q0712xrn2q2vkx = 8'd1;
localparam codaguzz0hwulmki8plk05a1tl   = 8'd2;

localparam ehf3lwj21fbudakfx9            = 3'd0;
localparam vgmgeaege4ia7hc           = 3'd1;
localparam lkdjbxd5kqnn9nb2p5y           = 3'd2;
localparam k1sebqfctqpk8z5tjg2           = 3'd3;
localparam tjmq_rg9o5kadjhk8_8j          = 3'd4;

localparam o59fpx2uri35181_3    = 32'h0c000067;
localparam l9p1t88zjkrw40pc19w    = 32'h0c000067; 
localparam zb7ej570mlfj5nga2iq9n    = 32'h0c000067; 
localparam ttjbn9c39ziunmsqvyt    = 32'h0c000067; 
localparam x43bxje5ood716p3ewb44    = 32'h0c000067; 

localparam v6a2pq_r9u9jjruu3_0   = 32'h10002823; 
localparam sbkhg6a0xgle32g3qh4p5   = 32'h10003823; 
localparam zqadrc1g014wtff      = 32'h00100073; 
localparam lw1dbr_2sxgdvqw4ag9      = 32'h00100073; 
localparam ojkmt8smt2g3rt9_r      = 32'h00100073; 
localparam b8fuv4qamrktz5      = 32'h00100073; 
localparam mphvh77x3qvz64dve6ar  = 32'h11002003; 
localparam qfki0v58jfcm7t_7a_  = 32'h11003003; 
localparam hk1d50nomn852ogmbwe     = 32'h00100073; 
localparam vc0w4jfxcmp1r_kb9     = 32'h00100073; 
localparam xyg1xr26xs6qt6mw     = 32'h00100073; 
localparam l82h342indxya4fnbl3     = 32'h00100073; 

localparam rm8dp943k0hbg_qy7gz      = 32'h7b241073; 
localparam ro0dzuoqm2k_us      = 32'h00002473; 
localparam z1z04a0vufecicvf7   = 32'h10802823; 
localparam gikah_txr49gtlzegcmj   = 32'h10803823; 
localparam f6nmwrhtc_gb4ykzjj      = 32'h7b202473; 
localparam z9jwkhk9cwds_v5ubn      = 32'h00100073; 
localparam d_ig0fq99exm8z4jy     = 32'h7b241073; 
localparam pc77kpt0abvc6o3xhgn7i  = 32'h11002403; 
localparam eniodzjwoauk00u11m  = 32'h11003403; 
localparam ak7gz0yi0kxpw8z7     = 32'h00041073; 
localparam kdz_pr5joy8wipqla_     = 32'h7b202473; 
localparam sgc8ol5jlaevuv07     = 32'h00100073; 

localparam pf3vmukxzld2et0wh_   = 32'h10002827; 
localparam bkietnnm_hbspgy2ur2sjf   = 32'h10003827;
localparam k9h3cv1wrsp7a7wpw      = 32'h00100073; 
localparam tkkhwilip2oxzggnzi      = 32'h00100073; 
localparam oc9r5_g2zdczf3p4f      = 32'h00100073; 
localparam u5ys83_oeisyxjd5e2v      = 32'h00100073; 
localparam kd7okwnxh7t20omqd410  = 32'h11002007; 
localparam r74d5l3oriykht4fyweu_hg  = 32'h11003007;
localparam x6227zjrpjm3mdfsc     = 32'h00100073; 
localparam oq0sa356rzsq90uwe     = 32'h00100073; 
localparam k3jcnoac4dv7nmf1rd     = 32'h00100073; 
localparam wr9dvag5mtzl3g_o     = 32'h00100073; 

localparam n8p49ekdadplzitwuu1             = 32'h7b241073; 
localparam mawisj0ia103jmgb54l             = 32'h7b349073; 
localparam u1o80zaq399be4zdsvr          = 32'h11402403; 
localparam xiiana7rbmfi_g5nq46cdn          = 32'h11803403;
localparam yoi2vbg6_iuvbpeeb15wz9g          = 32'h00040483; 
localparam ivqg_9qn9_lamvdwj0p          = 32'h11000483; 
localparam j5xthrnyb6jds0ekx7sf1e9u          = 32'h10900823; 
localparam cl_om0j9wxjp0pjuxnvy0rhv          = 32'h00940023; 
localparam z27u882vc07txf4814             = 32'h04c00067; 
localparam tvzm54h6oon_p38x36tt_3i55    = 32'h00040413; 
localparam tcmkcr01iujkuillkgfv418hq0dn = 32'h10802a23; 
localparam gvthnhy9isgbkedr5_xx_vhuxqi5d4n69 = 32'h10803c23;
localparam ge__d50r7pvcz6gf5nlm7bpgkq    = 32'h04c00067; 

localparam wmampknl  = 32'h00000023;    

localparam iz1a4m352icv   = 3'd2;

localparam h7qm4gdchgihbuedfbw = 7'h20;
localparam hs8t66qyp4msmj09sw2f = 7'h21;
localparam df826w0tr0ujt7no0z_0 = 7'h22;
localparam kq1q6g2z5s8vy9k299 = 7'h23;
localparam o0b3kayk7gpelof4ct = 7'h24;
localparam z33hhrxaoe7pynkmajp = 7'h25;
localparam e5e_dbyenxum0n6fkma5 = 7'h26;
localparam f9c4ft2ssszfdi08g80izc = 7'h27;
localparam gi5jphcqr7h5thk_51pyd = 7'h28;
localparam ddhlrph4_v54mbed5s = 7'h29;
localparam skp_pdoqmdedyfu_n7gaim= 7'h2a;
localparam pag68qsx0tzz0rfi62_k= 7'h2b;
localparam y7gg_6j22rearaq_a17d= 7'h2c;
localparam hqy0tjlggju7tzcwj5w= 7'h2d;
localparam min8yg2hamzo88dzhaf= 7'h2e;
localparam uffmjzklgdk28p9xvwyua8= 7'h2f;

localparam gixg8zsazjmz1x_brls  = 7'h30;
localparam ufd6dm208s7jyarlo651ta  = 7'h31;
localparam hzzi56ur3pc3ozd55y9  = 7'h32;
localparam grybk8armp6w_25n2athlf  = 7'h33;
localparam zvqpf_dzodsppyt2sy_  = 7'h34;
localparam kknbs_o3gqn0uzb6uxydb  = 7'h35;
localparam t9kao6jz00ceq9met6r  = 7'h36;
localparam bk1_dfc2yewnml9b67xq  = 7'h37;
localparam vdoigs60y4azen6d3tcs  = 7'h38;
localparam ui48c9q5f2turr4gak47g  = 7'h39;
localparam ytd01d3exnn7ehvy8m4gi = 7'h3a;
localparam ohbi7syrfghop_1ei_7_v = 7'h3b;
localparam fpg_uog8qlop0ciegpq = 7'h3c;
localparam c1lm4w95w1htl5nau42b = 7'h3d;
localparam xvf_oe_m8metbe7ln0og8m7x = 7'h3e;
localparam ougtjwdhlld141546ol2ns = 7'h3f;

localparam km0i5rel2kki7saovbnju   = 7'h40;
localparam yupij6i5uojje3u3bdgiy5= 7'h41;
localparam yhf4gk3fjs1g0c7vmxpfv  = 7'h42;
localparam mjsby4jqzutfz8ukh   = 7'h43;


localparam qj3a7cq7w0bujncuh	= 7'h44;
localparam mt_9sbagghbuv5a	= 7'h45;
localparam uqw9t32734czfnllj	= 7'h46;
localparam uvrkvxlxjv2ua24u	= 7'h47;
localparam u62d_7aeq5rs779p	= 7'h48;
localparam gn9rrcsi47vfyzz	= 7'h49;
localparam qrwi8l03c71sin9ruze	= 7'h4a;
localparam k7w_di6hk2v68wdy6_8	= 7'h4b;

localparam axd20af5hznmm5	= 32'h00100073;

localparam pn11iufvnvon1yjbw   = 3;
localparam sctcxvmp891m32rpg4w    = 3'b000;
localparam iyneurriss9qaw5wv5vz   = 3'b001;
localparam ldooojs2eemqgx70     = 3'b011;
localparam p_n8ldx18y53b6dr_6     = 3'b010;
localparam i2hy3177smkb_6w99thp  = 3'b110;












wire [smfpyk6-1:0] v91_a0d_e2l7g2npx2;
wire [smfpyk6-1:0] ua3hwncs2rj394m9h37;
wire [smfpyk6-1:0] ddm8a15ioc926sq2d;
wire [smfpyk6-1:0] a7pselnd0w05duz_ivqvp;
wire [smfpyk6-1:0] kq95iaja2o219ajkg2_jfny5v;
wire [smfpyk6-1:0] wxul7qtqbzvhly_rlbtr4lica;

wire        xgi_ovaieihs4f;

wire [31:0] r65hrblk6cfz_;     
wire [31:0] q7xpkacoiqp__elsg;    
wire [31:0] tchrn3tov0okb6f;     
wire [31:0] ws9kutgi4r0wui1;      
wire [31:0] y80_gmc7mbs2g68;      
wire [31:0] rwyvi96_wuktwcs65;      
wire [31:0] dr8lpark3fykgiqvl;      
wire [31:0] s51p9m5pter6agwkfmi;  
wire [31:0] lu2p7m5sdkbd;     
wire [31:0] stcjaa1sbc18df8;   
wire [31:0] hq9truyassja3d8s;      
wire [31:0] kg9c2fr3o4t1l2_udn; 
wire [11:0] cluaz37po70qc66wuio;
wire [15:0] xmgisya42ikqz7vaea3lpoj;

wire [2:0] iro64ooeeusz4ro;
wire [2:0] b69xflf6dvza7n0;
wire       zlzdpgdm7uynjpt_tg;

wire [31:0] roo2isb7xjjd372j766;  
wire [31:0] osmjr77x4r43r658pa;  
wire [31:0] h0s2y_7k2obvxraruu45;  
wire [31:0] rewvin436j1jc4w;  

wire [31:0] ajymk4x2v3;        
wire [31:0] mlyn8clead;        
wire [31:0] g2544euz9jpuu9;        
wire [31:0] rw_eqfvro8;        


wire [31:0] dmi_progbuf0; 
wire [31:0] i053jzqawhse;     
wire [31:0] tg3msrog_0bv;     
wire [31:0] g30pvzblnaf83zh;     
wire [31:0] j2juyav34kkmuqd;     
wire [31:0] watz9oqgogsyjeo;     
wire [31:0] kriizvysvcfvd;     
wire [31:0] l97zx3ot2wagshr9;     
wire [31:0] heiy5swkajxipcai;     
wire [31:0] etxdm_c986j2h;     
wire [31:0] iw9ukx193kjidkn;     
wire [31:0] hwwlvkrpw_rd1;     
wire [31:0] b81eb_9kn7xgu725;     
wire [31:0] rj3ujsskxnsw3;     
wire [31:0] fp511hjp_uccxk4;     
wire [31:0] dde_945nq4horxo;     



wire  [31:0] gsmp8y890cng;         
wire  [31:0] y2bt8u7bruuxsctix;   
wire  [31:0] zbawca6o200bvbpa1b6;   
wire  [31:0] bxlgqasel4nu6fjtmnt;   
wire  [31:0] e7wcd07jh85sk_hny6;   
wire  [31:0] oqevdjmfdhtvo;      
wire  [31:0] o12utn841wpwhrex;      
wire  [31:0] ayv5i_2icurn_;      
wire  [31:0] ue0zf04oji91y_44;      

wire        k53u3hfcf_oxdneqvc;
wire        prkl04ot6l0th2kjj3lensn;
wire        hoj1dk896qa8vjbobz;

wire        bf0mjxu4_jjk1oq;
wire        j3_0mc1_bfh0;

wire [31:0] hs4cmw6ypuuets98;

wire [31:0] xcgzxr3t0rc1243;
wire [31:0] f0ggwdo3sb91;
wire [31:0] cz26a1huhfl0;
wire [31:0] v7on9ph3nyz9r0;

wire [2:0]  yqdpagjrodj;
wire [2:0]  ikkfsfp;
wire [2:0]  bghtgz;
wire        wl4tlno7ko = yqdpagjrodj != sctcxvmp891m32rpg4w;
wire [9:0]  aswynak3c52xoo5;
wire [1023:0] oht8t1ux9vjcpjl842vlmyq = 1024'd1 << aswynak3c52xoo5;



wire [31:0] k42ki1zy09wlmo2;
wire [31:0] y8bs2_4f4deqi4oqg;
wire [31:0] ho5oon65ncaswgb0lj5;
wire [31:0] myuss9m1qp8gey0847r;
wire [31:0] axg6blt2b1j88hjl4_;
wire [31:0] l14fz29ful6_0ky8jl;
wire [31:0] zzsj3yl_71x_1q2lh09b;
wire [31:0] vw8sa1crlzg24r4;
wire [31:0] e0nj0rk_rp0knkls;
wire [31:0] r_tf74b2bwwlb6s1wi;
wire [31:0] xade4a80z8ri9n6tfuin4;
wire [31:0] s6ecnce9dbhjl8lyg3s7s;
wire [31:0] rfhaugdrqwldacohp91;
wire [31:0] e1ptokxdw97811mlgkh;
wire [31:0] ly2r1ofg_z2vx4ron71;
wire [31:0] zx1kehbfsf4fsgtm5;



wire          f6umtn3v33g4;
wire          i2r6o0rnjrg_t8c65;
wire    [9:0] hnvgp5pvvjoaa527;
wire [1023:0] amjh0bop7ptd8znl3hi = 1024'd1 << hnvgp5pvvjoaa527;
wire [1023:0] u5p7r7vyhmyho6aa;
wire [1023:0] duox68l_r_f8nou99k2;
wire [1023:0] n2y0qyph75pffp3dwwf80;
wire [1023:0] qfy5nt0fzqzm85nkaj;
wire          wse0ogbls179;
wire          f_bjjlctco54pp3;


wire [31:0] nd7gkqyz8zkdg3;
wire ai18gqgs_7ews5o;
wire ci1v3d4sfydbh_sz;

wire	[63:0]			qvpivcc8d7j57jlwl;
wire	[8:2]			uqi13ctmbgrce5j9;
wire	[2:0]			yygzyugpvajoy2ito;
wire	[8:2]			bf2jgqu2qq_lbyd;
wire	[63:0]			vq_q6kxvnkkqf2;




wire lypfqocyyrqu   = (yqdpagjrodj == sctcxvmp891m32rpg4w);
wire ebc4u4oafhzae  = (yqdpagjrodj == iyneurriss9qaw5wv5vz);
wire kjd3v6ed24ptvm    = (yqdpagjrodj == ldooojs2eemqgx70);
wire rknmpp444d3ijb    = (yqdpagjrodj == p_n8ldx18y53b6dr_6);
wire y4o106ig3ae61 = (yqdpagjrodj == i2hy3177smkb_6w99thp);

wire	arfgqzn8b91r3e;
wire	bfdnuw8phzaai12zaen;
wire	glencod3i3o7mjo7n25;
wire	pqyrjnamrpuq0yq9ny4;

wire	u06qbygttylwtj63blcgmn;
wire	d65omgobthbz58hr4v6c8vye;
wire	xjstumkuxktuwybrt70f09d;
wire	oq56n5j5gd3i2trf1n23;
wire	rgr3u9u7smu2_9zb3od6u4;
wire  [7:0] qxlm3tn20surby98;
wire [31:0] dk5qlcqv4hzz3221yncmzmjpc;
wire [31:0] p009emefkiuou558jih1od36;

wire  [9:0] zsnjingqe8568rcb3etc0gud;
wire        eayknskh17rtgo6n7hxacs7;
wire        qfk9f0qt00j7_h08dsa;
wire [31:0] c3b14wbbm2jilagqe = {21'd0, eayknskh17rtgo6n7hxacs7, zsnjingqe8568rcb3etc0gud} | {16'h0, arfgqzn8b91r3e, {15{~qfk9f0qt00j7_h08dsa}}};
wire [31:0] hn_zgnzhnj4hl = 32'd0;
wire [31:0] l5hh1f8jbhu6 = 32'd0;
wire [31:0] us8z6yxgvplahq18t = 32'd0;

wire        tf1byd_17w8d_ypae4v;
wire        p1yn5zqqxm8yw8ox;
wire        h3e4drj186x9hakap0e;
wire        uev0sc6o93o2rcvvy3p;
wire        lxnlpqnqclk48r5;
wire        w6r9d62ex8olvrj0zfd7;
wire        qcv2n1t0m8gvo5cto;
wire        w3f078jh09ukd9z_24;

wire [7:0]  hypvwiccin6_ahhv_    = hq9truyassja3d8s[31:24];
wire [2:0]  se0uenxs        = hq9truyassja3d8s[22:20]; 
wire        c5wsbnd7s80w3    = hq9truyassja3d8s[18];
wire        t3x39m8_1mr3    = hq9truyassja3d8s[17];
wire        hs0_yb7rhjcb       = hq9truyassja3d8s[16];
wire [15:0] r534zqz5n5zn       = hq9truyassja3d8s[15:0];
wire        o1gtiubjijenv6  = hq9truyassja3d8s[23]; 
wire [2:0]  fobztko7kz04d     = hq9truyassja3d8s[22:20];
wire        dxbb_aq_7hh19futiev = hq9truyassja3d8s[19];

wire [7:0]  he9dr9my5qt0vrui = hs4cmw6ypuuets98[31:24];
wire        o2cn09h2l79zhpeg8t7t      = (hypvwiccin6_ahhv_    == ab7kwrui0s1r8kz79uhlqz7r5mr4);
wire        iuasmef2ixpgpp9wrfgatqf    = (hypvwiccin6_ahhv_    == kq0d6o4iyx1q0712xrn2q2vkx);
wire        ook1gy0486_unhf32zio3qj7_w = (he9dr9my5qt0vrui == kq0d6o4iyx1q0712xrn2q2vkx);
wire        tbldq1rirf40guoxqqaheb      = (hypvwiccin6_ahhv_    == codaguzz0hwulmki8plk05a1tl);
wire        xl9kvstr9tbbh6vaejjlks7bkz   = o2cn09h2l79zhpeg8t7t | iuasmef2ixpgpp9wrfgatqf |
                                      (tbldq1rirf40guoxqqaheb & !o1gtiubjijenv6 & (fobztko7kz04d < tjmq_rg9o5kadjhk8_8j));
wire        i38u6n1ltlug0pip9m_;
wire        umwi6wlplo34froaxm6t = xl9kvstr9tbbh6vaejjlks7bkz & i38u6n1ltlug0pip9m_;
wire        krbd9wuik05rhl6vnfy5vh;

wire [31:0] jdv2ldkc9_q;
wire [31:0] mrse_xs0n5gn;
wire [31:0] qqgwfuykbb;
wire [31:0] tp7gcrgcgawl;
wire [31:0] atyzruk57fe;
wire [31:0] xwh383jprd;
wire [31:0] fsq3dvu1_f7r;
wire [31:0] swxb1euiqwukq;
wire [31:0] p05lkgp9i7yf5v7kf6ezjh;
wire [31:0] idw6r8r6c3kgxzbgpueg_5p;
wire [31:0] vochzpcnthf8mdr3hu6v4gd;
wire [31:0] twt3do1dqemkx_6d0fk5vtpv;
wire [31:0] trklo3qzr4u7a5f82_vg3j;
wire [31:0] fw0a5zyieal7nklrb8k_dcxx;
wire [31:0] lt3terzuwdjdjc96d_zwesq;
wire [31:0] lbjdrod2knedotqaks4ipqaa;
wire [31:0] r0ok7yh87dtunpb0fudogp4k;
wire [31:0] eltv7ctz_s7iqg4smemy0v7r0j;
wire [31:0] sp1_1j2w5w86h50jnnmw8xt;
wire [31:0] pgnid94xfwqpnd4n8a6ycd;
wire [31:0] pio7c42xp4l1mb_fskjs8uov6;

wire [31:0] aexbky0mi1u2lm2 = (se0uenxs == iz1a4m352icv) ? mphvh77x3qvz64dve6ar : qfki0v58jfcm7t_7a_; 
wire [31:0] r59f3p56s5agr3vv  = (se0uenxs == iz1a4m352icv) ? v6a2pq_r9u9jjruu3_0  : sbkhg6a0xgle32g3qh4p5;
wire [31:0] z7wp33594clq7ibe = (se0uenxs == iz1a4m352icv) ? kd7okwnxh7t20omqd410 : r74d5l3oriykht4fyweu_hg;
wire [31:0] l1u_dqv1wdbramd9a  = (se0uenxs == iz1a4m352icv) ? pf3vmukxzld2et0wh_  : bkietnnm_hbspgy2ur2sjf;

wire [2:0]  l8ptm_lp0j77nau_bwl1jt = {hs0_yb7rhjcb,r534zqz5n5zn[12],r534zqz5n5zn[5]};
assign p05lkgp9i7yf5v7kf6ezjh = (l8ptm_lp0j77nau_bwl1jt == 3'b000) ? rm8dp943k0hbg_qy7gz :
                               (l8ptm_lp0j77nau_bwl1jt == 3'b001) ? rm8dp943k0hbg_qy7gz :
                               (l8ptm_lp0j77nau_bwl1jt == 3'b010) ? (r59f3p56s5agr3vv | {7'd0, r534zqz5n5zn[4:0], 20'd0}) :
                               (l8ptm_lp0j77nau_bwl1jt == 3'b011) ? (l1u_dqv1wdbramd9a | {7'd0, r534zqz5n5zn[4:0], 20'd0}) :
                               (l8ptm_lp0j77nau_bwl1jt == 3'b100) ? d_ig0fq99exm8z4jy :
                               (l8ptm_lp0j77nau_bwl1jt == 3'b101) ? d_ig0fq99exm8z4jy :
                               (l8ptm_lp0j77nau_bwl1jt == 3'b110) ? (aexbky0mi1u2lm2 | {20'd0, r534zqz5n5zn[4:0], 7'd0}) :
                               (z7wp33594clq7ibe | {20'd0, r534zqz5n5zn[4:0], 7'd0});

















wire [31:0] x5ccz3mwtq7rnf3zf1 = (se0uenxs == iz1a4m352icv) ? pc77kpt0abvc6o3xhgn7i : eniodzjwoauk00u11m;
wire [2:0] sk6mnvnxbbqq6w0ji5j62a = {hs0_yb7rhjcb,r534zqz5n5zn[12],r534zqz5n5zn[5]};

assign idw6r8r6c3kgxzbgpueg_5p = (sk6mnvnxbbqq6w0ji5j62a == 3'b000) ? (ro0dzuoqm2k_us | {r534zqz5n5zn[11:0],20'd0}) :
                               (sk6mnvnxbbqq6w0ji5j62a == 3'b001) ? (ro0dzuoqm2k_us | {r534zqz5n5zn[11:0],20'd0}) :
                               (sk6mnvnxbbqq6w0ji5j62a == 3'b010) ? (c5wsbnd7s80w3 ? l9p1t88zjkrw40pc19w : zqadrc1g014wtff) :
                               (sk6mnvnxbbqq6w0ji5j62a == 3'b011) ? (c5wsbnd7s80w3 ? l9p1t88zjkrw40pc19w : k9h3cv1wrsp7a7wpw) :
                               (sk6mnvnxbbqq6w0ji5j62a == 3'b100) ? (x5ccz3mwtq7rnf3zf1) :
                               (sk6mnvnxbbqq6w0ji5j62a == 3'b101) ? (x5ccz3mwtq7rnf3zf1) :
                               (sk6mnvnxbbqq6w0ji5j62a == 3'b110) ? (c5wsbnd7s80w3 ? l9p1t88zjkrw40pc19w : hk1d50nomn852ogmbwe) :
                               (c5wsbnd7s80w3 ? l9p1t88zjkrw40pc19w : x6227zjrpjm3mdfsc);


















wire [31:0] zmfnwoy4sy7m9ek  = (se0uenxs == iz1a4m352icv) ? z1z04a0vufecicvf7  : gikah_txr49gtlzegcmj;
wire [2:0] qed08jt0swd30yj3tbm3pp = {hs0_yb7rhjcb,r534zqz5n5zn[12],r534zqz5n5zn[5]};

assign vochzpcnthf8mdr3hu6v4gd = (qed08jt0swd30yj3tbm3pp == 3'b000) ? zmfnwoy4sy7m9ek : 
                               (qed08jt0swd30yj3tbm3pp == 3'b001) ? zmfnwoy4sy7m9ek : 
                               (qed08jt0swd30yj3tbm3pp == 3'b010) ? lw1dbr_2sxgdvqw4ag9 : 
                               (qed08jt0swd30yj3tbm3pp == 3'b011) ? tkkhwilip2oxzggnzi : 
                               (qed08jt0swd30yj3tbm3pp == 3'b100) ? ak7gz0yi0kxpw8z7 | {r534zqz5n5zn[11:0],20'd0} :
                               (qed08jt0swd30yj3tbm3pp == 3'b101) ? ak7gz0yi0kxpw8z7 | {r534zqz5n5zn[11:0],20'd0} : 
                               (qed08jt0swd30yj3tbm3pp == 3'b110) ? vc0w4jfxcmp1r_kb9 : 
                               (oq0sa356rzsq90uwe);

















wire [2:0] pj2atqm338pqv_diim85 = {hs0_yb7rhjcb,r534zqz5n5zn[12],r534zqz5n5zn[5]};

assign twt3do1dqemkx_6d0fk5vtpv = (pj2atqm338pqv_diim85 == 3'b000) ? f6nmwrhtc_gb4ykzjj : 
                               (pj2atqm338pqv_diim85 == 3'b001) ? f6nmwrhtc_gb4ykzjj : 
                               (pj2atqm338pqv_diim85 == 3'b010) ? ojkmt8smt2g3rt9_r : 
                               (pj2atqm338pqv_diim85 == 3'b011) ? oc9r5_g2zdczf3p4f : 
                               (pj2atqm338pqv_diim85 == 3'b100) ? kdz_pr5joy8wipqla_ : 
                               (pj2atqm338pqv_diim85 == 3'b101) ? kdz_pr5joy8wipqla_ : 
                               (pj2atqm338pqv_diim85 == 3'b110) ? xyg1xr26xs6qt6mw :
                               (k3jcnoac4dv7nmf1rd);

















wire [2:0] d6t8jbw4yj18hw7azral = {hs0_yb7rhjcb,r534zqz5n5zn[12],r534zqz5n5zn[5]};

assign trklo3qzr4u7a5f82_vg3j = (d6t8jbw4yj18hw7azral == 3'b000) ? (c5wsbnd7s80w3 ? x43bxje5ood716p3ewb44 : z9jwkhk9cwds_v5ubn) : 
                               (d6t8jbw4yj18hw7azral == 3'b001) ? (c5wsbnd7s80w3 ? x43bxje5ood716p3ewb44 : z9jwkhk9cwds_v5ubn) : 
                               (d6t8jbw4yj18hw7azral == 3'b010) ? (b8fuv4qamrktz5) : 
                               (d6t8jbw4yj18hw7azral == 3'b011) ? (u5ys83_oeisyxjd5e2v) : 
                               (d6t8jbw4yj18hw7azral == 3'b100) ? (c5wsbnd7s80w3 ? x43bxje5ood716p3ewb44 : sgc8ol5jlaevuv07) : 
                               (d6t8jbw4yj18hw7azral == 3'b101) ? (c5wsbnd7s80w3 ? x43bxje5ood716p3ewb44 : sgc8ol5jlaevuv07) : 
                               (d6t8jbw4yj18hw7azral == 3'b110) ? (l82h342indxya4fnbl3) :
                               (wr9dvag5mtzl3g_o);

















assign fw0a5zyieal7nklrb8k_dcxx = n8p49ekdadplzitwuu1;
assign lt3terzuwdjdjc96d_zwesq = mawisj0ia103jmgb54l;

assign lbjdrod2knedotqaks4ipqaa = xiiana7rbmfi_g5nq46cdn;
assign r0ok7yh87dtunpb0fudogp4k = (hs0_yb7rhjcb)? ivqg_9qn9_lamvdwj0p | {17'd0, fobztko7kz04d, 12'd0} :
                                            yoi2vbg6_iuvbpeeb15wz9g | {17'd0, fobztko7kz04d, 12'd0} ;
assign eltv7ctz_s7iqg4smemy0v7r0j = (hs0_yb7rhjcb)? cl_om0j9wxjp0pjuxnvy0rhv | {17'd0, fobztko7kz04d, 12'd0} :
                                            j5xthrnyb6jds0ekx7sf1e9u | {17'd0, fobztko7kz04d, 12'd0} ;  
assign sp1_1j2w5w86h50jnnmw8xt = (dxbb_aq_7hh19futiev)? (tvzm54h6oon_p38x36tt_3i55 | (32'h100000 << fobztko7kz04d)) : z27u882vc07txf4814;
assign pgnid94xfwqpnd4n8a6ycd = (fobztko7kz04d ==  k1sebqfctqpk8z5tjg2)? gvthnhy9isgbkedr5_xx_vhuxqi5d4n69 : tcmkcr01iujkuillkgfv418hq0dn;
assign pio7c42xp4l1mb_fskjs8uov6 = ge__d50r7pvcz6gf5nlm7bpgkq;

assign jdv2ldkc9_q = tbldq1rirf40guoxqqaheb ? fw0a5zyieal7nklrb8k_dcxx :
                   o2cn09h2l79zhpeg8t7t ? (t3x39m8_1mr3 ? p05lkgp9i7yf5v7kf6ezjh : 
	                                (c5wsbnd7s80w3 ? o59fpx2uri35181_3 : axd20af5hznmm5)) :
		                        o59fpx2uri35181_3;
assign mrse_xs0n5gn = tbldq1rirf40guoxqqaheb ? lt3terzuwdjdjc96d_zwesq : idw6r8r6c3kgxzbgpueg_5p;
assign qqgwfuykbb = tbldq1rirf40guoxqqaheb ? lbjdrod2knedotqaks4ipqaa : vochzpcnthf8mdr3hu6v4gd;
assign tp7gcrgcgawl = tbldq1rirf40guoxqqaheb ? r0ok7yh87dtunpb0fudogp4k : twt3do1dqemkx_6d0fk5vtpv;
assign atyzruk57fe = tbldq1rirf40guoxqqaheb ? eltv7ctz_s7iqg4smemy0v7r0j : trklo3qzr4u7a5f82_vg3j;
assign xwh383jprd = tbldq1rirf40guoxqqaheb ? sp1_1j2w5w86h50jnnmw8xt : axd20af5hznmm5;
assign fsq3dvu1_f7r = tbldq1rirf40guoxqqaheb ? pgnid94xfwqpnd4n8a6ycd : axd20af5hznmm5;
assign swxb1euiqwukq = tbldq1rirf40guoxqqaheb ? pio7c42xp4l1mb_fskjs8uov6 : axd20af5hznmm5;

localparam p0t159zwkkyyulx = 2'b00;
localparam kapv0q86iup = 2'b01;
localparam g9rl8dm8yn = 2'b00;
assign xgi_ovaieihs4f = jutj9q2kpi & hy7ogyog4pk_4i[1] & nrxv3rneu2438;

wire ysbkkifl78x_74yihmmou_m = nrxv3rneu2438;
wire puuni4ssasd4hxb9e5wwye  = xgi_ovaieihs4f;
wire b5xt1a6vsi17t78i;

ux607_gnrl_dfflr #(1)    p0usxt4w9fjp6w3u3kob6r1864(ysbkkifl78x_74yihmmou_m, puuni4ssasd4hxb9e5wwye, b5xt1a6vsi17t78i, gf33atgy, hfocw7va5_);
  
wire dq9zivc29hucjvuprdn8r4 = nrxv3rneu2438;
wire h8jw2c5eb33jzodbvcr  = e_pz9vwnoa1r523;
wire jvottutw7zyalqe;

ux607_gnrl_dfflr #(1)    uovpoacn0sok4bfth5b(dq9zivc29hucjvuprdn8r4, h8jw2c5eb33jzodbvcr, jvottutw7zyalqe, gf33atgy, hfocw7va5_);

wire nbekcn12qcmiu1khw1p = nrxv3rneu2438;
wire [8:2] nkbk7uazihufpo9bg  = ehdeq25ha[8:2];
wire [8:2] cohyjbtg_qyh;

ux607_gnrl_dfflr #(7)    rk4vlae8x3rs28s9kthp1(nbekcn12qcmiu1khw1p, nkbk7uazihufpo9bg, cohyjbtg_qyh, gf33atgy, hfocw7va5_);











wire eui3agxj55ryll499;

wire qv2gqnqu4n7y26eo1sz0quji = (hy7ogyog4pk_4i[1]==1'b0);
wire nefljqb0lyofqktzke6vjt8woprdggdmz8 = jvottutw7zyalqe & b5xt1a6vsi17t78i & !e_pz9vwnoa1r523;
assign eui3agxj55ryll499 = qv2gqnqu4n7y26eo1sz0quji | !nefljqb0lyofqktzke6vjt8woprdggdmz8;

wire c11wmha0o0y3y_r2hw = 1'b1;
wire h1b8r20c_rynl_bg3udlvr = eui3agxj55ryll499;

ux607_gnrl_dfflrs #(1)    x39eptcbrfepf_pg5973xwj(c11wmha0o0y3y_r2hw, h1b8r20c_rynl_bg3udlvr, f2r3r2mwmdler, gf33atgy, hfocw7va5_);










assign o4hlkc18armddz = g9rl8dm8yn;

assign roo2isb7xjjd372j766 = 32'd0;
assign osmjr77x4r43r658pa = 32'd0;
assign h0s2y_7k2obvxraruu45 = 32'd0;
assign rewvin436j1jc4w = 32'd0;












assign k53u3hfcf_oxdneqvc    = b5xt1a6vsi17t78i & jvottutw7zyalqe & (cohyjbtg_qyh == wjwm0mmb8kdtc38hmvxcg7);
assign hoj1dk896qa8vjbobz     = b5xt1a6vsi17t78i & jvottutw7zyalqe & (cohyjbtg_qyh == jcqkgadqjnp1br60kcm7);

wire   s6m193phbzzswom34s   = b5xt1a6vsi17t78i & jvottutw7zyalqe & (cohyjbtg_qyh == xpf4_70tcyabeblxkt7aob2y);
wire   bxgr20exryirwahrpndyb8w14mai   = ~wl4tlno7ko & s6m193phbzzswom34s;
wire   src1s9kkdw9sn9kvu6z4      = b5xt1a6vsi17t78i & jvottutw7zyalqe & (cohyjbtg_qyh == bcei3m4eneqv0kswce_6);
wire   ohlejrcx6cdwmphlr      = b5xt1a6vsi17t78i & ((cohyjbtg_qyh == ggr6ql2zj7x40114w) |
                                                  (cohyjbtg_qyh == tcnwfsqopcq2kj) |
						  (cohyjbtg_qyh == ab_j1frhbffg57rc) |
						  (cohyjbtg_qyh == jim0ddiqnav_mr) |
						  (cohyjbtg_qyh == m0jpn5dn80dsf2q) |
						  (cohyjbtg_qyh == zxe9_q2s5fzxgu_k38) |
						  (cohyjbtg_qyh == va10rh7n02nkb6) |
						  (cohyjbtg_qyh == dmgo2idd7_vdsdnnaq3) |
						  (cohyjbtg_qyh == jbtj7er6n1t919tqlx) |
						  (cohyjbtg_qyh == qz57tyn0hruiw2xcq) |
						  (cohyjbtg_qyh == kfpiwe2xk_8vve0)|
						  (cohyjbtg_qyh == esrb21vaoahytvbimz));

wire   k9ddbzzry2og0lep5n5t6dc37_; 
wire   xl9_scab2526apfj3i0f8vd6 = b5xt1a6vsi17t78i & jvottutw7zyalqe & (cohyjbtg_qyh == rzuyw47p7ehj1uy43z4w9l63d3);
wire   utec8wet9b5ke5gtbnr__oo1hi7395v = ~wl4tlno7ko & xl9_scab2526apfj3i0f8vd6;

wire   heq7laaei2amn9igl2        = ~wl4tlno7ko & b5xt1a6vsi17t78i & jvottutw7zyalqe & (cohyjbtg_qyh == ggr6ql2zj7x40114w) | tf1byd_17w8d_ypae4v;
wire   ldbdzv1slpkxnh        = ~wl4tlno7ko & b5xt1a6vsi17t78i & jvottutw7zyalqe & (cohyjbtg_qyh == tcnwfsqopcq2kj) | p1yn5zqqxm8yw8ox;
wire   r7195x8bumqznsl        = ~wl4tlno7ko & b5xt1a6vsi17t78i & jvottutw7zyalqe & (cohyjbtg_qyh == ab_j1frhbffg57rc) | h3e4drj186x9hakap0e;
wire   wputl8m_xeys6yd2_        = ~wl4tlno7ko & b5xt1a6vsi17t78i & jvottutw7zyalqe & (cohyjbtg_qyh == jim0ddiqnav_mr) | uev0sc6o93o2rcvvy3p;

wire   hrxvvr_jkklnx6btx7 = b5xt1a6vsi17t78i &
	(
		((d8panmbslrc4xeco > 0 ) &  (cohyjbtg_qyh == ggr6ql2zj7x40114w    ) & cluaz37po70qc66wuio[0]    ) |
		((d8panmbslrc4xeco > 1 ) &  (cohyjbtg_qyh == tcnwfsqopcq2kj    ) & cluaz37po70qc66wuio[1]    ) |
		((d8panmbslrc4xeco > 2 ) &  (cohyjbtg_qyh == ab_j1frhbffg57rc    ) & cluaz37po70qc66wuio[2]    ) |
		((d8panmbslrc4xeco > 3 ) &  (cohyjbtg_qyh == jim0ddiqnav_mr    ) & cluaz37po70qc66wuio[3]    ) |
		((yv13_lx8u9yhr8p6i > 0 ) & (cohyjbtg_qyh == u_cztegv7294f0w2ck ) & xmgisya42ikqz7vaea3lpoj[0] ) |
		((yv13_lx8u9yhr8p6i > 1 ) & (cohyjbtg_qyh == ew_k_8affyv8ltn2n9t ) & xmgisya42ikqz7vaea3lpoj[1] ) |
		((yv13_lx8u9yhr8p6i > 2 ) & (cohyjbtg_qyh == c2pgc56ortybp6qk31tah2 ) & xmgisya42ikqz7vaea3lpoj[2] ) |
		((yv13_lx8u9yhr8p6i > 3 ) & (cohyjbtg_qyh == vojasz8wlqnrlmd7irtxe ) & xmgisya42ikqz7vaea3lpoj[3] ) |
		((yv13_lx8u9yhr8p6i > 4 ) & (cohyjbtg_qyh == bhmgs3vgnseqkofaq ) & xmgisya42ikqz7vaea3lpoj[4] ) |
		((yv13_lx8u9yhr8p6i > 5 ) & (cohyjbtg_qyh == v1p67sbkplioln574gw ) & xmgisya42ikqz7vaea3lpoj[5] ) |
		((yv13_lx8u9yhr8p6i > 6 ) & (cohyjbtg_qyh == s8hr7m7qhl3pqnt89tus ) & xmgisya42ikqz7vaea3lpoj[6] ) |
		((yv13_lx8u9yhr8p6i > 7 ) & (cohyjbtg_qyh == z6pqul13taj_bw4t8yli ) & xmgisya42ikqz7vaea3lpoj[7] ) |
		((yv13_lx8u9yhr8p6i > 8 ) & (cohyjbtg_qyh == hvhnim02z6srj83lugw ) & xmgisya42ikqz7vaea3lpoj[8] ) |
		((yv13_lx8u9yhr8p6i > 9 ) & (cohyjbtg_qyh == v7um53_ht6a2cwt6ubl2u5 ) & xmgisya42ikqz7vaea3lpoj[9] ) |
		((yv13_lx8u9yhr8p6i > 10) & (cohyjbtg_qyh == usr_d4ztbwfqnw1ksw) & xmgisya42ikqz7vaea3lpoj[10]) |
		((yv13_lx8u9yhr8p6i > 11) & (cohyjbtg_qyh == s8z4ks84p0yw2dqwwu) & xmgisya42ikqz7vaea3lpoj[11]) |
		((yv13_lx8u9yhr8p6i > 12) & (cohyjbtg_qyh == fbu4pj38gfgemse5eu) & xmgisya42ikqz7vaea3lpoj[12]) |
		((yv13_lx8u9yhr8p6i > 13) & (cohyjbtg_qyh == vf67ei0xuhdiywaae5mejm) & xmgisya42ikqz7vaea3lpoj[13]) |
		((yv13_lx8u9yhr8p6i > 14) & (cohyjbtg_qyh == p_0cn2roe14mgc29a_0h) & xmgisya42ikqz7vaea3lpoj[14]) |
		((yv13_lx8u9yhr8p6i > 15) & (cohyjbtg_qyh == oo6atcmpor7odv_pblz40y) & xmgisya42ikqz7vaea3lpoj[15]) 
	) 
	& !wl4tlno7ko & (iro64ooeeusz4ro == 3'd0);


wire   y6iognrzzx70lo41     = ~wl4tlno7ko & b5xt1a6vsi17t78i & jvottutw7zyalqe & (cohyjbtg_qyh == u_cztegv7294f0w2ck);
wire   ycy9ybsio5u2sv_u     = ~wl4tlno7ko & b5xt1a6vsi17t78i & jvottutw7zyalqe & (cohyjbtg_qyh == ew_k_8affyv8ltn2n9t);
wire   r7cb6vtpb7f_9k0ptq4vt     = ~wl4tlno7ko & b5xt1a6vsi17t78i & jvottutw7zyalqe & (cohyjbtg_qyh == c2pgc56ortybp6qk31tah2);
wire   b1kr1ktqldmq7upcm3     = ~wl4tlno7ko & b5xt1a6vsi17t78i & jvottutw7zyalqe & (cohyjbtg_qyh == vojasz8wlqnrlmd7irtxe);
wire   kjohxrar_xfy5le716     = ~wl4tlno7ko & b5xt1a6vsi17t78i & jvottutw7zyalqe & (cohyjbtg_qyh == bhmgs3vgnseqkofaq);
wire   wahk2cmvu9oez0oyj8pnb     = ~wl4tlno7ko & b5xt1a6vsi17t78i & jvottutw7zyalqe & (cohyjbtg_qyh == v1p67sbkplioln574gw);
wire   sque8cegtpz7u4p_     = ~wl4tlno7ko & b5xt1a6vsi17t78i & jvottutw7zyalqe & (cohyjbtg_qyh == s8hr7m7qhl3pqnt89tus);
wire   efr5v0_6lmocr1v3s     = ~wl4tlno7ko & b5xt1a6vsi17t78i & jvottutw7zyalqe & (cohyjbtg_qyh == z6pqul13taj_bw4t8yli);
wire   ov9xy25sj0yngtmtlrp     = ~wl4tlno7ko & b5xt1a6vsi17t78i & jvottutw7zyalqe & (cohyjbtg_qyh == hvhnim02z6srj83lugw);
wire   g83t3072np0dxqlin     = ~wl4tlno7ko & b5xt1a6vsi17t78i & jvottutw7zyalqe & (cohyjbtg_qyh == v7um53_ht6a2cwt6ubl2u5);
wire   ycnyqhwxogfwpkhhmqfqp     = ~wl4tlno7ko & b5xt1a6vsi17t78i & jvottutw7zyalqe & (cohyjbtg_qyh == usr_d4ztbwfqnw1ksw);
wire   k7hc4wdxsdztmi0wby5ut     = ~wl4tlno7ko & b5xt1a6vsi17t78i & jvottutw7zyalqe & (cohyjbtg_qyh == s8z4ks84p0yw2dqwwu);
wire   vo0qs9ay_75sue1lt     = ~wl4tlno7ko & b5xt1a6vsi17t78i & jvottutw7zyalqe & (cohyjbtg_qyh == fbu4pj38gfgemse5eu);
wire   s24gshk_q37q79nz9qukuv     = ~wl4tlno7ko & b5xt1a6vsi17t78i & jvottutw7zyalqe & (cohyjbtg_qyh == vf67ei0xuhdiywaae5mejm);
wire   wkpckbb4zbinpn7mx0cdo     = ~wl4tlno7ko & b5xt1a6vsi17t78i & jvottutw7zyalqe & (cohyjbtg_qyh == p_0cn2roe14mgc29a_0h);
wire   xy8ch1odd_pqev5h59zx6     = ~wl4tlno7ko & b5xt1a6vsi17t78i & jvottutw7zyalqe & (cohyjbtg_qyh == oo6atcmpor7odv_pblz40y);

wire   pf4xyp48dd4kkmpy5ab    = b5xt1a6vsi17t78i & ( (cohyjbtg_qyh == u_cztegv7294f0w2ck)
                                                  | (cohyjbtg_qyh == ew_k_8affyv8ltn2n9t)
                                                  | (cohyjbtg_qyh == c2pgc56ortybp6qk31tah2)
                                                  | (cohyjbtg_qyh == vojasz8wlqnrlmd7irtxe)
                                                  | (cohyjbtg_qyh == bhmgs3vgnseqkofaq)
                                                  | (cohyjbtg_qyh == v1p67sbkplioln574gw)
                                                  | (cohyjbtg_qyh == s8hr7m7qhl3pqnt89tus)
                                                  | (cohyjbtg_qyh == z6pqul13taj_bw4t8yli)
                                                  | (cohyjbtg_qyh == hvhnim02z6srj83lugw)
                                                  | (cohyjbtg_qyh == v7um53_ht6a2cwt6ubl2u5)
                                                  | (cohyjbtg_qyh == usr_d4ztbwfqnw1ksw)
                                                  | (cohyjbtg_qyh == s8z4ks84p0yw2dqwwu)
                                                  | (cohyjbtg_qyh == fbu4pj38gfgemse5eu)
                                                  | (cohyjbtg_qyh == vf67ei0xuhdiywaae5mejm)
                                                  | (cohyjbtg_qyh == p_0cn2roe14mgc29a_0h)
                                                  | (cohyjbtg_qyh == oo6atcmpor7odv_pblz40y)
                                                  );

wire   jqecsbcna9xks4236v7y;
wire   bg6j3mh0cbpsnjsw8;
wire   g3ss6oez6hga6h4sc;
wire   bpf8y70t6yfklo_g8w2vz;
wire   wmao806lq98cxpivg;
wire   d65wnf88ntcgv6j5aqzdd;
wire   zyrzsibwzfi9i9wbbf;
wire   lu303j9kh0__1tuhdc3wn1;
wire   meq51ng31supqk_vkxuh;
wire   vhake2p_2q859v6b79w9bt;
wire   nimnckhhiicxl3my3yxx;
wire   yi1sq51qvk1rehte9p8_;
wire   lapvh12sh70dkfu0lnktk5;
wire   ts8jeswko5lfbpmtqe;
wire   yjole_26w_x6maqonk;
wire   oj1yq4vf080z10xcce;

wire   pize1u2oxu5xj00 = y6iognrzzx70lo41 | jqecsbcna9xks4236v7y;
wire   oap_3j1l7iu77qz = ycy9ybsio5u2sv_u | bg6j3mh0cbpsnjsw8;
wire   a1lc422n48q68c7 = r7cb6vtpb7f_9k0ptq4vt | g3ss6oez6hga6h4sc;
wire   yrsrzj9xgtahq9zah = b1kr1ktqldmq7upcm3 | bpf8y70t6yfklo_g8w2vz;
wire   a3ahayu4bahs = kjohxrar_xfy5le716 | wmao806lq98cxpivg;
wire   jowfj_v52hdqypc = wahk2cmvu9oez0oyj8pnb | d65wnf88ntcgv6j5aqzdd;
wire   zhrzwed1qf5xclzq0 = sque8cegtpz7u4p_ | zyrzsibwzfi9i9wbbf;
wire   e8i6of8n537o = efr5v0_6lmocr1v3s | lu303j9kh0__1tuhdc3wn1;
wire   h5cykrla39c8zlmr = ov9xy25sj0yngtmtlrp | meq51ng31supqk_vkxuh;
wire   iwmac56d70_7 = g83t3072np0dxqlin | vhake2p_2q859v6b79w9bt;
wire   fbcol2fiz4_dakl6 = ycnyqhwxogfwpkhhmqfqp | nimnckhhiicxl3my3yxx;
wire   okw64jbuomhjb3l9he = k7hc4wdxsdztmi0wby5ut | yi1sq51qvk1rehte9p8_;
wire   xdx6hvlnkbknoa_m = vo0qs9ay_75sue1lt | lapvh12sh70dkfu0lnktk5;
wire   dzcjaphosa9ch = s24gshk_q37q79nz9qukuv | ts8jeswko5lfbpmtqe;
wire   dxhr63c235702bgyoa = wkpckbb4zbinpn7mx0cdo | yjole_26w_x6maqonk;
wire   kt7so0oerx68ydrpz = xy8ch1odd_pqev5h59zx6 | oj1yq4vf080z10xcce;


wire   ip8r6j4zqf0c24uw3v_j5     = b5xt1a6vsi17t78i & jvottutw7zyalqe & (cohyjbtg_qyh == zym_cwfh2nuxo_oxcw6bw);

wire   ka6mrfj_02knc55k6         = b5xt1a6vsi17t78i & jvottutw7zyalqe & (cohyjbtg_qyh == qnwyvxc9qyjqiu);
wire   od6u7rr1fxvo091a298   = b5xt1a6vsi17t78i & jvottutw7zyalqe & (cohyjbtg_qyh == co7pv8p2kbxe610a1fd6iz);
wire   fp20b2_fx9jb40co6__3   = b5xt1a6vsi17t78i & jvottutw7zyalqe & (cohyjbtg_qyh == jscy4q366gyq9lj13lo9r_t);
wire   iy011s14bjaestsjehfc   = b5xt1a6vsi17t78i & jvottutw7zyalqe & (cohyjbtg_qyh == gdv3d9wl61p6agakjyorlu6);
wire   m9xf9uxglv4neo5ivk3   = b5xt1a6vsi17t78i & jvottutw7zyalqe & (cohyjbtg_qyh == gv3onvtfu_6pjps2fsz57vdz);
wire   gvbp1k6dl4r0o3hg6n      = b5xt1a6vsi17t78i & jvottutw7zyalqe & (cohyjbtg_qyh == jebjru_ggwvrtiwo8i);
wire   kits5q7f_cnh6v1l      = b5xt1a6vsi17t78i & jvottutw7zyalqe & (cohyjbtg_qyh == gzcyq45ld9_ynnk5);
wire   vzl0_w7ht4urni897h3      = b5xt1a6vsi17t78i & jvottutw7zyalqe & (cohyjbtg_qyh == lm2c1fdkx8du93b_9);
wire   ppt849kffgp8e6pv9j      = b5xt1a6vsi17t78i & jvottutw7zyalqe & (cohyjbtg_qyh == g11_czp4uyqfn8ri);
wire   j0d0ajxf_i5ihg3yt95      = xgi_ovaieihs4f    & ~e_pz9vwnoa1r523   & (ehdeq25ha[8:2] == jebjru_ggwvrtiwo8i);

assign bf0mjxu4_jjk1oq      = k53u3hfcf_oxdneqvc & ph7jz_7_o_welqv[28] & ph7jz_7_o_welqv[0];


assign hs4cmw6ypuuets98      = ph7jz_7_o_welqv;

assign xcgzxr3t0rc1243        = tf1byd_17w8d_ypae4v ? (qvpivcc8d7j57jlwl[31:0] & dk5qlcqv4hzz3221yncmzmjpc) : ph7jz_7_o_welqv;
assign f0ggwdo3sb91        = p1yn5zqqxm8yw8ox ? (oq56n5j5gd3i2trf1n23 ? (qvpivcc8d7j57jlwl[vmw6vavuv7md5-1:vmw6vavuv7md5-32] & p009emefkiuou558jih1od36): (qvpivcc8d7j57jlwl[31:0] & dk5qlcqv4hzz3221yncmzmjpc)) : ph7jz_7_o_welqv;
assign cz26a1huhfl0        = h3e4drj186x9hakap0e ? (qvpivcc8d7j57jlwl[31:0] & dk5qlcqv4hzz3221yncmzmjpc) : ph7jz_7_o_welqv;
assign v7on9ph3nyz9r0        = uev0sc6o93o2rcvvy3p ? (oq56n5j5gd3i2trf1n23 ? (qvpivcc8d7j57jlwl[vmw6vavuv7md5-1:vmw6vavuv7md5-32] & p009emefkiuou558jih1od36): (qvpivcc8d7j57jlwl[31:0] & dk5qlcqv4hzz3221yncmzmjpc)) : ph7jz_7_o_welqv;


assign k42ki1zy09wlmo2     = jqecsbcna9xks4236v7y ? qvpivcc8d7j57jlwl[31:0] : ph7jz_7_o_welqv;
assign y8bs2_4f4deqi4oqg     = bg6j3mh0cbpsnjsw8 ? (oq56n5j5gd3i2trf1n23 ? qvpivcc8d7j57jlwl[vmw6vavuv7md5-1:vmw6vavuv7md5-32] : qvpivcc8d7j57jlwl[31:0]) : ph7jz_7_o_welqv;
assign ho5oon65ncaswgb0lj5     = g3ss6oez6hga6h4sc ? qvpivcc8d7j57jlwl[31:0] : ph7jz_7_o_welqv;
assign myuss9m1qp8gey0847r     = bpf8y70t6yfklo_g8w2vz ? (oq56n5j5gd3i2trf1n23 ? qvpivcc8d7j57jlwl[vmw6vavuv7md5-1:vmw6vavuv7md5-32] : qvpivcc8d7j57jlwl[31:0]) : ph7jz_7_o_welqv;
assign axg6blt2b1j88hjl4_     = wmao806lq98cxpivg ? qvpivcc8d7j57jlwl[31:0] : ph7jz_7_o_welqv;
assign l14fz29ful6_0ky8jl     = d65wnf88ntcgv6j5aqzdd ? (oq56n5j5gd3i2trf1n23 ? qvpivcc8d7j57jlwl[vmw6vavuv7md5-1:vmw6vavuv7md5-32] : qvpivcc8d7j57jlwl[31:0]) : ph7jz_7_o_welqv;
assign zzsj3yl_71x_1q2lh09b     = zyrzsibwzfi9i9wbbf ? qvpivcc8d7j57jlwl[31:0] : ph7jz_7_o_welqv;
assign vw8sa1crlzg24r4     = lu303j9kh0__1tuhdc3wn1 ? (oq56n5j5gd3i2trf1n23 ? qvpivcc8d7j57jlwl[vmw6vavuv7md5-1:vmw6vavuv7md5-32] : qvpivcc8d7j57jlwl[31:0]) : ph7jz_7_o_welqv;

assign e0nj0rk_rp0knkls     = meq51ng31supqk_vkxuh ? qvpivcc8d7j57jlwl[31:0] : ph7jz_7_o_welqv;
assign r_tf74b2bwwlb6s1wi     = vhake2p_2q859v6b79w9bt ? (oq56n5j5gd3i2trf1n23 ? qvpivcc8d7j57jlwl[vmw6vavuv7md5-1:vmw6vavuv7md5-32] : qvpivcc8d7j57jlwl[31:0]) : ph7jz_7_o_welqv;
assign xade4a80z8ri9n6tfuin4     = nimnckhhiicxl3my3yxx ? qvpivcc8d7j57jlwl[31:0] : ph7jz_7_o_welqv;
assign s6ecnce9dbhjl8lyg3s7s     = yi1sq51qvk1rehte9p8_ ? (oq56n5j5gd3i2trf1n23 ? qvpivcc8d7j57jlwl[vmw6vavuv7md5-1:vmw6vavuv7md5-32] : qvpivcc8d7j57jlwl[31:0]) : ph7jz_7_o_welqv;
assign rfhaugdrqwldacohp91     = lapvh12sh70dkfu0lnktk5 ? qvpivcc8d7j57jlwl[31:0] : ph7jz_7_o_welqv;
assign e1ptokxdw97811mlgkh     = ts8jeswko5lfbpmtqe ? (oq56n5j5gd3i2trf1n23 ? qvpivcc8d7j57jlwl[vmw6vavuv7md5-1:vmw6vavuv7md5-32] : qvpivcc8d7j57jlwl[31:0]) : ph7jz_7_o_welqv;
assign ly2r1ofg_z2vx4ron71     = yjole_26w_x6maqonk ? qvpivcc8d7j57jlwl[31:0] : ph7jz_7_o_welqv;
assign zx1kehbfsf4fsgtm5     = oj1yq4vf080z10xcce ? (oq56n5j5gd3i2trf1n23 ? qvpivcc8d7j57jlwl[vmw6vavuv7md5-1:vmw6vavuv7md5-32] : qvpivcc8d7j57jlwl[31:0]) : ph7jz_7_o_welqv;



localparam ooxsa7fkpkg7s0no142 = 4'd2;

wire       ywxqdtlc1lq30jgk8mu9;
wire       dj_0z4kpnkm667my96de;
wire       dc05a4etne0pkj7u9_nb;
wire       pqteh7_cyvhhbcf4;
wire       e6_o9xin1wu8kylws9m;
wire       gj_o1f7vjh3bs5_rkd65mtg;
wire       l8d6kinl1s6rh6ha;
wire       k68x_2_wxidbic0ld_;
wire       s942sghng1f2y8;
wire       svgpgd1koc7jztn7h2;
wire       pd9da145nlzxwlaua8;
wire       cp0_pk_fscb9h1z;
wire       zy51q_pbb9tfrc_of = 1'b1;
wire       qmur7eb6mi4y = 1'b0;
wire       a5ee5u9gnomn5itad6c8 = 1'b1;
wire       dd2_ly9t687r6v_wa = 1'b0;
wire [3:0] czyq3s7omblo1 = ooxsa7fkpkg7s0no142;

wire	   [smfpyk6-1:0] u9eb3j3kbeih0qsei71;
wire	   [smfpyk6-1:0] byyagfto1uztznf7eh;
wire	   [smfpyk6-1:0] i_1o22g1okmq7xskth;
wire	   [smfpyk6-1:0] hod7aki51hhxhaobdn;


wire       [smfpyk6-1:0] okvgcb6z3u4;
wire	   [smfpyk6-1:0] uxfmt_p8696p685;
wire	   [smfpyk6-1:0] xcl486gg7mcx74msnzz;
wire	               h90anyh0t2067aaxikbb;

wire	   [smfpyk6-1:0] c_d83vejsnlgx1b750;
wire	   [smfpyk6-1:0] g9_nradsie9gn_rr4o;
wire	               wv03_r28177pyhq87q_eku;

wire	   [smfpyk6-1:0] df7442xh1y14cj3o6qx;
wire	   [smfpyk6-1:0] je9cia8z8gc_arzaynhtmf;
wire	   [smfpyk6-1:0] r2vx5irgc6jszc2q1zg9;
wire	   [smfpyk6-1:0] tekott495862wlgwpec4r;

wire       [smfpyk6-1:0] k_g1vkidq8p8y6ghnxc4;


wire                   km788k575stdqjlb_qqfypq;
wire             [9:0] sv2fooskb173c3b58;
wire             [9:0] rir_sifntdbcly7vezk338qsh3 = sv2fooskb173c3b58 + 10'd1;
wire             [9:0] tgw362y_u7jxvpdu2t3c;
wire                   v5ciuvu6m6lmww03;

ux607_gnrl_dffr #(smfpyk6) furx7g3xqed0ewcynrhyurt8zqaj (u_ll4hq1b12s2i1       , v91_a0d_e2l7g2npx2, gf33atgy, hfocw7va5_);
ux607_gnrl_dffr #(smfpyk6) gvlkbzd8kjv7032zvdsg2k9pcu (v91_a0d_e2l7g2npx2 , ua3hwncs2rj394m9h37, gf33atgy, hfocw7va5_);

ux607_gnrl_dffr #(smfpyk6) fepf5oe26unwf5xb1kwbijn1zo_a (w41ourymsjpvm8q1e       , kq95iaja2o219ajkg2_jfny5v, dk2xhkj77a, hfocw7va5_);
ux607_gnrl_dffr #(smfpyk6) rjs4b9__csxvkgkiisif7ibq81a (kq95iaja2o219ajkg2_jfny5v , wxul7qtqbzvhly_rlbtr4lica, dk2xhkj77a, hfocw7va5_);

ux607_gnrl_dffr #(smfpyk6) n1aujcpj84c4v92ciz_ut9 (z5w8jrogg064jr       , ddm8a15ioc926sq2d, gf33atgy, hfocw7va5_);
ux607_gnrl_dffr #(smfpyk6) c13909eu7n5_uq41f4q6h69 (ddm8a15ioc926sq2d , a7pselnd0w05duz_ivqvp, gf33atgy, hfocw7va5_);

ux607_gnrl_dffr #(smfpyk6) k7wdbwroa2yfv26olf8b (byyagfto1uztznf7eh , u9eb3j3kbeih0qsei71, dk2xhkj77a, hfocw7va5_);











































assign u5p7r7vyhmyho6aa[smfpyk6-1:0]  = a7pselnd0w05duz_ivqvp[smfpyk6-1:0];
assign duox68l_r_f8nou99k2[smfpyk6-1:0] = ua3hwncs2rj394m9h37[smfpyk6-1:0];
assign n2y0qyph75pffp3dwwf80[smfpyk6-1:0] = u9eb3j3kbeih0qsei71[smfpyk6-1:0];
assign qfy5nt0fzqzm85nkaj[smfpyk6-1:0] = df7442xh1y14cj3o6qx[smfpyk6-1:0];

generate
if (smfpyk6 < 1024) begin : trtvthzs0bo5bhr0o62w9gwf70s
	assign u5p7r7vyhmyho6aa[1023:smfpyk6]    = {(1024-smfpyk6){1'b0}};
	assign duox68l_r_f8nou99k2[1023:smfpyk6]   = {(1024-smfpyk6){1'b0}};
	assign n2y0qyph75pffp3dwwf80[1023:smfpyk6] = {(1024-smfpyk6){1'b0}};
	assign qfy5nt0fzqzm85nkaj[1023:smfpyk6] = {(1024-smfpyk6){1'b0}};
end
endgenerate

wire   j3hs6x_gr14ms2c_qp91   = |ua3hwncs2rj394m9h37;

assign byyagfto1uztznf7eh  = hod7aki51hhxhaobdn | (~i_1o22g1okmq7xskth & u9eb3j3kbeih0qsei71);
assign hod7aki51hhxhaobdn = wxul7qtqbzvhly_rlbtr4lica;
assign i_1o22g1okmq7xskth = {smfpyk6{j3_0mc1_bfh0}} &  amjh0bop7ptd8znl3hi[smfpyk6-1:0];

assign dj_0z4kpnkm667my96de  = ywxqdtlc1lq30jgk8mu9;
assign pqteh7_cyvhhbcf4   = dc05a4etne0pkj7u9_nb;
assign gj_o1f7vjh3bs5_rkd65mtg = e6_o9xin1wu8kylws9m;
assign k68x_2_wxidbic0ld_     = l8d6kinl1s6rh6ha;
assign svgpgd1koc7jztn7h2     = s942sghng1f2y8;
assign cp0_pk_fscb9h1z      = pd9da145nlzxwlaua8;

assign ywxqdtlc1lq30jgk8mu9      = n2y0qyph75pffp3dwwf80[hnvgp5pvvjoaa527];
assign dc05a4etne0pkj7u9_nb      = qfy5nt0fzqzm85nkaj[hnvgp5pvvjoaa527];
wire   gds4le09zm4ap5uqms88_s = (hnvgp5pvvjoaa527 >= smfpyk6[9:0]);
wire   jozps8luysq4zqusxi0     = duox68l_r_f8nou99k2[hnvgp5pvvjoaa527];
wire   qp4697adqzamoa1l7o93     = ~u5p7r7vyhmyho6aa[hnvgp5pvvjoaa527];
wire   ja02quqb6_fw73n11w_l      =  u5p7r7vyhmyho6aa[hnvgp5pvvjoaa527];

ux607_gnrl_dffr #(1) pliwsgyugyhal96t1kxpi_175t (gds4le09zm4ap5uqms88_s , e6_o9xin1wu8kylws9m, gf33atgy, hfocw7va5_);

ux607_gnrl_dffr #(1) yt02lvyovf3udlzivjwe8_ (jozps8luysq4zqusxi0 , l8d6kinl1s6rh6ha, gf33atgy, hfocw7va5_);

ux607_gnrl_dffr #(1) qd8rizzzip9hzvzroq49 (qp4697adqzamoa1l7o93 , s942sghng1f2y8, gf33atgy, hfocw7va5_);

ux607_gnrl_dffr #(1) jfr_xh6zx_r9xymhy_glopj (ja02quqb6_fw73n11w_l , pd9da145nlzxwlaua8, gf33atgy, hfocw7va5_);





































assign r65hrblk6cfz_[31:27] = 5'd0;
assign r65hrblk6cfz_[26:24] = 3'd0;	
assign r65hrblk6cfz_[23]    = 1'd0;
assign r65hrblk6cfz_[22]    = 1'b1;	
assign r65hrblk6cfz_[21:20] = 2'd0;
assign r65hrblk6cfz_[19]    = ywxqdtlc1lq30jgk8mu9;
assign r65hrblk6cfz_[18]    = dj_0z4kpnkm667my96de;
assign r65hrblk6cfz_[17]    = dc05a4etne0pkj7u9_nb;
assign r65hrblk6cfz_[16]    = pqteh7_cyvhhbcf4;
assign r65hrblk6cfz_[15]    = e6_o9xin1wu8kylws9m;
assign r65hrblk6cfz_[14]    = gj_o1f7vjh3bs5_rkd65mtg;
assign r65hrblk6cfz_[13]    = l8d6kinl1s6rh6ha;
assign r65hrblk6cfz_[12]    = k68x_2_wxidbic0ld_;
assign r65hrblk6cfz_[11]    = s942sghng1f2y8;
assign r65hrblk6cfz_[10]    = svgpgd1koc7jztn7h2;
assign r65hrblk6cfz_[9]     = pd9da145nlzxwlaua8;
assign r65hrblk6cfz_[8]     = cp0_pk_fscb9h1z;
assign r65hrblk6cfz_[7]     = zy51q_pbb9tfrc_of;
assign r65hrblk6cfz_[6]     = qmur7eb6mi4y;
assign r65hrblk6cfz_[5]     = a5ee5u9gnomn5itad6c8;
assign r65hrblk6cfz_[4]     = dd2_ly9t687r6v_wa;
assign r65hrblk6cfz_[3:0]   = czyq3s7omblo1;


assign q7xpkacoiqp__elsg[31]    = 1'b0;
assign q7xpkacoiqp__elsg[30]    = 1'b0;
assign q7xpkacoiqp__elsg[29]    = 1'b0;	
assign q7xpkacoiqp__elsg[28]    = 1'b0;	
assign q7xpkacoiqp__elsg[27]    = 1'b0;
assign q7xpkacoiqp__elsg[26]    = 1'b0;	
assign q7xpkacoiqp__elsg[25:16] = hnvgp5pvvjoaa527;
assign q7xpkacoiqp__elsg[1]     = wse0ogbls179;

wire wgfaj9bbjo8xrhim;
wire h2nbgy9dwca7fcjfc6;

assign q7xpkacoiqp__elsg[0]     = h2nbgy9dwca7fcjfc6;
assign q7xpkacoiqp__elsg[4]     = wgfaj9bbjo8xrhim;
assign q7xpkacoiqp__elsg[3:2]   = 2'd0;
assign q7xpkacoiqp__elsg[15:5]  = 11'd0;

assign o59nl09azxaz = f_bjjlctco54pp3; 
assign nm83rtc_qty = wse0ogbls179; 

wire			jp0vvpklui3rxd2lpke313;
wire			eavu1m98r0wej0agclq01_27do;
wire			qigehcjj73tai4iqvn11v;
wire			krvdn1vymr7rwz7cp3fvd8di;

wire       [smfpyk6-1:0]	dyaqvcnm3xjd57ga;
wire       [smfpyk6-1:0]	tyg4te0t3o8p00bpz7m3;

assign dyaqvcnm3xjd57ga =   ({smfpyk6{jp0vvpklui3rxd2lpke313}} & amjh0bop7ptd8znl3hi[smfpyk6-1:0])
		       | (~({smfpyk6{qigehcjj73tai4iqvn11v}} & amjh0bop7ptd8znl3hi[smfpyk6-1:0]) & io5ukym11gp2utw);
assign tyg4te0t3o8p00bpz7m3 = (~f_bjjlctco54pp3) ? {smfpyk6{1'b0}} : dyaqvcnm3xjd57ga;

assign eavu1m98r0wej0agclq01_27do = ph7jz_7_o_welqv[0] & ph7jz_7_o_welqv[3] & k53u3hfcf_oxdneqvc;
assign krvdn1vymr7rwz7cp3fvd8di = ph7jz_7_o_welqv[0] & ph7jz_7_o_welqv[2] & k53u3hfcf_oxdneqvc;



ux607_gnrl_dffr #(smfpyk6) ijas7s58tl_jz5tom (tyg4te0t3o8p00bpz7m3 , io5ukym11gp2utw, gf33atgy, hfocw7va5_);

ux607_gnrl_dffr #(1)     m2xgz8727qawomlzvsdfwcai (eavu1m98r0wej0agclq01_27do , jp0vvpklui3rxd2lpke313, gf33atgy, hfocw7va5_);
ux607_gnrl_dffr #(1)     aa629_len9drtgpz3kgrbb26fhx (krvdn1vymr7rwz7cp3fvd8di , qigehcjj73tai4iqvn11v, gf33atgy, hfocw7va5_);

wire d0ddeoh4di2fegf = ph7jz_7_o_welqv[31] & ph7jz_7_o_welqv[0];
wire dlqbcohfwpnt989j0nz69m = ph7jz_7_o_welqv[30] & ph7jz_7_o_welqv[0];
wire [9:0] b3nao_oc31uvz0nru = ph7jz_7_o_welqv[25:16] & {10{ph7jz_7_o_welqv[0]}};
wire d86bb1j5ii3kdwg7yfqg = ph7jz_7_o_welqv[1] & ph7jz_7_o_welqv[0];

ux607_gnrl_dfflr #(1)    g_bvwhuwyadfif0sg8sisr  (k53u3hfcf_oxdneqvc, d0ddeoh4di2fegf  , f6umtn3v33g4  , gf33atgy, hfocw7va5_);
ux607_gnrl_dfflr #(1)    til9we_0t7_9fnz48tt9rp1e(k53u3hfcf_oxdneqvc, dlqbcohfwpnt989j0nz69m, i2r6o0rnjrg_t8c65, gf33atgy, hfocw7va5_);
ux607_gnrl_dfflr #(10)   p6cf_rxitij1_98164i  (k53u3hfcf_oxdneqvc, b3nao_oc31uvz0nru  , hnvgp5pvvjoaa527  , gf33atgy, hfocw7va5_);
ux607_gnrl_dfflr #(1)    knlgixfr_0vpjzin0l (k53u3hfcf_oxdneqvc, d86bb1j5ii3kdwg7yfqg , wse0ogbls179 , gf33atgy, hfocw7va5_);

wire jbb4reujnm78vxv3;
wire wp01tn3udyi;
wire hdgmfjosptbbbdrm;
wire ro10qraedfbfwyu;


  ux607_gnrl_sync # (
  .DP(2),
  .DW(1)
  ) xiswdbhmedbakiav7(
      .din_a    (v66uy2mvzfhls6   ),
      .dout     (jbb4reujnm78vxv3),
      .clk      (dk2xhkj77a        ),
      .rst_n    (hfocw7va5_        ) 
  );

assign wp01tn3udyi = jbb4reujnm78vxv3 & wgfaj9bbjo8xrhim;
ux607_gnrl_dffr #(1) he1p__6jv30rolixi (wp01tn3udyi, hdgmfjosptbbbdrm , dk2xhkj77a, hfocw7va5_);
assign ro10qraedfbfwyu = wp01tn3udyi ^ hdgmfjosptbbbdrm;

ux607_gnrl_dfflr #(1) cj5z3gi02_1efxcvnjf6e07 (k53u3hfcf_oxdneqvc, ph7jz_7_o_welqv[4], wgfaj9bbjo8xrhim, gf33atgy, hfocw7va5_);

wire o5ja8v5rdov6rjj80tjucm;
wire [14:0] wpxle7je_f7gca4ksk;
wire [14:0] fwskutqvos0y64s08oycuj2 = 
	(wgfaj9bbjo8xrhim == 1'b0 || b5xt1a6vsi17t78i == 1'b1)   ? {1'b0, {14{1'b0}}}: 
	(ro10qraedfbfwyu  == 1'b1 && o5ja8v5rdov6rjj80tjucm == 1'b0)? wpxle7je_f7gca4ksk + 1'b1: 
	                                                        wpxle7je_f7gca4ksk; 
ux607_gnrl_dffr #(14 + 1) x4fo_my5564_tw_xuf_30zu0m (fwskutqvos0y64s08oycuj2, wpxle7je_f7gca4ksk, dk2xhkj77a, hfocw7va5_);
assign o5ja8v5rdov6rjj80tjucm = wpxle7je_f7gca4ksk[14];

ux607_gnrl_dfflr #(1)    x1xy2p1gi52uyenka9j3d (k53u3hfcf_oxdneqvc, ph7jz_7_o_welqv[0]    , h2nbgy9dwca7fcjfc6, gf33atgy, hfocw7va5_);
assign f_bjjlctco54pp3 =   o5ja8v5rdov6rjj80tjucm? 1'b0: h2nbgy9dwca7fcjfc6;








































ux607_gnrl_dffr #(1)     cu2mh686avy5o5x9g567         (bf0mjxu4_jjk1oq , j3_0mc1_bfh0, gf33atgy, hfocw7va5_);
ux607_gnrl_dffr #(1)     gytrx8gkm60rtjlay_ougx77x3 (k53u3hfcf_oxdneqvc , prkl04ot6l0th2kjj3lensn, gf33atgy, hfocw7va5_);

















ux607_gnrl_dfflr #(smfpyk6)     o6lgren3tni7al0pgzadn7   (h90anyh0t2067aaxikbb  , xcl486gg7mcx74msnzz   , uxfmt_p8696p685   , gf33atgy, hfocw7va5_);
ux607_gnrl_dfflr #(smfpyk6)     l6woqnizbt2j05cyvxgms0lt (wv03_r28177pyhq87q_eku, g9_nradsie9gn_rr4o , c_d83vejsnlgx1b750 , gf33atgy, hfocw7va5_);
ux607_gnrl_dffrs #(smfpyk6)     cs232zc182_bina03bd1gx (je9cia8z8gc_arzaynhtmf, df7442xh1y14cj3o6qx    , gf33atgy, hfocw7va5_);
ux607_gnrl_dffr #(smfpyk6)      k2wqdvqyxcs1t_        (okvgcb6z3u4      , o0pri6gw33y, gf33atgy, hfocw7va5_);





























assign h90anyh0t2067aaxikbb    = prkl04ot6l0th2kjj3lensn | ~f_bjjlctco54pp3;
assign xcl486gg7mcx74msnzz    = ( amjh0bop7ptd8znl3hi[smfpyk6-1:0] & {smfpyk6{f6umtn3v33g4}}   & {smfpyk6{f_bjjlctco54pp3}})
                          | (~amjh0bop7ptd8znl3hi[smfpyk6-1:0] & uxfmt_p8696p685           & {smfpyk6{f_bjjlctco54pp3}})
			  ;
assign wv03_r28177pyhq87q_eku  = prkl04ot6l0th2kjj3lensn | ~f_bjjlctco54pp3;
assign g9_nradsie9gn_rr4o  = ( amjh0bop7ptd8znl3hi[smfpyk6-1:0] & {smfpyk6{i2r6o0rnjrg_t8c65}} & {smfpyk6{f_bjjlctco54pp3}})
                          | (~amjh0bop7ptd8znl3hi[smfpyk6-1:0] & c_d83vejsnlgx1b750         & {smfpyk6{f_bjjlctco54pp3}})
			  ;


wire  [1023:0] lrtmvfndgc0qjeri7vt = 1024'd1 << qvpivcc8d7j57jlwl[9:0];

assign r2vx5irgc6jszc2q1zg9 = lrtmvfndgc0qjeri7vt[smfpyk6-1:0] & c_d83vejsnlgx1b750[smfpyk6-1:0] & {smfpyk6{qcv2n1t0m8gvo5cto}};
assign tekott495862wlgwpec4r = (amjh0bop7ptd8znl3hi[smfpyk6-1:0] & {smfpyk6{i2r6o0rnjrg_t8c65 & prkl04ot6l0th2kjj3lensn}})	
                          | {smfpyk6{~f_bjjlctco54pp3}};
assign je9cia8z8gc_arzaynhtmf  = ~tekott495862wlgwpec4r & (df7442xh1y14cj3o6qx |  r2vx5irgc6jszc2q1zg9);

assign okvgcb6z3u4 = uxfmt_p8696p685 | k_g1vkidq8p8y6ghnxc4;

ux607_gnrl_dfflr #(10)     ybuxueg6wd1klv6mxra81x3nm4a (km788k575stdqjlb_qqfypq, tgw362y_u7jxvpdu2t3c , sv2fooskb173c3b58 , gf33atgy, hfocw7va5_);








wire [1023:0] yb654zmcg4h8c21uh3_xo8v1n;
assign yb654zmcg4h8c21uh3_xo8v1n[smfpyk6-1:0] =  c_d83vejsnlgx1b750[smfpyk6-1:0] & ~uxfmt_p8696p685[smfpyk6-1:0] & ~df7442xh1y14cj3o6qx[smfpyk6-1:0];

generate
if (smfpyk6 < 1024) begin : slwa97c5fe_l8qordzzd6eugg7hlrsz89cgb
	assign yb654zmcg4h8c21uh3_xo8v1n[1023:smfpyk6] = {(1024-smfpyk6){1'b0}};
end
endgenerate

assign v5ciuvu6m6lmww03 = yb654zmcg4h8c21uh3_xo8v1n[sv2fooskb173c3b58];

assign km788k575stdqjlb_qqfypq = ~f_bjjlctco54pp3 | (~v5ciuvu6m6lmww03 & |yb654zmcg4h8c21uh3_xo8v1n);
assign tgw362y_u7jxvpdu2t3c = (f_bjjlctco54pp3 & (rir_sifntdbcly7vezk338qsh3 != smfpyk6[9:0])) ?  rir_sifntdbcly7vezk338qsh3 : 10'd0;


assign tchrn3tov0okb6f[31:24] = 8'd0;
assign tchrn3tov0okb6f[23:20] = 4'd2;	
assign tchrn3tov0okb6f[19:17] = 3'd0;
assign tchrn3tov0okb6f[16]    = 1'b1;	
assign tchrn3tov0okb6f[15:12] = 4'd4;	
assign tchrn3tov0okb6f[11:0]  = {3'b000, qj3a7cq7w0bujncuh,2'b00};	

wire [1023:0] ghtqd4su_73qa2_mn843e;
wire [31:0]   vdgq54scrsea23 [31:0];
wire [31:0]   poaip4n8_6sk4wngow0k [31:0];
wire [31:0]   tm5axyn4g64fiyd0;
wire [31:0]   ssxbsxqu8jyx08tyf;



assign ghtqd4su_73qa2_mn843e[smfpyk6-1:0] = a7pselnd0w05duz_ivqvp[smfpyk6-1:0];

generate
if (smfpyk6 < 1024) begin : u94nir8u1qjx5kuduxv8g4ze0za4jg
	assign ghtqd4su_73qa2_mn843e[1023:smfpyk6] = {(1024-smfpyk6){1'b0}};
end
endgenerate

genvar i;
generate
	for (i=0; i<32; i=i+1) begin : y47ukd5nk5u11e
		assign vdgq54scrsea23[i] = ghtqd4su_73qa2_mn843e[i*32+32-1 : i*32];
		assign poaip4n8_6sk4wngow0k[i] = vdgq54scrsea23[i];
	end
endgenerate


assign ws9kutgi4r0wui1     = poaip4n8_6sk4wngow0k[hnvgp5pvvjoaa527[9:5]];




generate
	for (i=0; i<32; i=i+1) begin : v9cbwwfcr1b4c
		assign tm5axyn4g64fiyd0[i] = &poaip4n8_6sk4wngow0k[i];  
	end
endgenerate

assign ssxbsxqu8jyx08tyf = tm5axyn4g64fiyd0;
assign y80_gmc7mbs2g68     = (smfpyk6 > 32) ? ssxbsxqu8jyx08tyf : 32'b0;


assign rwyvi96_wuktwcs65     = 32'b0;


assign dr8lpark3fykgiqvl     = 32'b0;

assign s51p9m5pter6agwkfmi = 32'd0;
assign lu2p7m5sdkbd = 32'd0;


wire	[31:0]	c60vhelr4y2rwt9h_czqh   = yv13_lx8u9yhr8p6i;
wire	[31:0]	bq_nf94_buw8y4s71ahj_a_1t = d8panmbslrc4xeco;

assign stcjaa1sbc18df8[31:29] = 3'd0;
assign stcjaa1sbc18df8[28:24] = c60vhelr4y2rwt9h_czqh[4:0];
assign stcjaa1sbc18df8[23:13] = 11'd0;
assign stcjaa1sbc18df8[12]    = wl4tlno7ko;
assign stcjaa1sbc18df8[11]    = 1'b0;
assign stcjaa1sbc18df8[10:8]  = iro64ooeeusz4ro;
assign stcjaa1sbc18df8[7:5]  = 3'd0;
assign stcjaa1sbc18df8[4:0]  = bq_nf94_buw8y4s71ahj_a_1t[4:0];

wire       lp9sg9fpufpewvq4c = (~f_bjjlctco54pp3) | zlzdpgdm7uynjpt_tg;
wire [2:0] nzboxl6w7dnaie = (~f_bjjlctco54pp3) ? 3'd0 : b69xflf6dvza7n0;

ux607_gnrl_dfflr #(3)     v6h0xfsju50scc4w0f (lp9sg9fpufpewvq4c, nzboxl6w7dnaie , iro64ooeeusz4ro , gf33atgy, hfocw7va5_);







































wire jyrh1m9mjbf9l4drus = qcv2n1t0m8gvo5cto & (qvpivcc8d7j57jlwl[9:0] == aswynak3c52xoo5[9:0]);
wire tpiou8668hwj    = w6r9d62ex8olvrj0zfd7 & ((oq56n5j5gd3i2trf1n23 ? qvpivcc8d7j57jlwl[vmw6vavuv7md5-23:vmw6vavuv7md5-32] : qvpivcc8d7j57jlwl[9:0]) == aswynak3c52xoo5[9:0]);

wire qmc6cb9fgpzenmn5y1q = lypfqocyyrqu;
wire [pn11iufvnvon1yjbw-1:0] dfammclc11scjo = (k9ddbzzry2og0lep5n5t6dc37_ | hrxvvr_jkklnx6btx7) ? iyneurriss9qaw5wv5vz : sctcxvmp891m32rpg4w;

wire ln3j6633fy9dn0a9lzh = ebc4u4oafhzae;
wire [pn11iufvnvon1yjbw-1:0] qcvbxek5nak_3kg = umwi6wlplo34froaxm6t ? ldooojs2eemqgx70 : sctcxvmp891m32rpg4w;

wire sep9pg4c7osixv8n = kjd3v6ed24ptvm;
wire [pn11iufvnvon1yjbw-1:0] cc3x320l97fzil = lxnlpqnqclk48r5 ? p_n8ldx18y53b6dr_6 : ldooojs2eemqgx70;

wire ddkfjvirafklpe2n2ob = rknmpp444d3ijb;
wire [pn11iufvnvon1yjbw-1:0] cl1fukzehij9dr4 = tpiou8668hwj ? (iuasmef2ixpgpp9wrfgatqf ? i2hy3177smkb_6w99thp : sctcxvmp891m32rpg4w) : p_n8ldx18y53b6dr_6;

wire s_z38uf568t4qu9sim1 = y4o106ig3ae61;
wire [pn11iufvnvon1yjbw-1:0] gj3_s9piinfa55 = jyrh1m9mjbf9l4drus ? sctcxvmp891m32rpg4w : i2hy3177smkb_6w99thp;

assign ikkfsfp =   ({pn11iufvnvon1yjbw{qmc6cb9fgpzenmn5y1q  }} & dfammclc11scjo  )
                 | ({pn11iufvnvon1yjbw{ln3j6633fy9dn0a9lzh }} & qcvbxek5nak_3kg )
                 | ({pn11iufvnvon1yjbw{sep9pg4c7osixv8n   }} & cc3x320l97fzil   )
                 | ({pn11iufvnvon1yjbw{ddkfjvirafklpe2n2ob   }} & cl1fukzehij9dr4   )
                 | ({pn11iufvnvon1yjbw{s_z38uf568t4qu9sim1}} & gj3_s9piinfa55)
                 ;

assign bghtgz = ((~f_bjjlctco54pp3) | wse0ogbls179) ? sctcxvmp891m32rpg4w : ikkfsfp;


ux607_gnrl_dfflr #(pn11iufvnvon1yjbw) qzb2adc0i_qg (1'b1, bghtgz, yqdpagjrodj, gf33atgy, hfocw7va5_);

assign bfdnuw8phzaai12zaen = rknmpp444d3ijb & w3f078jh09ukd9z_24;
assign glencod3i3o7mjo7n25 = tpiou8668hwj | wse0ogbls179;
assign pqyrjnamrpuq0yq9ny4  = bfdnuw8phzaai12zaen | (~glencod3i3o7mjo7n25 & arfgqzn8b91r3e);

wire b8yd4qt8bkhjrkvp = (~f_bjjlctco54pp3) ? 1'b0 : pqyrjnamrpuq0yq9ny4;

ux607_gnrl_dffl #(1) qquxe3hnzsxo3os (1'b1, b8yd4qt8bkhjrkvp, arfgqzn8b91r3e, gf33atgy, hfocw7va5_);










assign k9ddbzzry2og0lep5n5t6dc37_ = src1s9kkdw9sn9kvu6z4 & !wl4tlno7ko & (iro64ooeeusz4ro == 3'd0);

wire o124_op876pzcfi01b = k9ddbzzry2og0lep5n5t6dc37_ | (~f_bjjlctco54pp3);
wire [31:0] orqx5c5dk3t30g8445 = (~f_bjjlctco54pp3) ? 32'b0 : hs4cmw6ypuuets98;

wire a0gjphesi80nf8t4lvia = k9ddbzzry2og0lep5n5t6dc37_ | (~f_bjjlctco54pp3);
wire [9:0] prfxgeshmxayfj9 = (~f_bjjlctco54pp3) ? 10'b0 : hnvgp5pvvjoaa527;












ux607_gnrl_dffl #(32) lm_z9rh3w7_v54ac7ieuh (o124_op876pzcfi01b, orqx5c5dk3t30g8445, hq9truyassja3d8s, gf33atgy, hfocw7va5_);
ux607_gnrl_dffl #(10) p49iopwglxv7f45aqpobn (a0gjphesi80nf8t4lvia, prfxgeshmxayfj9, aswynak3c52xoo5, gf33atgy, hfocw7va5_);

localparam nbonmp8swjf2mgut        = 3'd0;
localparam creudrkk5x09rp        = 3'd1;
localparam crbggp3xcrjnllx5k4g = 3'd2;
localparam xmmu_lvl5192zd0t   = 3'd3;
localparam cxyxb7iduoropwijhyb  = 3'd4;
localparam bx7mo2mgyawwbwslm       = 3'd7;

wire kkb1acu9jvs6z4mupj8g        = (src1s9kkdw9sn9kvu6z4 | hrxvvr_jkklnx6btx7 | ohlejrcx6cdwmphlr | pf4xyp48dd4kkmpy5ab | s6m193phbzzswom34s | xl9_scab2526apfj3i0f8vd6) & wl4tlno7ko;

assign i38u6n1ltlug0pip9m_ = (o2cn09h2l79zhpeg8t7t   &  krbd9wuik05rhl6vnfy5vh)
                          | (iuasmef2ixpgpp9wrfgatqf & ~krbd9wuik05rhl6vnfy5vh)
                          | (tbldq1rirf40guoxqqaheb   &  krbd9wuik05rhl6vnfy5vh);

wire agmfdaem7i7u_tfp = ebc4u4oafhzae & ~umwi6wlplo34froaxm6t;
wire yi5ch5xrql2ssq_xjs14 = w3f078jh09ukd9z_24;

wire [2:0] gc3n9et6yw79py = iro64ooeeusz4ro[2:0] & ~ph7jz_7_o_welqv[10:8];

assign zlzdpgdm7uynjpt_tg = bxgr20exryirwahrpndyb8w14mai | kkb1acu9jvs6z4mupj8g | agmfdaem7i7u_tfp | yi5ch5xrql2ssq_xjs14;
assign b69xflf6dvza7n0 = bxgr20exryirwahrpndyb8w14mai     ? gc3n9et6yw79py     :
		       (iro64ooeeusz4ro != 3'd0)   ? iro64ooeeusz4ro         :
		       kkb1acu9jvs6z4mupj8g        ? creudrkk5x09rp        :
		       yi5ch5xrql2ssq_xjs14   ? xmmu_lvl5192zd0t   :
		       ~xl9kvstr9tbbh6vaejjlks7bkz ? crbggp3xcrjnllx5k4g :
		       ~i38u6n1ltlug0pip9m_    ? cxyxb7iduoropwijhyb  :
						bx7mo2mgyawwbwslm;

assign k_g1vkidq8p8y6ghnxc4 = oht8t1ux9vjcpjl842vlmyq[smfpyk6-1:0] & {smfpyk6{(yqdpagjrodj == ldooojs2eemqgx70) & iuasmef2ixpgpp9wrfgatqf}};

assign krbd9wuik05rhl6vnfy5vh = |(a7pselnd0w05duz_ivqvp[smfpyk6-1:0] & oht8t1ux9vjcpjl842vlmyq[smfpyk6-1:0]);

assign qfk9f0qt00j7_h08dsa   = kjd3v6ed24ptvm | y4o106ig3ae61 | v5ciuvu6m6lmww03;
assign zsnjingqe8568rcb3etc0gud = (kjd3v6ed24ptvm | y4o106ig3ae61) ?  aswynak3c52xoo5 : sv2fooskb173c3b58;
assign eayknskh17rtgo6n7hxacs7  = ~kjd3v6ed24ptvm;

assign kg9c2fr3o4t1l2_udn[11:0]  = cluaz37po70qc66wuio;
assign kg9c2fr3o4t1l2_udn[15:12] = 4'd0;
assign kg9c2fr3o4t1l2_udn[31:16] = xmgisya42ikqz7vaea3lpoj;

generate
if (d8panmbslrc4xeco > 0) begin : f53coqlt0ckb140qbcc









        wire [d8panmbslrc4xeco-1:0] rv1hcr_7yt8876a1_jpo;
        wire [d8panmbslrc4xeco-1:0] snl7vxp_nf2hg7759nuls2kwi;
        wire u13o9kcllpgr756jrne2s420 = utec8wet9b5ke5gtbnr__oo1hi7395v;
        wire vsa1ioy4ls45okvn20aanrtutp = ~f_bjjlctco54pp3;
        wire dol8_l4yrxzfwdrdai2gtj9mch = u13o9kcllpgr756jrne2s420 | vsa1ioy4ls45okvn20aanrtutp;
        assign snl7vxp_nf2hg7759nuls2kwi = vsa1ioy4ls45okvn20aanrtutp ? {d8panmbslrc4xeco{1'b0}} : ph7jz_7_o_welqv[d8panmbslrc4xeco-1:0];
        ux607_gnrl_dffl #(d8panmbslrc4xeco)    pqy5kgyf32ytjj51eaxvl01n0  (dol8_l4yrxzfwdrdai2gtj9mch, snl7vxp_nf2hg7759nuls2kwi, rv1hcr_7yt8876a1_jpo, gf33atgy, hfocw7va5_);   
        assign cluaz37po70qc66wuio[d8panmbslrc4xeco-1:0]   = rv1hcr_7yt8876a1_jpo;
end
if (d8panmbslrc4xeco < 12) begin : am984i72yytt5vuvlxvmuxeq3z
	assign cluaz37po70qc66wuio[11:d8panmbslrc4xeco] = {(12-d8panmbslrc4xeco){1'b0}};
end
endgenerate

generate
if (yv13_lx8u9yhr8p6i > 0) begin : iwu334qxpanzbwbuzwvvu









        wire [yv13_lx8u9yhr8p6i-1:0] qo208zzbmp5xo6xd0y3dvm7s9;
        wire [yv13_lx8u9yhr8p6i-1:0] f9w70migyhh_t24gw67o5pmgtk2gqm;
        wire f7b9usnivlk584_5_k7xkordqdmccq = utec8wet9b5ke5gtbnr__oo1hi7395v;
        wire b4j_7fkuanfojsz9awcxq30_ljkqauo = ~f_bjjlctco54pp3;
        wire eiiql4vh9e2sqisryvcm5wqbw688c9 = f7b9usnivlk584_5_k7xkordqdmccq | b4j_7fkuanfojsz9awcxq30_ljkqauo;
        assign f9w70migyhh_t24gw67o5pmgtk2gqm = b4j_7fkuanfojsz9awcxq30_ljkqauo ? {yv13_lx8u9yhr8p6i{1'b0}} : ph7jz_7_o_welqv[(yv13_lx8u9yhr8p6i+16-1):16];
        ux607_gnrl_dffl #(yv13_lx8u9yhr8p6i)    ts5_skdjb8189qqk5uu253z8u  (eiiql4vh9e2sqisryvcm5wqbw688c9, f9w70migyhh_t24gw67o5pmgtk2gqm, qo208zzbmp5xo6xd0y3dvm7s9, gf33atgy, hfocw7va5_);
        assign xmgisya42ikqz7vaea3lpoj[yv13_lx8u9yhr8p6i-1:0] = qo208zzbmp5xo6xd0y3dvm7s9;
end
if (yv13_lx8u9yhr8p6i < 16) begin : jem2ui5s73d1tek9ab2005q_3p1h2ti7
	assign xmgisya42ikqz7vaea3lpoj[15:yv13_lx8u9yhr8p6i] = {(16-yv13_lx8u9yhr8p6i){1'b0}};
end
endgenerate

generate
if (d8panmbslrc4xeco > 0) begin : e8k15bror5jxl









wire [31:0] wpa8fofepv5mc4bm;
wire r9jq_n3uxzxc_n = heq7laaei2amn9igl2;
wire js4opspbn48g8o_6_ = ~f_bjjlctco54pp3;
wire j5e1idqvzaqsvomrk = r9jq_n3uxzxc_n | js4opspbn48g8o_6_;
assign wpa8fofepv5mc4bm = js4opspbn48g8o_6_ ? 32'b0 : xcgzxr3t0rc1243;

ux607_gnrl_dffl #(32)    eoz3b7jtog30ln  (j5e1idqvzaqsvomrk, wpa8fofepv5mc4bm, ajymk4x2v3, gf33atgy, hfocw7va5_);   
end
else begin : spayea75kbpdkcrkd2da45
	assign ajymk4x2v3 = 32'h0;
end
endgenerate

generate
if (d8panmbslrc4xeco > 1) begin : a5jiyfx4v3v7a









wire [31:0] j4i_a02nt9s1jazpo;
wire grr4fdk_k5hn5 = ldbdzv1slpkxnh;
wire tt72z6vyzoymwd46 = ~f_bjjlctco54pp3;
wire pc36ugbjnhr_zqyn = grr4fdk_k5hn5 | tt72z6vyzoymwd46;
assign j4i_a02nt9s1jazpo = tt72z6vyzoymwd46 ? 32'b0 : f0ggwdo3sb91;

ux607_gnrl_dffl #(32)    k3cjokxauvg4ql  (pc36ugbjnhr_zqyn, j4i_a02nt9s1jazpo, mlyn8clead, gf33atgy, hfocw7va5_);   
end
else begin : rifj8nqd6jd39j1ltym1n
	assign mlyn8clead = 32'h0;
end
endgenerate

generate
if (d8panmbslrc4xeco > 2) begin : sc1_fi8ah7zo65









wire [31:0] qkgg41flvh3z8;
wire zlglfnfynrfyd0h = r7195x8bumqznsl;
wire y2dq54n16clzikwibs = ~f_bjjlctco54pp3;
wire kjk3ty8x6kj7on = zlglfnfynrfyd0h | y2dq54n16clzikwibs;
assign qkgg41flvh3z8 = y2dq54n16clzikwibs ? 32'b0 : cz26a1huhfl0;

ux607_gnrl_dffl #(32)    yb7iwvzff164rqyf5h  (kjk3ty8x6kj7on, qkgg41flvh3z8, g2544euz9jpuu9, gf33atgy, hfocw7va5_);   
end
else begin : a_5irptbn70elegi1cps1ixs
	assign g2544euz9jpuu9 = 32'h0;
end
endgenerate

generate
if (d8panmbslrc4xeco > 3) begin : jsfl6kn4sug









wire [31:0] eh_8pem54alrt8;
wire emdq_pzlbxkrb = wputl8m_xeys6yd2_;
wire o6c320w1h6gf0 = ~f_bjjlctco54pp3;
wire yhlh3ux0xc0ky = emdq_pzlbxkrb | o6c320w1h6gf0;
assign eh_8pem54alrt8 = o6c320w1h6gf0 ? 32'b0 : v7on9ph3nyz9r0;

ux607_gnrl_dffl #(32)    e7h81e7kzbijto5vj8  (yhlh3ux0xc0ky, eh_8pem54alrt8, rw_eqfvro8, gf33atgy, hfocw7va5_);   
end
else begin : nbr7yggeidui44rf_4po31a
	assign rw_eqfvro8 = 32'h0;
end
endgenerate

generate
if (yv13_lx8u9yhr8p6i > 0) begin : h4mgqyh1ap3v









	wire [31:0] qe6q8vtd81px5fdd4dm;
	wire [31:0] h1r1e3yme6d2803x4qcqgc;
	wire x_vq6j7wrow94k8wg0z85cv2b = pize1u2oxu5xj00;
	wire qfr6_s0nept4ttu0bbxvz8 = ~f_bjjlctco54pp3;
	wire qv0arao_uvwvj6s8sb0y01 = x_vq6j7wrow94k8wg0z85cv2b | qfr6_s0nept4ttu0bbxvz8;
	assign h1r1e3yme6d2803x4qcqgc = qfr6_s0nept4ttu0bbxvz8 ? 32'b0 : k42ki1zy09wlmo2;
	ux607_gnrl_dffl #(32)    avetb7ssuno357vhlgdz  (qv0arao_uvwvj6s8sb0y01, h1r1e3yme6d2803x4qcqgc, qe6q8vtd81px5fdd4dm, gf33atgy, hfocw7va5_);   
	assign dmi_progbuf0 = qe6q8vtd81px5fdd4dm;
end
else begin : hub9h_9vy22jnqwamr4eer0h
	assign dmi_progbuf0 = axd20af5hznmm5;
end
endgenerate

generate
if (yv13_lx8u9yhr8p6i > 1) begin : tdvzq_pa4y0f3qni









	wire [31:0] awz652bc_sgy_rxi7;
	wire [31:0] zfekbezddye98jy1_8yrc1vfh;
	wire czbzajow3k0qkoqs7nt9ojm = oap_3j1l7iu77qz;
	wire u3_q7ig0_xm0en1qqrea = ~f_bjjlctco54pp3;
	wire iqx9r51u_tdko8oqarrwjz = czbzajow3k0qkoqs7nt9ojm | u3_q7ig0_xm0en1qqrea;
	assign zfekbezddye98jy1_8yrc1vfh = u3_q7ig0_xm0en1qqrea ? 32'b0 : y8bs2_4f4deqi4oqg;
	ux607_gnrl_dffl #(32)    bzf_9k7yt6j6aemjtblx96  (iqx9r51u_tdko8oqarrwjz, zfekbezddye98jy1_8yrc1vfh, awz652bc_sgy_rxi7, gf33atgy, hfocw7va5_);   
	assign i053jzqawhse = awz652bc_sgy_rxi7;
end
else begin : fmziwb5okvue8d151yewl7
	assign i053jzqawhse = axd20af5hznmm5;
end
endgenerate

generate
if (yv13_lx8u9yhr8p6i > 2) begin : wg_tlc34_vmnqsi4t









	wire [31:0] y1ykc1s0syzyajwoy7azm;
	wire [31:0] ezrfsvo7h40t52lle0_rfvp;
	wire raayv5c_g05m_o08ts1mzej = a1lc422n48q68c7;
	wire jwgq_s78l8cv12_b06idfd = ~f_bjjlctco54pp3;
	wire w6anmg21emi2og0lr39ndd0 = raayv5c_g05m_o08ts1mzej | jwgq_s78l8cv12_b06idfd;
	assign ezrfsvo7h40t52lle0_rfvp = jwgq_s78l8cv12_b06idfd ? 32'b0 : ho5oon65ncaswgb0lj5;
	ux607_gnrl_dffl #(32)    mn7v7ef1a3gm36apaa4ude  (w6anmg21emi2og0lr39ndd0, ezrfsvo7h40t52lle0_rfvp, y1ykc1s0syzyajwoy7azm, gf33atgy, hfocw7va5_);   
	assign tg3msrog_0bv = y1ykc1s0syzyajwoy7azm;
end
else begin : imkq7twgxtoon8x7iutuw4iql
	assign tg3msrog_0bv = axd20af5hznmm5;
end
endgenerate

generate
if (yv13_lx8u9yhr8p6i > 3) begin : i73on5yc4ki_wwxku









	wire [31:0] jgor81ql97tin6wl;
	wire [31:0] f45xuws1hbl0zlw9sziuk;
	wire j1kephsnnn_ttot22nxyu = yrsrzj9xgtahq9zah;
	wire w3tf7zsiutsun03yae9ap = ~f_bjjlctco54pp3;
	wire deydxh9yva6qndk5tjp95sz1r = j1kephsnnn_ttot22nxyu | w3tf7zsiutsun03yae9ap;
	assign f45xuws1hbl0zlw9sziuk = w3tf7zsiutsun03yae9ap ? 32'b0 : myuss9m1qp8gey0847r;
	ux607_gnrl_dffl #(32)    z5e8a8ltkn30gqep9ll  (deydxh9yva6qndk5tjp95sz1r, f45xuws1hbl0zlw9sziuk, jgor81ql97tin6wl, gf33atgy, hfocw7va5_);   
	assign g30pvzblnaf83zh = jgor81ql97tin6wl;
end
else begin : e7v01i3wma0q2tgw4ffdmoyw
	assign g30pvzblnaf83zh = axd20af5hznmm5;
end
endgenerate

generate
if (yv13_lx8u9yhr8p6i > 4) begin : r82dt15hekscfnean









	wire [31:0] qwy_h41h8d6fwxkh0;
	wire [31:0] chmxjhx_3jou2bsh2s57;
	wire t4o6qsuixop7u4tiiz8d3gt7 = a3ahayu4bahs;
	wire ckxl7omxo9_yxgep8iogqfruo = ~f_bjjlctco54pp3;
	wire g81nwl7vmf36c6eya6f4 = t4o6qsuixop7u4tiiz8d3gt7 | ckxl7omxo9_yxgep8iogqfruo;
	assign chmxjhx_3jou2bsh2s57 = ckxl7omxo9_yxgep8iogqfruo ? 32'b0 : axg6blt2b1j88hjl4_;
	ux607_gnrl_dffl #(32)    w7g4mlh5glmkbumf7m  (g81nwl7vmf36c6eya6f4, chmxjhx_3jou2bsh2s57, qwy_h41h8d6fwxkh0, gf33atgy, hfocw7va5_);   
	assign j2juyav34kkmuqd = qwy_h41h8d6fwxkh0;
end
else begin : pfrbfvt27v4ne25le_6w_nbq
	assign j2juyav34kkmuqd = axd20af5hznmm5;
end
endgenerate

generate
if (yv13_lx8u9yhr8p6i > 5) begin : xtoflf195rbbbn2









	wire [31:0] qezocale5gdsiq1dve;
	wire [31:0] gu2bog7gks5ism9fgeo3;
	wire ojmsplrq5tp65lg64p82 = jowfj_v52hdqypc;
	wire nj5sk5rwsdxpz012fskat2 = ~f_bjjlctco54pp3;
	wire n460l_h28pzkjb1gnnh9ry = ojmsplrq5tp65lg64p82 | nj5sk5rwsdxpz012fskat2;
	assign gu2bog7gks5ism9fgeo3 = nj5sk5rwsdxpz012fskat2 ? 32'b0 : l14fz29ful6_0ky8jl;
	ux607_gnrl_dffl #(32)    su01slzjr15pv6j3camnf  (n460l_h28pzkjb1gnnh9ry, gu2bog7gks5ism9fgeo3, qezocale5gdsiq1dve, gf33atgy, hfocw7va5_);   
	assign watz9oqgogsyjeo = qezocale5gdsiq1dve;
end
else begin : knwuxbkr5delfshw7t91vs5qk9
	assign watz9oqgogsyjeo = axd20af5hznmm5;
end
endgenerate

generate
if (yv13_lx8u9yhr8p6i > 6) begin : en2rnw9qhoko5pid









	wire [31:0] etyua9o05qdmvwi_ln4_;
	wire [31:0] yw5gu5_wildyh2e1bosv0;
	wire w947hub9x9pv_poajt6nw_e9g = zhrzwed1qf5xclzq0;
	wire jikvxlukftcnszhu3c4r9 = ~f_bjjlctco54pp3;
	wire nw1w_vu68omvlkwf23qqwbi = w947hub9x9pv_poajt6nw_e9g | jikvxlukftcnszhu3c4r9;
	assign yw5gu5_wildyh2e1bosv0 = jikvxlukftcnszhu3c4r9 ? 32'b0 : zzsj3yl_71x_1q2lh09b;
	ux607_gnrl_dffl #(32)    yl0e6jbe77bppfv3cmu2  (nw1w_vu68omvlkwf23qqwbi, yw5gu5_wildyh2e1bosv0, etyua9o05qdmvwi_ln4_, gf33atgy, hfocw7va5_);   
	assign kriizvysvcfvd = etyua9o05qdmvwi_ln4_;
end
else begin : oghvhizaluexlilgt7j2wfn
	assign kriizvysvcfvd = axd20af5hznmm5;
end
endgenerate

generate
if (yv13_lx8u9yhr8p6i > 7) begin : nqn7au0o0dyjk3oz









	wire [31:0] cjc77_489itlzftbb30;
	wire [31:0] zksw9d_3avz8wipzk6smli;
	wire dokt2qu1jjknqa6siwdumdan = e8i6of8n537o;
	wire aywikc_l_xtbcsdbxar55w6 = ~f_bjjlctco54pp3;
	wire h3yivlljkniy8ccttagjv7t = dokt2qu1jjknqa6siwdumdan | aywikc_l_xtbcsdbxar55w6;
	assign zksw9d_3avz8wipzk6smli = aywikc_l_xtbcsdbxar55w6 ? 32'b0 : vw8sa1crlzg24r4;
	ux607_gnrl_dffl #(32)    mkwohlqgwm92kmd_haf  (h3yivlljkniy8ccttagjv7t, zksw9d_3avz8wipzk6smli, cjc77_489itlzftbb30, gf33atgy, hfocw7va5_);   
	assign l97zx3ot2wagshr9 = cjc77_489itlzftbb30;
end
else begin : ditwpqq0yav_1euor7dvzn_2
	assign l97zx3ot2wagshr9 = axd20af5hznmm5;
end
endgenerate

generate
if (yv13_lx8u9yhr8p6i > 8) begin : jf4p3wkixbcc37pb0









	wire [31:0] fd5d0c5qn_cr48dza;
	wire [31:0] a98j2n5cz6d9ok52pfds4p1;
	wire cj_ow_snhn9sh3owfqeoeqe2e = h5cykrla39c8zlmr;
	wire n46mj4k5ziuljiy012tsnehoa = ~f_bjjlctco54pp3;
	wire oo3j_s5y4jak8eygiezbsqm = cj_ow_snhn9sh3owfqeoeqe2e | n46mj4k5ziuljiy012tsnehoa;
	assign a98j2n5cz6d9ok52pfds4p1 = n46mj4k5ziuljiy012tsnehoa ? 32'b0 : e0nj0rk_rp0knkls;
	ux607_gnrl_dffl #(32)    wnhvrtx9d_vhedsc78n5f  (oo3j_s5y4jak8eygiezbsqm, a98j2n5cz6d9ok52pfds4p1, fd5d0c5qn_cr48dza, gf33atgy, hfocw7va5_);   
	assign heiy5swkajxipcai = fd5d0c5qn_cr48dza;
end
else begin : c9ljhylqjjtf915vkvwhmpsw4oq
	assign heiy5swkajxipcai = axd20af5hznmm5;
end
endgenerate

generate
if (yv13_lx8u9yhr8p6i > 9) begin : mzanpak2u5v0









	wire [31:0] ilqrtadbxc5plrd0zm;
	wire [31:0] kjda_dy1oocmtnvntlo15m;
	wire vni7_daoeoz23ddng46hqacy = iwmac56d70_7;
	wire aqhi4t0_n2awyb3xw4od = ~f_bjjlctco54pp3;
	wire xkvimq9a6vycta3a1c42c = vni7_daoeoz23ddng46hqacy | aqhi4t0_n2awyb3xw4od;
	assign kjda_dy1oocmtnvntlo15m = aqhi4t0_n2awyb3xw4od ? 32'b0 : r_tf74b2bwwlb6s1wi;
	ux607_gnrl_dffl #(32)    opt_mrl3mn82s9182pnq6  (xkvimq9a6vycta3a1c42c, kjda_dy1oocmtnvntlo15m, ilqrtadbxc5plrd0zm, gf33atgy, hfocw7va5_);   
	assign etxdm_c986j2h = ilqrtadbxc5plrd0zm;
end
else begin : ul_6hqe2iklycmlhc7ijg3he
	assign etxdm_c986j2h = axd20af5hznmm5;
end
endgenerate

generate
if (yv13_lx8u9yhr8p6i > 10) begin : l2k0os6yjoebbhmez









	wire [31:0] uc0rvlnsz8o7_e3gv;
	wire [31:0] pd605484f4b717w3vbp9w;
	wire qs5uj20nikv1kdi63cc79 = fbcol2fiz4_dakl6;
	wire dvbe_if1418e5f2mtwn20sez4 = ~f_bjjlctco54pp3;
	wire wjgotxegsk4rv9za6hgiutr2oq = qs5uj20nikv1kdi63cc79 | dvbe_if1418e5f2mtwn20sez4;
	assign pd605484f4b717w3vbp9w = dvbe_if1418e5f2mtwn20sez4 ? 32'b0 : xade4a80z8ri9n6tfuin4;
	ux607_gnrl_dffl #(32)    szkmr19ojqqm1hx9_87967  (wjgotxegsk4rv9za6hgiutr2oq, pd605484f4b717w3vbp9w, uc0rvlnsz8o7_e3gv, gf33atgy, hfocw7va5_);   
	assign iw9ukx193kjidkn = uc0rvlnsz8o7_e3gv;
end
else begin : gvqruao06_bkn0wvnvlybud_
	assign iw9ukx193kjidkn = axd20af5hznmm5;
end
endgenerate

generate
if (yv13_lx8u9yhr8p6i > 11) begin : t0mvoq0cnoxq53i6









	wire [31:0] b8l5jwkx6198m97ihdr;
	wire [31:0] ulcduqialh2qylqsqq7tpzxx;
	wire h59uththpyzf5m6v1cn8z5wiph = okw64jbuomhjb3l9he;
	wire feo6hkovaxpdmfux07ra4sroyg = ~f_bjjlctco54pp3;
	wire n8y_z8v7i0r_f04akni8v = h59uththpyzf5m6v1cn8z5wiph | feo6hkovaxpdmfux07ra4sroyg;
	assign ulcduqialh2qylqsqq7tpzxx = feo6hkovaxpdmfux07ra4sroyg ? 32'b0 : s6ecnce9dbhjl8lyg3s7s;
	ux607_gnrl_dffl #(32)    fkt7njei2t6vgkehjea  (n8y_z8v7i0r_f04akni8v, ulcduqialh2qylqsqq7tpzxx, b8l5jwkx6198m97ihdr, gf33atgy, hfocw7va5_);   
	assign hwwlvkrpw_rd1 = b8l5jwkx6198m97ihdr;
end
else begin : v7c5wg7afj47m_mvkyicufh
	assign hwwlvkrpw_rd1 = axd20af5hznmm5;
end
endgenerate

generate
if (yv13_lx8u9yhr8p6i > 12) begin : dc2ay7lr8f6vniz9dm









	wire [31:0] tim3s8_3w3sskbq_68ajj;
	wire [31:0] p2m97fa4jf06jb4dlf9x4wnmd;
	wire p7nzvfgaeowekms05lyy1bs = xdx6hvlnkbknoa_m;
	wire a3wpnjclcf41sukcsozhcs = ~f_bjjlctco54pp3;
	wire m_1cjt8g6cho1yvhw37gu = p7nzvfgaeowekms05lyy1bs | a3wpnjclcf41sukcsozhcs;
	assign p2m97fa4jf06jb4dlf9x4wnmd = a3wpnjclcf41sukcsozhcs ? 32'b0 : rfhaugdrqwldacohp91;
	ux607_gnrl_dffl #(32)    wcjjdniqo8f0xbz0nz6m7  (m_1cjt8g6cho1yvhw37gu, p2m97fa4jf06jb4dlf9x4wnmd, tim3s8_3w3sskbq_68ajj, gf33atgy, hfocw7va5_);   
	assign b81eb_9kn7xgu725 = tim3s8_3w3sskbq_68ajj;
end
else begin : jky6xgptu8u2hymqaxbi82w
	assign b81eb_9kn7xgu725 = axd20af5hznmm5;
end
endgenerate

generate
if (yv13_lx8u9yhr8p6i > 13) begin : sd_yggqk61_oztavq









	wire [31:0] i08fbp3msw2y3z_0z;
	wire [31:0] r0rjdm5_vlxlwbndmh8cn;
	wire ab1sbtrz74nfr620lck1t3fdu = dzcjaphosa9ch;
	wire d8x87v42_ce88oex3byjxo0u_ = ~f_bjjlctco54pp3;
	wire r33j0f7ga679l_5uvafrzs3 = ab1sbtrz74nfr620lck1t3fdu | d8x87v42_ce88oex3byjxo0u_;
	assign r0rjdm5_vlxlwbndmh8cn = d8x87v42_ce88oex3byjxo0u_ ? 32'b0 : e1ptokxdw97811mlgkh;
	ux607_gnrl_dffl #(32)    iadj3yyzjy4df4_9a4a3  (r33j0f7ga679l_5uvafrzs3, r0rjdm5_vlxlwbndmh8cn, i08fbp3msw2y3z_0z, gf33atgy, hfocw7va5_);   
	assign rj3ujsskxnsw3 = i08fbp3msw2y3z_0z;
end
else begin : pfawa6b51sh02kinexdv3o0l
	assign rj3ujsskxnsw3 = axd20af5hznmm5;
end
endgenerate

generate
if (yv13_lx8u9yhr8p6i > 14) begin : y0sdhaeej20xzr









	wire [31:0] bd6aymk92snjoqmny;
	wire [31:0] pmz9xmgb4jm18t0056ew7z13;
	wire o7vmc2gdqnv5b7jhcz5jr5xe = dxhr63c235702bgyoa;
	wire hh6vv2r5ej0_x7dgyj4fg = ~f_bjjlctco54pp3;
	wire yy4o6fshdqqe6_tqvxo0j = o7vmc2gdqnv5b7jhcz5jr5xe | hh6vv2r5ej0_x7dgyj4fg;
	assign pmz9xmgb4jm18t0056ew7z13 = hh6vv2r5ej0_x7dgyj4fg ? 32'b0 : ly2r1ofg_z2vx4ron71;
	ux607_gnrl_dffl #(32)    b2hvdksd_58ni0hvff  (yy4o6fshdqqe6_tqvxo0j, pmz9xmgb4jm18t0056ew7z13, bd6aymk92snjoqmny, gf33atgy, hfocw7va5_);   
	assign fp511hjp_uccxk4 = bd6aymk92snjoqmny;
end
else begin : g8tzy7vvvq92qmr7tqryrlfi
	assign fp511hjp_uccxk4 = axd20af5hznmm5;
end
endgenerate

generate
if (yv13_lx8u9yhr8p6i > 15) begin : hi9fatevmzg3fbw3m









	wire [31:0] t4hfbwcy0flj4nwzol;
	wire [31:0] gx27urorckh49sygbj8k3;
	wire o4iphbo705ph_pwrjrhef_hf = kt7so0oerx68ydrpz;
	wire t5qjpe73j3j0_ob_8tay8e4ftl = ~f_bjjlctco54pp3;
	wire ywwbvqkt7x13fcwkrkxd11qj = o4iphbo705ph_pwrjrhef_hf | t5qjpe73j3j0_ob_8tay8e4ftl;
	assign gx27urorckh49sygbj8k3 = t5qjpe73j3j0_ob_8tay8e4ftl ? 32'b0 : zx1kehbfsf4fsgtm5;
	ux607_gnrl_dffl #(32)    asdu4xot08z_cedp630fa  (ywwbvqkt7x13fcwkrkxd11qj, gx27urorckh49sygbj8k3, t4hfbwcy0flj4nwzol, gf33atgy, hfocw7va5_);   
	assign dde_945nq4horxo = t4hfbwcy0flj4nwzol;
end
else begin : eyg1ynpkjqbozjddchjb4lywz27e
	assign dde_945nq4horxo = axd20af5hznmm5;
end
endgenerate

































































































































































































































































































































































































































































































































































































































































































































































    
    
    
    
    
    
    localparam nssj8f0leerxslqz4v8f   = ((x5jl_73d_gruzgtcqu >=8));
    localparam t7jihcw5qjd4jvy9zkj  = ((x5jl_73d_gruzgtcqu >=16));
    localparam qf78j99hr5frn3oel037nu6  = ((x5jl_73d_gruzgtcqu >=32));
    localparam suokhv_cmzokm2mfitte  = ((x5jl_73d_gruzgtcqu >=64));
    localparam hyiaal7cwi_arst3fu0ui6x = ((x5jl_73d_gruzgtcqu >=128));
    localparam coskgmnlindpe = uaue4a0q4yu2u48[6:0];
    localparam d6fo1cizl8a07v1hoq17k   = 3'd0;
    localparam z68iccz0j602b2m9uekd7utr  = 3'd1;
    localparam tzfebftjmirx__sl5mroslq  = 3'd2;
    localparam obhfbd2skwiz5h4ycuhz8qc  = 3'd3;
    localparam nflkoqm4ystz_8qmgpml7smfy = 3'd4;
    
    genvar ly3dor8, mijwlia0, oily7;
    
    wire		f7d3dgllmdd700u391;
    wire		codzot9zq_4cz1;
    wire	[2:0]	yl_oakyedt10di1;
    
    wire		nijvffj_k83iteeb61;
    wire		y98wkjik72p2pi;
    wire	[127:0]	z1h6n4git1qfcautzkf7d;
    wire	[127:0]	sb0_ui0s9qs02p22r_1;
    wire	[127:0]	p1dv438hc3p6b3cc_o;
    wire		qdso0sntbt33twwh90;
    
    wire		t_wng_z1d0pxhdoop;
    wire		m9yqdzp8_4fxtud;
    wire		u_jpz86m2q4328du_;
    wire		jtszu4eoodrwh;
    wire		w_0muls__b8v_;
    wire		mtlruvvjhcvzf6;
    wire		zs1r9hd1d1_p;
    wire		xkda0fom0vel4oensw7;
    wire		i4oiz2wl_m8q5y00l76bwi;
    wire		kp5ybypb04805jmkg3619oh3s8;
    wire		jfo4e1ypekb5lfzzx39_4ru0;
    
    assign f7d3dgllmdd700u391    = gsmp8y890cng[20];
    assign codzot9zq_4cz1    = gsmp8y890cng[15];
    assign yl_oakyedt10di1	 = gsmp8y890cng[19:17];
    assign u_jpz86m2q4328du_	 = codzot9zq_4cz1 & j0d0ajxf_i5ihg3yt95;
    assign t_wng_z1d0pxhdoop	 = f7d3dgllmdd700u391 & od6u7rr1fxvo091a298;
    assign jtszu4eoodrwh	 = gvbp1k6dl4r0o3hg6n & ~zs1r9hd1d1_p;
    assign w_0muls__b8v_	 = (u_jpz86m2q4328du_ | m9yqdzp8_4fxtud) & ~zs1r9hd1d1_p;  
    assign mtlruvvjhcvzf6    = (jtszu4eoodrwh | w_0muls__b8v_);
    assign zs1r9hd1d1_p	 = (|gsmp8y890cng[14:12]) | gsmp8y890cng[22];
    
    assign p1dv438hc3p6b3cc_o  = {e7wcd07jh85sk_hny6, bxlgqasel4nu6fjtmnt, zbawca6o200bvbpa1b6, y2bt8u7bruuxsctix};

    
    assign jfo4e1ypekb5lfzzx39_4ru0 = (~f_bjjlctco54pp3) | (k53u3hfcf_oxdneqvc & ~ph7jz_7_o_welqv[0]);

    ux607_gnrl_dfflr #(1)  ogd1v8_p2oah2oxa1cwzw(1'b1, t_wng_z1d0pxhdoop, m9yqdzp8_4fxtud, gf33atgy, hfocw7va5_);

    
    
    wire h5maomnmovgqtb7 = fkm9up63o1aeauaqhjb & to_1lv9wnb3vmu6tvz5rc;
    wire jlwst2h0gt_6sp4da7gy = mtlruvvjhcvzf6 & ~xkda0fom0vel4oensw7 & ~jfo4e1ypekb5lfzzx39_4ru0;
    wire np3rynbqfba2mhmaun = h5maomnmovgqtb7 | jfo4e1ypekb5lfzzx39_4ru0;
    wire mldtc9sn3m60x9eriw8l = jlwst2h0gt_6sp4da7gy | np3rynbqfba2mhmaun;
    wire kx6z_pkj5wh_h7itxw = jlwst2h0gt_6sp4da7gy | (~np3rynbqfba2mhmaun);
    wire y0mgg9563m7xd4dskx;

    ux607_gnrl_dfflr #(1)   hycfz6ca4__q_27i9gh(mldtc9sn3m60x9eriw8l, kx6z_pkj5wh_h7itxw, y0mgg9563m7xd4dskx, gf33atgy, hfocw7va5_);
    
    assign fkm9up63o1aeauaqhjb = y0mgg9563m7xd4dskx;

    
    generate
	for (mijwlia0 = 0; mijwlia0 < uaue4a0q4yu2u48; mijwlia0=mijwlia0+32) begin: ynfao2sqi01suenjeegep_nu3ixh3dn_e7
		if ((mijwlia0+32) > uaue4a0q4yu2u48) begin: w4zpdu7boerc0qgii4k
			assign ju1kbeplcqy314lfj4[uaue4a0q4yu2u48-1:mijwlia0] = p1dv438hc3p6b3cc_o[uaue4a0q4yu2u48-1:mijwlia0];
		end
		else begin: g2tj0mp44e0uoxjsml4u
			assign ju1kbeplcqy314lfj4[(mijwlia0+31):mijwlia0] = p1dv438hc3p6b3cc_o[(mijwlia0+31):mijwlia0];
		end
	end
    endgenerate

    
    wire t8mvp5u93cjjm46h96 = jtszu4eoodrwh & ~xkda0fom0vel4oensw7 & ~jfo4e1ypekb5lfzzx39_4ru0;
    wire l1re437rmtafyidg_d9i6 = h5maomnmovgqtb7 | jfo4e1ypekb5lfzzx39_4ru0;
    wire yri8j450f6yd15apx06an = t8mvp5u93cjjm46h96 | l1re437rmtafyidg_d9i6;
    wire xnkju15pbe57c605uih = t8mvp5u93cjjm46h96 | (~l1re437rmtafyidg_d9i6);
    wire wit2mn0vwyc6onh0rc;

    ux607_gnrl_dfflr #(1)   voftzz7jdk6n483wflv4ypkl(yri8j450f6yd15apx06an, xnkju15pbe57c605uih, wit2mn0vwyc6onh0rc, gf33atgy, hfocw7va5_);
	
    assign r985fbe5k7hgzaq9i = ~wit2mn0vwyc6onh0rc;

    wire begwifcc9uvdqcg58d7rdxg8 = h5maomnmovgqtb7 | jfo4e1ypekb5lfzzx39_4ru0;
    wire sysgroia33amo29u859qc6qb;
    
    ux607_gnrl_dfflr #(1)   y8fgvm0oig9gdwg82lkmgh0m9j15l7(begwifcc9uvdqcg58d7rdxg8, wit2mn0vwyc6onh0rc, sysgroia33amo29u859qc6qb, gf33atgy, hfocw7va5_);
	
    
    assign bb04gpwotp2s6c7_p1gqkq = st4f16aums5; 

    
    assign sqmey185cu3mtixhl = p05ld2ghmwh; 

    
    assign rffcsd1o699ytclmx = 1'b1;  

    
    generate
	for (ly3dor8 = 0; ly3dor8 < x5jl_73d_gruzgtcqu; ly3dor8 = ly3dor8+32) begin: kahh1n4_12oqaw2yngibs48uxiziy6fd3
		assign lbr88vbqtg8rht7320frde[(ly3dor8+31):ly3dor8] = sb0_ui0s9qs02p22r_1[(ly3dor8+31):ly3dor8];
	end
    endgenerate

    
    wire [2:0]  ogc4vnz46z9rgvvncyy76lzb1 = (x5jl_73d_gruzgtcqu == 32) ? {1'b0,p1dv438hc3p6b3cc_o[1:0]} : p1dv438hc3p6b3cc_o[2:0];
    wire [15:0] sujr5m8l4oxl6iwk31;
    assign sujr5m8l4oxl6iwk31 = (yl_oakyedt10di1[1:0] == 2'b00) ? (16'h0001 <<  ogc4vnz46z9rgvvncyy76lzb1[2:0]) : 
                               (yl_oakyedt10di1[1:0] == 2'b01) ? (16'h0003 << {ogc4vnz46z9rgvvncyy76lzb1[2:1], 1'b0}) :
                               (yl_oakyedt10di1[1:0] == 2'b10) ? (16'h000f << {ogc4vnz46z9rgvvncyy76lzb1[2:2], 2'b0}) :
                               (yl_oakyedt10di1[1:0] == 2'b11) ? (16'h00ff) :
                               16'h0;

    assign g7qq38mx3d58n1b15kcia = wit2mn0vwyc6onh0rc ? sujr5m8l4oxl6iwk31[8-1:0] : 8'b0;

    
    assign demg_fwfkmaeawq30t = 1'b0; 

    
    assign grtb6ypa0px2gi1c = 1'b0; 

    
    assign f128d8ws0seoihu1 = yl_oakyedt10di1[1:0]; 

    
    wire kgv6f0xs6zr5ne3lzaw = m2r7mfmq3afdd1ine & nhafiywg3hg_52kogwh;
	assign nijvffj_k83iteeb61 = kgv6f0xs6zr5ne3lzaw;
	assign y98wkjik72p2pi   = xrqayy6vigrw66z8a;
	assign qdso0sntbt33twwh90 = kgv6f0xs6zr5ne3lzaw & (~sysgroia33amo29u859qc6qb);

    
    assign nhafiywg3hg_52kogwh = 1'b1; 

    
    wire [127:0] hqt6iij0v5y9iz0du4f_k;
    generate
	for (oily7 = 0; oily7 < 128; oily7=oily7+32) begin: ona78a__wof6ge1o2rhx98rf5h1na
		if (oily7 < x5jl_73d_gruzgtcqu) begin: n8p9u3x3it2fanvruq1z46lp6u21
			assign hqt6iij0v5y9iz0du4f_k[(oily7+31):oily7] = drz92qecqx_qtxwro[(oily7+31):oily7];
		end
		else begin: vbj6gcpt5a5xnwn9tfvw1vwau8b_xu1w1
			assign hqt6iij0v5y9iz0du4f_k[(oily7+31):oily7] = drz92qecqx_qtxwro[31:0];
		end
	end
    endgenerate
	assign z1h6n4git1qfcautzkf7d[31:0]   = hqt6iij0v5y9iz0du4f_k[31:0];
	assign z1h6n4git1qfcautzkf7d[63:32]  = hqt6iij0v5y9iz0du4f_k[63:32];
	assign z1h6n4git1qfcautzkf7d[95:64]  = hqt6iij0v5y9iz0du4f_k[95:64];
	assign z1h6n4git1qfcautzkf7d[127:96] = (x5jl_73d_gruzgtcqu == 64) ? hqt6iij0v5y9iz0du4f_k[63:32] : hqt6iij0v5y9iz0du4f_k[127:96];


	reg  [31:0] om4i8b1g4ffpkkjkse91;   
	reg  [31:0] sf14ab4y4pwg9uzf7ei;   
	reg  [31:0] at1z83ksz098eaaw45zorq;   
	reg  [31:0] pmxmx6g704kt9ffe_k3gsb4;   
	reg  [31:0] ln0owurz2hrjqyzt;      
	reg  [31:0] jy3u2zz45w3qt2o8ueas;      
	reg  [31:0] riur0xm9vgi7prn;      
	reg  [31:0] g4n2d80tx347g5d;      

	wire [31:0] cf1p9na3s94mkxr663b;
	wire [31:0] b2kif3s0l5f10gxlqp;
	wire [31:0] chxwpklhgug7nuaerfmj;
	wire [31:0] vhvg6pli9i9rtyr0gpued;
	wire [31:0] asuxi27dz56cq9qk1q6;
	wire [31:0] shq4l11_gkpyac;
	wire [31:0] zaqsdqqsq29r81i;
	wire [31:0] lbwqg4gjtgckn2f;
	wire [31:0] j3chbw93vus855iltfv4p;
	wire [31:0] d6y6mbjwlwbautf9;
	wire [31:0] a2uofg5xxki0oe1xex155;
	wire [31:0] cjg6agdce9fgz9d1hl0v;
	reg  [31:0] xwe5116fdnncgl5_idf0q;
	wire [31:0] xoviomvc7o7y87p3yap;
	wire [31:0] rfdqkys5p2ujup5_mm2n;
	wire [31:0] owcemq5_leom8y6ncl;

	wire [2:0]	xuzpr_ag_zzjjlhleh = 3'd1;
	reg		    shsgn99xfgm_falbwej9r;
	reg		    dlgkkhcodyhtm4ue;
	reg		    erplkdk9eejnm26v2q9axu;
	reg	 [2:0]	a91q0mpju3lvvuyy;
	reg		    sbn67m1e906fpvnin8pxq;
	reg		    c9fbc2_3b0q24_wa9w84pk;
	reg	 [2:0]	nwrntu_ns6js9tio;
	wire [6:0]	kz_vf5v7hkz3     = coskgmnlindpe;
	wire		ntt3vblrcouy6if54la = hyiaal7cwi_arst3fu0ui6x;
	wire		l36ob57itxhda2q  = suokhv_cmzokm2mfitte;
	wire		jij19fj8jksetx4  = qf78j99hr5frn3oel037nu6;
	wire		ivo3nt6en_d1s4fnn  = t7jihcw5qjd4jvy9zkj;
	wire		msljxv405r4t1rbl   = nssj8f0leerxslqz4v8f;

	wire		q3jh_tep8g0mk7m2ohvp;
	wire		gw5bpkb0gwli80bq;
	wire		p60i1235jw07wggo07zuxm;
	wire [2:0]	c9jvr8hzwcs0svgzgj4x;
	wire		nkqcgp9gxttikxmttl77t7sx;
	wire		z1uojli46j34r_32meos9;

	wire [2:0]	szmaji702081lti_h0qux;
	wire		vcedcqevwspfk05rtor3;
	wire		zzzclorwnw16vf8;
	wire		u5mjc2lh222oaobj;
	wire		btob5wz940x35dypuh;
	wire		hyqrpuxs_jhuma9ai4f9f;
	wire		dnah6nc0fw8ts_1ltvjz;
	wire [4:0]	wvyzyntlw4ro36s310tyw;

	wire [2:0]	bjkw1ffrzjhax1g63pke;
	wire		pnghshojyfxwjqjregrnf;

	wire		ssay1k38w94lso_;

	wire		alpkrgsdgm3z2_llqs9wc;
	wire		h7bf8fgzcxv2nr5q_g4nygf5c;
	wire		xt_seq2pq4js8rmtsz;
	wire		idbkyxhyplh8ik16cau;
	
	wire [127:0] elm1vif4d_10b1_g8_2;
	wire [127:0] jd3bx8g5usv4rwh4;
	wire [31:0]	z8heidfnfd6oy8;
	wire		doaxea8vme8i1z;
	wire		xuea1_k_eg81xsp7;
	wire		ub0do2eia4_zpjgutcd;
	wire		ooobnffsf8o6qo9i;
	wire		wlhp1d9_0qsm5__;
	wire		zz9n5bfhur01yx;
	wire		w2bzlpz5nmwdb2d;
	wire		tdjiiekyziosyf;
	wire		p6rade23wlwj8tphay;
	wire		qrsc_8c1f0s50ogii;
	wire		hehn594ckxi95te8;
	wire		czya52zksuaqev;

	reg	 [15:0]	cn8y8j2rziuq8l;
	wire [15:0]	z54sfjatc1sac9pfiv;
	reg		    k8f9lz_optfi4vcf;
	reg		    u3x9iybnpf8suar92;
	reg		    sb57m7q7jimdmg_;
	reg		    op9rx4p45h29r;
	wire		s93zuexjncoy1wmij4u;
	wire		d5g9bjqnj4hlkaa8tl1v;
	wire		q1o9g4lcei7dy3z1;
	wire		tljwcx5n4m9ruiltki;
	wire		otd6qmzkpph;
	wire [31:0]	vkb6t1zon4pxe;
	wire [31:0]	a0o2jippaa1o7rp5;
	wire [31:0]	cguui3s6gp4x7;
	wire [31:0]	rbaif3vx037msdnd;

	always @(posedge gf33atgy or negedge hfocw7va5_) begin
		if (!hfocw7va5_) begin
			dlgkkhcodyhtm4ue	 <= 1'b0;
			shsgn99xfgm_falbwej9r <= 1'b0;
		end
		else if (jfo4e1ypekb5lfzzx39_4ru0) begin
			dlgkkhcodyhtm4ue	 <= 1'b0;
			shsgn99xfgm_falbwej9r <= 1'b0;
		end
		else begin
			dlgkkhcodyhtm4ue	 <= gw5bpkb0gwli80bq;
			shsgn99xfgm_falbwej9r <= q3jh_tep8g0mk7m2ohvp;
		end
	end

	always @(posedge gf33atgy or negedge hfocw7va5_) begin
		if (!hfocw7va5_) begin
			nwrntu_ns6js9tio	 <= 3'd0;
		end
		else if (jfo4e1ypekb5lfzzx39_4ru0) begin
			nwrntu_ns6js9tio	 <= 3'd0;
		end
		else if (pnghshojyfxwjqjregrnf) begin
			nwrntu_ns6js9tio	 <= bjkw1ffrzjhax1g63pke;
		end
	end

	always @(posedge gf33atgy or negedge hfocw7va5_) begin
		if (!hfocw7va5_) begin
			erplkdk9eejnm26v2q9axu    <= 1'b0;
			a91q0mpju3lvvuyy	     <= tzfebftjmirx__sl5mroslq;
			sbn67m1e906fpvnin8pxq <= 1'b0;
			c9fbc2_3b0q24_wa9w84pk    <= 1'b0;
			u3x9iybnpf8suar92	     <= 1'b0;
			sb57m7q7jimdmg_	     <= 1'b0;
			k8f9lz_optfi4vcf	     <= 1'b0;
			op9rx4p45h29r	     <= 1'b0;
		end
		else if (jfo4e1ypekb5lfzzx39_4ru0) begin
			erplkdk9eejnm26v2q9axu    <= 1'b0;
			a91q0mpju3lvvuyy	     <= tzfebftjmirx__sl5mroslq;
			sbn67m1e906fpvnin8pxq <= 1'b0;
			c9fbc2_3b0q24_wa9w84pk    <= 1'b0;
			u3x9iybnpf8suar92	     <= 1'b0;
			sb57m7q7jimdmg_	     <= 1'b0;
			k8f9lz_optfi4vcf	     <= 1'b0;
			op9rx4p45h29r	     <= 1'b0;
		end
		else if (ka6mrfj_02knc55k6) begin
			erplkdk9eejnm26v2q9axu    <= p60i1235jw07wggo07zuxm;
			a91q0mpju3lvvuyy	     <= c9jvr8hzwcs0svgzgj4x;
			sbn67m1e906fpvnin8pxq <= nkqcgp9gxttikxmttl77t7sx;
			c9fbc2_3b0q24_wa9w84pk    <= z1uojli46j34r_32meos9;
			u3x9iybnpf8suar92	     <= d5g9bjqnj4hlkaa8tl1v;
			sb57m7q7jimdmg_	     <= q1o9g4lcei7dy3z1;
			k8f9lz_optfi4vcf	     <= s93zuexjncoy1wmij4u;
			op9rx4p45h29r	     <= tljwcx5n4m9ruiltki;
		end
	end

	always @(posedge gf33atgy or negedge hfocw7va5_) begin
		if (!hfocw7va5_) begin
			om4i8b1g4ffpkkjkse91 <= 32'd0;
		end
		else if (!o59nl09azxaz) begin
			om4i8b1g4ffpkkjkse91 <= 32'd0;
		end
		else if (doaxea8vme8i1z) begin
			om4i8b1g4ffpkkjkse91 <= cf1p9na3s94mkxr663b;
		end
	end
	
	always @(posedge gf33atgy or negedge hfocw7va5_) begin
		if (!hfocw7va5_) begin
			sf14ab4y4pwg9uzf7ei <= 32'd0;
		end
		else if (!o59nl09azxaz) begin
			sf14ab4y4pwg9uzf7ei <= 32'd0;
		end
		else if (xuea1_k_eg81xsp7) begin
			sf14ab4y4pwg9uzf7ei <= b2kif3s0l5f10gxlqp;
		end
	end

	always @(posedge gf33atgy or negedge hfocw7va5_) begin
		if (!hfocw7va5_) begin
			at1z83ksz098eaaw45zorq <= 32'd0;
		end
		else if (!o59nl09azxaz) begin
			at1z83ksz098eaaw45zorq <= 32'd0;
		end
		else if (ub0do2eia4_zpjgutcd) begin
			at1z83ksz098eaaw45zorq <= chxwpklhgug7nuaerfmj;
		end
	end
	
	always @(posedge gf33atgy or negedge hfocw7va5_) begin
		if (!hfocw7va5_) begin
			pmxmx6g704kt9ffe_k3gsb4 <= 32'd0;
		end
		else if (!o59nl09azxaz) begin
			pmxmx6g704kt9ffe_k3gsb4 <= 32'd0;
		end
		else if (ooobnffsf8o6qo9i) begin
			pmxmx6g704kt9ffe_k3gsb4 <= vhvg6pli9i9rtyr0gpued;
		end
	end

	always @(posedge gf33atgy or negedge hfocw7va5_) begin
		if (!hfocw7va5_) begin
			cn8y8j2rziuq8l <= 16'd0;
		end
		else if (!o59nl09azxaz) begin
			cn8y8j2rziuq8l <= 16'd0;
		end
		else if (otd6qmzkpph) begin
			cn8y8j2rziuq8l <= z54sfjatc1sac9pfiv;
		end
	end

	always @(posedge gf33atgy or negedge hfocw7va5_) begin
		if (!hfocw7va5_) begin
			ln0owurz2hrjqyzt <= 32'd0;
		end
		else if (!o59nl09azxaz) begin
			ln0owurz2hrjqyzt <= 32'd0;
		end
		else if (wlhp1d9_0qsm5__) begin
			ln0owurz2hrjqyzt <= asuxi27dz56cq9qk1q6;
		end
	end
	
	always @(posedge gf33atgy or negedge hfocw7va5_) begin
		if (!hfocw7va5_) begin
			jy3u2zz45w3qt2o8ueas <= 32'd0;
		end
		else if (!o59nl09azxaz) begin
			jy3u2zz45w3qt2o8ueas <= 32'd0;
		end
		else if (zz9n5bfhur01yx) begin
			jy3u2zz45w3qt2o8ueas <= shq4l11_gkpyac;
		end
	end
	
	always @(posedge gf33atgy or negedge hfocw7va5_) begin
		if (!hfocw7va5_) begin
			riur0xm9vgi7prn <= 32'd0;
		end
		else if (!o59nl09azxaz) begin
			riur0xm9vgi7prn <= 32'd0;
		end
		else if (w2bzlpz5nmwdb2d) begin
			riur0xm9vgi7prn <= zaqsdqqsq29r81i;
		end
	end
	
	always @(posedge gf33atgy or negedge hfocw7va5_) begin
		if (!hfocw7va5_) begin
			g4n2d80tx347g5d <= 32'd0;
		end
		else if (!o59nl09azxaz) begin
			g4n2d80tx347g5d <= 32'd0;
		end
		else if (tdjiiekyziosyf) begin
			g4n2d80tx347g5d <= lbwqg4gjtgckn2f;
		end
	end
	
	assign alpkrgsdgm3z2_llqs9wc = od6u7rr1fxvo091a298 & erplkdk9eejnm26v2q9axu;
	assign h7bf8fgzcxv2nr5q_g4nygf5c = j0d0ajxf_i5ihg3yt95    & c9fbc2_3b0q24_wa9w84pk;
	assign xt_seq2pq4js8rmtsz = (gvbp1k6dl4r0o3hg6n | alpkrgsdgm3z2_llqs9wc | h7bf8fgzcxv2nr5q_g4nygf5c) & jlwst2h0gt_6sp4da7gy;
	assign idbkyxhyplh8ik16cau = nijvffj_k83iteeb61;
	assign gw5bpkb0gwli80bq  = xt_seq2pq4js8rmtsz | (~idbkyxhyplh8ik16cau & dlgkkhcodyhtm4ue);

	assign ssay1k38w94lso_ = dlgkkhcodyhtm4ue & (alpkrgsdgm3z2_llqs9wc | h7bf8fgzcxv2nr5q_g4nygf5c);
	assign q3jh_tep8g0mk7m2ohvp     = (ka6mrfj_02knc55k6 & ph7jz_7_o_welqv[22])  ? 1'b0 : 
					 ssay1k38w94lso_ ? 1'b1 :
							   shsgn99xfgm_falbwej9r;
	assign p60i1235jw07wggo07zuxm    = ph7jz_7_o_welqv[20];
	assign c9jvr8hzwcs0svgzgj4x	       = ph7jz_7_o_welqv[19:17];
	assign nkqcgp9gxttikxmttl77t7sx = ph7jz_7_o_welqv[16];
	assign z1uojli46j34r_32meos9    = ph7jz_7_o_welqv[15];

	assign wvyzyntlw4ro36s310tyw  = {ntt3vblrcouy6if54la, l36ob57itxhda2q, jij19fj8jksetx4, ivo3nt6en_d1s4fnn, msljxv405r4t1rbl};

	assign szmaji702081lti_h0qux = nwrntu_ns6js9tio & ~ph7jz_7_o_welqv[14:12];
	assign vcedcqevwspfk05rtor3 = nijvffj_k83iteeb61 & y98wkjik72p2pi;

	assign zzzclorwnw16vf8    = (a91q0mpju3lvvuyy == z68iccz0j602b2m9uekd7utr) &   y2bt8u7bruuxsctix[0];
	assign u5mjc2lh222oaobj    = (a91q0mpju3lvvuyy == tzfebftjmirx__sl5mroslq) & (|y2bt8u7bruuxsctix[1:0]);
	assign btob5wz940x35dypuh    = (a91q0mpju3lvvuyy == obhfbd2skwiz5h4ycuhz8qc) & (|y2bt8u7bruuxsctix[2:0]);
	assign hyqrpuxs_jhuma9ai4f9f = ~dnah6nc0fw8ts_1ltvjz & (zzzclorwnw16vf8 | u5mjc2lh222oaobj | btob5wz940x35dypuh);
	assign dnah6nc0fw8ts_1ltvjz = ~|((5'b00001 << a91q0mpju3lvvuyy) & wvyzyntlw4ro36s310tyw);
	assign xkda0fom0vel4oensw7 = hyqrpuxs_jhuma9ai4f9f | dnah6nc0fw8ts_1ltvjz;
	assign i4oiz2wl_m8q5y00l76bwi = hyqrpuxs_jhuma9ai4f9f & mtlruvvjhcvzf6;
	assign kp5ybypb04805jmkg3619oh3s8 = dnah6nc0fw8ts_1ltvjz & mtlruvvjhcvzf6;
	assign pnghshojyfxwjqjregrnf = nijvffj_k83iteeb61 | ka6mrfj_02knc55k6 | i4oiz2wl_m8q5y00l76bwi | kp5ybypb04805jmkg3619oh3s8;
	assign bjkw1ffrzjhax1g63pke	= ({3{ka6mrfj_02knc55k6       }} & szmaji702081lti_h0qux)
				| ({3{vcedcqevwspfk05rtor3       }} & 3'd2)
				| ({3{i4oiz2wl_m8q5y00l76bwi    }} & 3'd3)
				| ({3{kp5ybypb04805jmkg3619oh3s8}} & 3'd4);

	assign doaxea8vme8i1z = od6u7rr1fxvo091a298 | (sbn67m1e906fpvnin8pxq & nijvffj_k83iteeb61);
	assign xuea1_k_eg81xsp7 = fp20b2_fx9jb40co6__3 | (sbn67m1e906fpvnin8pxq & nijvffj_k83iteeb61);
	assign ub0do2eia4_zpjgutcd = iy011s14bjaestsjehfc | (sbn67m1e906fpvnin8pxq & nijvffj_k83iteeb61);
	assign ooobnffsf8o6qo9i = m9xf9uxglv4neo5ivk3 | (sbn67m1e906fpvnin8pxq & nijvffj_k83iteeb61);

	assign z8heidfnfd6oy8 = (32'd1 << a91q0mpju3lvvuyy);
	assign elm1vif4d_10b1_g8_2 = {e7wcd07jh85sk_hny6, bxlgqasel4nu6fjtmnt, zbawca6o200bvbpa1b6, y2bt8u7bruuxsctix};
	assign jd3bx8g5usv4rwh4  = elm1vif4d_10b1_g8_2 + {96'd0, z8heidfnfd6oy8};
	
	assign cf1p9na3s94mkxr663b = od6u7rr1fxvo091a298 ? ph7jz_7_o_welqv : jd3bx8g5usv4rwh4[31:0];
	assign b2kif3s0l5f10gxlqp = (x5jl_73d_gruzgtcqu >= 64) ? (fp20b2_fx9jb40co6__3 ? ph7jz_7_o_welqv : jd3bx8g5usv4rwh4[63:32] ) : 32'h0; 
	assign chxwpklhgug7nuaerfmj = (x5jl_73d_gruzgtcqu > 64 ) ? (iy011s14bjaestsjehfc ? ph7jz_7_o_welqv : jd3bx8g5usv4rwh4[95:64] ) : 32'h0; 
	assign vhvg6pli9i9rtyr0gpued = (x5jl_73d_gruzgtcqu > 64 ) ? (m9xf9uxglv4neo5ivk3 ? ph7jz_7_o_welqv : jd3bx8g5usv4rwh4[127:96]) : 32'h0;

	assign j3chbw93vus855iltfv4p = ph7jz_7_o_welqv;
	assign d6y6mbjwlwbautf9 = ph7jz_7_o_welqv;
	assign a2uofg5xxki0oe1xex155 = ph7jz_7_o_welqv;
	assign cjg6agdce9fgz9d1hl0v = ph7jz_7_o_welqv;

	assign d5g9bjqnj4hlkaa8tl1v  = (c9jvr8hzwcs0svgzgj4x == tzfebftjmirx__sl5mroslq) & l36ob57itxhda2q;
	assign q1o9g4lcei7dy3z1  = (c9jvr8hzwcs0svgzgj4x == obhfbd2skwiz5h4ycuhz8qc) & ntt3vblrcouy6if54la;
	assign s93zuexjncoy1wmij4u = (c9jvr8hzwcs0svgzgj4x <  tzfebftjmirx__sl5mroslq);
	assign otd6qmzkpph       = gvbp1k6dl4r0o3hg6n & k8f9lz_optfi4vcf;
	assign z54sfjatc1sac9pfiv  = a91q0mpju3lvvuyy[0] ? ph7jz_7_o_welqv[15:0] : {ph7jz_7_o_welqv[7:0], ph7jz_7_o_welqv[7:0]};
	assign tljwcx5n4m9ruiltki	 = ~(s93zuexjncoy1wmij4u | d5g9bjqnj4hlkaa8tl1v | q1o9g4lcei7dy3z1);

	assign vkb6t1zon4pxe = ({32{ k8f9lz_optfi4vcf}} & {cn8y8j2rziuq8l, cn8y8j2rziuq8l})
			    | ({32{~k8f9lz_optfi4vcf}} & ln0owurz2hrjqyzt);

	assign a0o2jippaa1o7rp5 = ({32{k8f9lz_optfi4vcf}} & {cn8y8j2rziuq8l, cn8y8j2rziuq8l})
			    | ({32{u3x9iybnpf8suar92}}  & ln0owurz2hrjqyzt)
			    | ({32{(op9rx4p45h29r | sb57m7q7jimdmg_)}} & jy3u2zz45w3qt2o8ueas);

	assign cguui3s6gp4x7 = ({32{k8f9lz_optfi4vcf}} & {cn8y8j2rziuq8l, cn8y8j2rziuq8l})
			    | ({32{op9rx4p45h29r}}	    & riur0xm9vgi7prn)
			    | ({32{(u3x9iybnpf8suar92 | sb57m7q7jimdmg_)}} & ln0owurz2hrjqyzt);

	assign rbaif3vx037msdnd = ({32{k8f9lz_optfi4vcf}} & {cn8y8j2rziuq8l, cn8y8j2rziuq8l})
			    | ({32{u3x9iybnpf8suar92}}  & ln0owurz2hrjqyzt)
			    | ({32{sb57m7q7jimdmg_}}  & jy3u2zz45w3qt2o8ueas)
			    | ({32{op9rx4p45h29r}}	    & g4n2d80tx347g5d);

	assign sb0_ui0s9qs02p22r_1[31:0]   = vkb6t1zon4pxe;
	assign sb0_ui0s9qs02p22r_1[63:32]  = a0o2jippaa1o7rp5;
    	assign sb0_ui0s9qs02p22r_1[95:64]  = cguui3s6gp4x7; 
	assign sb0_ui0s9qs02p22r_1[127:96] = rbaif3vx037msdnd;

	always @* begin
		case (a91q0mpju3lvvuyy[2:0])
		3'b000: 
			case ({(y2bt8u7bruuxsctix[3] & ntt3vblrcouy6if54la), (y2bt8u7bruuxsctix[2] & l36ob57itxhda2q), y2bt8u7bruuxsctix[1:0]}) 
				4'b0000: xwe5116fdnncgl5_idf0q = {24'd0, z1h6n4git1qfcautzkf7d[7:0]};
				4'b0001: xwe5116fdnncgl5_idf0q = {24'd0, z1h6n4git1qfcautzkf7d[15:8]};
				4'b0010: xwe5116fdnncgl5_idf0q = {24'd0, z1h6n4git1qfcautzkf7d[23:16]};
				4'b0011: xwe5116fdnncgl5_idf0q = {24'd0, z1h6n4git1qfcautzkf7d[31:24]};
				4'b0100: xwe5116fdnncgl5_idf0q = {24'd0, z1h6n4git1qfcautzkf7d[39:32]};
				4'b0101: xwe5116fdnncgl5_idf0q = {24'd0, z1h6n4git1qfcautzkf7d[47:40]};
				4'b0110: xwe5116fdnncgl5_idf0q = {24'd0, z1h6n4git1qfcautzkf7d[55:48]};
				4'b0111: xwe5116fdnncgl5_idf0q = {24'd0, z1h6n4git1qfcautzkf7d[63:56]};
				4'b1000: xwe5116fdnncgl5_idf0q = {24'd0, z1h6n4git1qfcautzkf7d[71:64]};
				4'b1001: xwe5116fdnncgl5_idf0q = {24'd0, z1h6n4git1qfcautzkf7d[79:72]};
				4'b1010: xwe5116fdnncgl5_idf0q = {24'd0, z1h6n4git1qfcautzkf7d[87:80]};
				4'b1011: xwe5116fdnncgl5_idf0q = {24'd0, z1h6n4git1qfcautzkf7d[95:88]};
				4'b1100: xwe5116fdnncgl5_idf0q = {24'd0, z1h6n4git1qfcautzkf7d[103:96]};
				4'b1101: xwe5116fdnncgl5_idf0q = {24'd0, z1h6n4git1qfcautzkf7d[111:104]};
				4'b1110: xwe5116fdnncgl5_idf0q = {24'd0, z1h6n4git1qfcautzkf7d[119:112]};
				4'b1111: xwe5116fdnncgl5_idf0q = {24'd0, z1h6n4git1qfcautzkf7d[127:120]};
				default: xwe5116fdnncgl5_idf0q = 32'dx;
			endcase
		3'b001: 
			case (y2bt8u7bruuxsctix[3:1]) 
				3'b000: xwe5116fdnncgl5_idf0q = {16'd0, z1h6n4git1qfcautzkf7d[15:0]};	
				3'b001: xwe5116fdnncgl5_idf0q = {16'd0, z1h6n4git1qfcautzkf7d[31:16]};	
				3'b010: xwe5116fdnncgl5_idf0q = {16'd0, z1h6n4git1qfcautzkf7d[47:32]};	
				3'b011: xwe5116fdnncgl5_idf0q = {16'd0, z1h6n4git1qfcautzkf7d[63:48]};	
				3'b100: xwe5116fdnncgl5_idf0q = {16'd0, z1h6n4git1qfcautzkf7d[79:64]};	
				3'b101: xwe5116fdnncgl5_idf0q = {16'd0, z1h6n4git1qfcautzkf7d[95:80]};	
				3'b110: xwe5116fdnncgl5_idf0q = {16'd0, z1h6n4git1qfcautzkf7d[111:96]};	
				3'b111: xwe5116fdnncgl5_idf0q = {16'd0, z1h6n4git1qfcautzkf7d[127:112]};	
				default: xwe5116fdnncgl5_idf0q = 32'dx;
			endcase
		3'b010:
			case (y2bt8u7bruuxsctix[3:2])
				2'b00: xwe5116fdnncgl5_idf0q = z1h6n4git1qfcautzkf7d[31:0];
				2'b01: xwe5116fdnncgl5_idf0q = z1h6n4git1qfcautzkf7d[63:32];
				2'b10: xwe5116fdnncgl5_idf0q = z1h6n4git1qfcautzkf7d[95:64];
				2'b11: xwe5116fdnncgl5_idf0q = z1h6n4git1qfcautzkf7d[127:96];
			endcase
		
		3'b011:	xwe5116fdnncgl5_idf0q = z1h6n4git1qfcautzkf7d[31:0];
		3'b100:	xwe5116fdnncgl5_idf0q = z1h6n4git1qfcautzkf7d[31:0];
		default: xwe5116fdnncgl5_idf0q = z1h6n4git1qfcautzkf7d[31:0];
		endcase
	end
	
	assign xoviomvc7o7y87p3yap = (a91q0mpju3lvvuyy[2:0] == 3'b011) ? z1h6n4git1qfcautzkf7d[63:32] : 32'h0;
	assign rfdqkys5p2ujup5_mm2n = z1h6n4git1qfcautzkf7d[95:64];
	assign owcemq5_leom8y6ncl = z1h6n4git1qfcautzkf7d[127:96];

	assign p6rade23wlwj8tphay = qdso0sntbt33twwh90;
	assign qrsc_8c1f0s50ogii = qdso0sntbt33twwh90 & l36ob57itxhda2q;
	assign hehn594ckxi95te8 = qdso0sntbt33twwh90 & ntt3vblrcouy6if54la;
	assign czya52zksuaqev = qdso0sntbt33twwh90 & ntt3vblrcouy6if54la;

	assign asuxi27dz56cq9qk1q6 = gvbp1k6dl4r0o3hg6n ? j3chbw93vus855iltfv4p : xwe5116fdnncgl5_idf0q;
	assign shq4l11_gkpyac = (x5jl_73d_gruzgtcqu >= 64) ? (kits5q7f_cnh6v1l ? d6y6mbjwlwbautf9 : xoviomvc7o7y87p3yap) : 32'h0;
	assign zaqsdqqsq29r81i = (x5jl_73d_gruzgtcqu > 64 ) ? (vzl0_w7ht4urni897h3 ? a2uofg5xxki0oe1xex155 : rfdqkys5p2ujup5_mm2n) : 32'h0;
	assign lbwqg4gjtgckn2f = (x5jl_73d_gruzgtcqu > 64 ) ? (ppt849kffgp8e6pv9j ? cjg6agdce9fgz9d1hl0v : owcemq5_leom8y6ncl) : 32'h0;
	
	assign wlhp1d9_0qsm5__ =  gvbp1k6dl4r0o3hg6n | p6rade23wlwj8tphay;
	assign zz9n5bfhur01yx = (kits5q7f_cnh6v1l | qrsc_8c1f0s50ogii) & l36ob57itxhda2q;
	assign w2bzlpz5nmwdb2d = (vzl0_w7ht4urni897h3 | hehn594ckxi95te8) & ntt3vblrcouy6if54la;
	assign tdjiiekyziosyf = (ppt849kffgp8e6pv9j | czya52zksuaqev) & ntt3vblrcouy6if54la;

	assign gsmp8y890cng = {xuzpr_ag_zzjjlhleh, 6'd0, shsgn99xfgm_falbwej9r, dlgkkhcodyhtm4ue, erplkdk9eejnm26v2q9axu, a91q0mpju3lvvuyy, 
			   sbn67m1e906fpvnin8pxq, c9fbc2_3b0q24_wa9w84pk, nwrntu_ns6js9tio, kz_vf5v7hkz3, ntt3vblrcouy6if54la, 
			   l36ob57itxhda2q, jij19fj8jksetx4, ivo3nt6en_d1s4fnn, msljxv405r4t1rbl};
	assign y2bt8u7bruuxsctix = om4i8b1g4ffpkkjkse91;
	assign zbawca6o200bvbpa1b6 = sf14ab4y4pwg9uzf7ei;
	assign bxlgqasel4nu6fjtmnt = at1z83ksz098eaaw45zorq;
	assign e7wcd07jh85sk_hny6 = pmxmx6g704kt9ffe_k3gsb4;
	assign oqevdjmfdhtvo    = ln0owurz2hrjqyzt;
	assign o12utn841wpwhrex    = jy3u2zz45w3qt2o8ueas;
	assign ayv5i_2icurn_    = riur0xm9vgi7prn;
	assign ue0zf04oji91y_44    = g4n2d80tx347g5d;



assign ai18gqgs_7ews5o     = nrxv3rneu2438;
assign ci1v3d4sfydbh_sz     = ai18gqgs_7ews5o & xgi_ovaieihs4f & !e_pz9vwnoa1r523;










ux607_gnrl_dfflr #(32) tos5s69zwu98ow_bdn8y (ci1v3d4sfydbh_sz, nd7gkqyz8zkdg3, tigza5anv0i48c7, gf33atgy, hfocw7va5_);

wire njhx5n_op0yb7gm_vyl      = (ehdeq25ha[8:2] == jcqkgadqjnp1br60kcm7);
wire pdzwfy9pk3b5svl6cvcj     = (ehdeq25ha[8:2] == wjwm0mmb8kdtc38hmvxcg7);
wire z9jm0ut6nbh6kyp1l96h      = (ehdeq25ha[8:2] == r9pqyndxl9ydaeube81umk);
wire esss55cpr6isvlpd56m43      = (ehdeq25ha[8:2] == dakqe9s6bwbckfsw4zlpj);
wire tamcjleq42fhwopgxdo3_o6_3 = (ehdeq25ha[8:2] == aon_4_u6h74hgk3ispa3if13);
wire o6q8tmuwwf_toj3mda    = (ehdeq25ha[8:2] == aufn2qiboj8l12dufk0p);
wire nyy07ivb1kfodzq3ymtp    = (ehdeq25ha[8:2] == xpf4_70tcyabeblxkt7aob2y);
wire y82a2i5o124hqncb1       = (ehdeq25ha[8:2] == bcei3m4eneqv0kswce_6);
wire nlnjr9n0_cb_jpwdj_iqz  = (ehdeq25ha[8:2] == rzuyw47p7ehj1uy43z4w9l63d3);
wire u2ry39tw1_30gq05v3z   = (ehdeq25ha[8:2] == yi9jeqslby_o_kzsjsm3);
wire mb267xvi0ttvdtsowy_w0l   = (ehdeq25ha[8:2] == wu726eflupgjm7hs9uonaad7p);
wire by5mxc0x6bct82k436d2c   = (ehdeq25ha[8:2] == js76iv7t9nvkn6yv_4661);
wire gs7zpu8n6wq0oaf9qjij3s   = (ehdeq25ha[8:2] == fufl25ug_h3jqm3k9o_gkyii);
wire yu1649mlxykb6         = (ehdeq25ha[8:2] == ggr6ql2zj7x40114w);
wire e5y49nph_ez39         = (ehdeq25ha[8:2] == tcnwfsqopcq2kj);
wire twj2grwj9ljye         = (ehdeq25ha[8:2] == ab_j1frhbffg57rc);
wire okdzf57tgwjr0         = (ehdeq25ha[8:2] == jim0ddiqnav_mr);
wire tm1jmyv1gu61hwhy         = (ehdeq25ha[8:2] == m0jpn5dn80dsf2q);
wire nr3mm5k5r0zhti8fbk         = (ehdeq25ha[8:2] == zxe9_q2s5fzxgu_k38);
wire njzi0kzl3_32u         = (ehdeq25ha[8:2] == va10rh7n02nkb6);
wire kicvef_8sd32wv6baw         = (ehdeq25ha[8:2] == dmgo2idd7_vdsdnnaq3);
wire qnk_0bdroh3yfx         = (ehdeq25ha[8:2] == jbtj7er6n1t919tqlx);
wire stmesantvywf91         = (ehdeq25ha[8:2] == qz57tyn0hruiw2xcq);
wire qd94c12p5f6493es4bq        = (ehdeq25ha[8:2] == kfpiwe2xk_8vve0);
wire e96rsuov2npbrazf        = (ehdeq25ha[8:2] == esrb21vaoahytvbimz);
wire ljo1ulblsd9ddlraw      = (ehdeq25ha[8:2] == u_cztegv7294f0w2ck);
wire i2btk5ij_tlwjioph      = (ehdeq25ha[8:2] == ew_k_8affyv8ltn2n9t);
wire k_my464a4gmk4ccq      = (ehdeq25ha[8:2] == c2pgc56ortybp6qk31tah2);
wire lsu7l9vbkzofaw7xlpy      = (ehdeq25ha[8:2] == vojasz8wlqnrlmd7irtxe);
wire saair51so3vezkkotv3n      = (ehdeq25ha[8:2] == bhmgs3vgnseqkofaq);
wire s5hnsat0f7wga6234bpk      = (ehdeq25ha[8:2] == v1p67sbkplioln574gw);
wire gvr6fi5eto8aaefh      = (ehdeq25ha[8:2] == s8hr7m7qhl3pqnt89tus);
wire roqlp4oc_oc4_bys64j      = (ehdeq25ha[8:2] == z6pqul13taj_bw4t8yli);
wire rd948sx674bdnyiua6xnv      = (ehdeq25ha[8:2] == hvhnim02z6srj83lugw);
wire c0mkbgblwyte0k_wb42e9      = (ehdeq25ha[8:2] == v7um53_ht6a2cwt6ubl2u5);
wire kfe_2l1ed6qbodnnu0w     = (ehdeq25ha[8:2] == usr_d4ztbwfqnw1ksw);
wire jdpddsjp6d4r5b_l4_sfhe     = (ehdeq25ha[8:2] == s8z4ks84p0yw2dqwwu);
wire q5ahcshwwj4hl16cgoh     = (ehdeq25ha[8:2] == fbu4pj38gfgemse5eu);
wire t5n9owyrabs62s34r     = (ehdeq25ha[8:2] == vf67ei0xuhdiywaae5mejm);
wire fh4fqeqkuzkj1_qzlus     = (ehdeq25ha[8:2] == p_0cn2roe14mgc29a_0h);
wire ey5b48q1n0kyjfw6dts     = (ehdeq25ha[8:2] == oo6atcmpor7odv_pblz40y);
wire uopzrn1k0tyyuuoag      = (ehdeq25ha[8:2] == klufzp92vwn000j_r);
wire y55hvs7x7vwyenxfmng      = (ehdeq25ha[8:2] == if4yqcjnanofw8tsvk);
wire si3qepcci4hpr          = (ehdeq25ha[8:2] == qnwyvxc9qyjqiu);
wire n8g90nmtwa8dus48jrry    = (ehdeq25ha[8:2] == co7pv8p2kbxe610a1fd6iz);
wire zz0m5gqmwt888fwts07z    = (ehdeq25ha[8:2] == jscy4q366gyq9lj13lo9r_t);
wire weyklv5yeeuu_lsyxr    = (ehdeq25ha[8:2] == gdv3d9wl61p6agakjyorlu6);
wire czniuh3upbvbrzr73j3bm    = (ehdeq25ha[8:2] == gv3onvtfu_6pjps2fsz57vdz);
wire d17lzosigos84bs       = (ehdeq25ha[8:2] == jebjru_ggwvrtiwo8i);
wire tc1tnx0yx12b2pt       = (ehdeq25ha[8:2] == gzcyq45ld9_ynnk5);
wire c8wek614e1cnw5cswnnb       = (ehdeq25ha[8:2] == lm2c1fdkx8du93b_9);
wire mvi6qplppvv_nabjnkz       = (ehdeq25ha[8:2] == g11_czp4uyqfn8ri);
wire p5mbtrcu683_lxf38      = (ehdeq25ha[8:2] == mibasbdgzaznbi2ob);

assign nd7gkqyz8zkdg3 =   ({32{njhx5n_op0yb7gm_vyl     }} & r65hrblk6cfz_)
                       | ({32{pdzwfy9pk3b5svl6cvcj    }} & q7xpkacoiqp__elsg)
                       | ({32{z9jm0ut6nbh6kyp1l96h     }} & tchrn3tov0okb6f)
                       | ({32{esss55cpr6isvlpd56m43     }} & y80_gmc7mbs2g68)
                       | ({32{tamcjleq42fhwopgxdo3_o6_3}} & s51p9m5pter6agwkfmi)
                       | ({32{o6q8tmuwwf_toj3mda   }} & lu2p7m5sdkbd)
                       | ({32{nyy07ivb1kfodzq3ymtp   }} & stcjaa1sbc18df8)
                       | ({32{y82a2i5o124hqncb1      }} & hq9truyassja3d8s)
                       | ({32{nlnjr9n0_cb_jpwdj_iqz }} & kg9c2fr3o4t1l2_udn)
                       | ({32{u2ry39tw1_30gq05v3z  }} & roo2isb7xjjd372j766)
                       | ({32{mb267xvi0ttvdtsowy_w0l  }} & osmjr77x4r43r658pa)
                       | ({32{by5mxc0x6bct82k436d2c  }} & h0s2y_7k2obvxraruu45)
                       | ({32{gs7zpu8n6wq0oaf9qjij3s  }} & rewvin436j1jc4w)
                       | ({32{yu1649mlxykb6        }} & ajymk4x2v3)
                       | ({32{e5y49nph_ez39        }} & mlyn8clead)
                       | ({32{twj2grwj9ljye        }} & g2544euz9jpuu9)
                       | ({32{okdzf57tgwjr0        }} & rw_eqfvro8)
                       | ({32{tm1jmyv1gu61hwhy        }} & 32'b0)
                       | ({32{nr3mm5k5r0zhti8fbk        }} & 32'b0)
                       | ({32{njzi0kzl3_32u        }} & 32'b0)
                       | ({32{kicvef_8sd32wv6baw        }} & 32'b0)
                       | ({32{qnk_0bdroh3yfx        }} & 32'b0)
                       | ({32{stmesantvywf91        }} & 32'b0)
                       | ({32{qd94c12p5f6493es4bq       }} & 32'b0)
                       | ({32{e96rsuov2npbrazf       }} & 32'b0)
                       | ({32{ljo1ulblsd9ddlraw     }} & dmi_progbuf0)
                       | ({32{i2btk5ij_tlwjioph     }} & i053jzqawhse)
                       | ({32{k_my464a4gmk4ccq     }} & tg3msrog_0bv)
                       | ({32{lsu7l9vbkzofaw7xlpy     }} & g30pvzblnaf83zh)
                       | ({32{saair51so3vezkkotv3n     }} & j2juyav34kkmuqd)
                       | ({32{s5hnsat0f7wga6234bpk     }} & watz9oqgogsyjeo)
                       | ({32{gvr6fi5eto8aaefh     }} & kriizvysvcfvd)
                       | ({32{roqlp4oc_oc4_bys64j     }} & l97zx3ot2wagshr9)
                       | ({32{rd948sx674bdnyiua6xnv     }} & heiy5swkajxipcai)
                       | ({32{c0mkbgblwyte0k_wb42e9     }} & etxdm_c986j2h)
                       | ({32{kfe_2l1ed6qbodnnu0w    }} & iw9ukx193kjidkn)
                       | ({32{jdpddsjp6d4r5b_l4_sfhe    }} & hwwlvkrpw_rd1)
                       | ({32{q5ahcshwwj4hl16cgoh    }} & b81eb_9kn7xgu725)
                       | ({32{t5n9owyrabs62s34r    }} & rj3ujsskxnsw3)
                       | ({32{fh4fqeqkuzkj1_qzlus    }} & fp511hjp_uccxk4)
                       | ({32{ey5b48q1n0kyjfw6dts    }} & dde_945nq4horxo)
                       | ({32{uopzrn1k0tyyuuoag     }} & rwyvi96_wuktwcs65)
                       | ({32{y55hvs7x7vwyenxfmng     }} & dr8lpark3fykgiqvl)
                       | ({32{si3qepcci4hpr         }} & gsmp8y890cng)
                       | ({32{n8g90nmtwa8dus48jrry   }} & y2bt8u7bruuxsctix)
                       | ({32{zz0m5gqmwt888fwts07z   }} & zbawca6o200bvbpa1b6)
                       | ({32{weyklv5yeeuu_lsyxr   }} & bxlgqasel4nu6fjtmnt)
                       | ({32{czniuh3upbvbrzr73j3bm   }} & e7wcd07jh85sk_hny6)
                       | ({32{d17lzosigos84bs      }} & oqevdjmfdhtvo)
                       | ({32{tc1tnx0yx12b2pt      }} & o12utn841wpwhrex)
                       | ({32{c8wek614e1cnw5cswnnb      }} & ayv5i_2icurn_)
                       | ({32{mvi6qplppvv_nabjnkz      }} & ue0zf04oji91y_44)
                       | ({32{p5mbtrcu683_lxf38     }} & ws9kutgi4r0wui1)
                       ;





























































genvar pa3ohjp_zdvw6w;
generate
if (s_hrmp88w3m_7k29y == "uci2r") begin : yyhuj6991mc9ku920f1o
	wire                    vwylbr7u3j4mi5iqit_5h_x;
	wire [8:0]              ury740k32four;
	wire [2:0]              de3t2irquwko3atn67;
	wire                    rw6e7cvsxd4f40mig;

	wire [vmw6vavuv7md5-1:0]   f4jcdkmf2du_knygwtq08v;
	wire [vmw6vavuv7md5-1:0]   a04o140evqlw3mw;
	wire                    pkxkm53fkzwapatf0zsb_qhni;

	wire                    t2xogqackphhs2nom6;

	wire                    exjl1aq54hbbcjxy4n;
	wire                    s1m0779f4lb7mgzcrse70;
	wire                    evn1_dsee0mpk_woecwb4bm9tqp;

	ux607_gnrl_dffrs #(1) k35zllomktxb39ntbtd1 (s1m0779f4lb7mgzcrse70, exjl1aq54hbbcjxy4n, gf33atgy, hfocw7va5_);










	ux607_gnrl_dfflr #(9) gbcf66r8rybgjten (n2vqwxz4b7yahnp, evqksuwcgvwotl[8:0], ury740k32four, gf33atgy, hfocw7va5_);
	ux607_gnrl_dfflr #(3) tf4h8to_whij26jt (n2vqwxz4b7yahnp, qbiibzbu0j5xu, de3t2irquwko3atn67, gf33atgy, hfocw7va5_);
	ux607_gnrl_dfflr #(1) x_k2uio2in6wf0a4 (n2vqwxz4b7yahnp, ohod7vxvej8qwj, rw6e7cvsxd4f40mig, gf33atgy, hfocw7va5_);
	ux607_gnrl_dfflr #(1) fguxo23l3mygy3ziwvrnm3iw (n2vqwxz4b7yahnp, u06qbygttylwtj63blcgmn, vwylbr7u3j4mi5iqit_5h_x, gf33atgy, hfocw7va5_);
















	ux607_gnrl_dfflr #(vmw6vavuv7md5) uqrss2gp72jc6u67tz43t9 (xjstumkuxktuwybrt70f09d, f4jcdkmf2du_knygwtq08v, a04o140evqlw3mw, gf33atgy, hfocw7va5_);









	assign t2xogqackphhs2nom6 = tk2pf9erp83 & p9_huoh6oy1jai[1] & n2vqwxz4b7yahnp;
	assign u06qbygttylwtj63blcgmn = t2xogqackphhs2nom6 & ohod7vxvej8qwj;
	assign d65omgobthbz58hr4v6c8vye = vwylbr7u3j4mi5iqit_5h_x;
	assign oq56n5j5gd3i2trf1n23 = (de3t2irquwko3atn67 == 3'h3) | ((de3t2irquwko3atn67 < 3'h3) &  yygzyugpvajoy2ito[2]);
	assign rgr3u9u7smu2_9zb3od6u4  = (de3t2irquwko3atn67 == 3'h3) | ((de3t2irquwko3atn67 < 3'h3) & ~yygzyugpvajoy2ito[2]);
    assign qxlm3tn20surby98      = (de3t2irquwko3atn67 == 3'h3) ? 8'hff :
                                  (de3t2irquwko3atn67 == 3'h2) ? (8'h0f << {yygzyugpvajoy2ito[2:2],2'b0}) : 
                                  (de3t2irquwko3atn67 == 3'h1) ? (8'h03 << {yygzyugpvajoy2ito[2:1],1'b0}) : 
                                  (de3t2irquwko3atn67 == 3'h0) ? (8'h01 << {yygzyugpvajoy2ito[2:0]}) : 
                                  8'h00; 
    assign dk5qlcqv4hzz3221yncmzmjpc  = {{8{qxlm3tn20surby98[3]}}, {8{qxlm3tn20surby98[2]}}, {8{qxlm3tn20surby98[1]}}, {8{qxlm3tn20surby98[0]}}};
    assign p009emefkiuou558jih1od36 = {{8{qxlm3tn20surby98[7]}}, {8{qxlm3tn20surby98[6]}}, {8{qxlm3tn20surby98[5]}}, {8{qxlm3tn20surby98[4]}}};

	assign evn1_dsee0mpk_woecwb4bm9tqp = (p9_huoh6oy1jai[1]==1'b0);
	assign s1m0779f4lb7mgzcrse70    =  evn1_dsee0mpk_woecwb4bm9tqp | ~u06qbygttylwtj63blcgmn;

	assign v5jhtjwnqklb6oje85 = exjl1aq54hbbcjxy4n;

	assign pkxkm53fkzwapatf0zsb_qhni = (vmw6vavuv7md5 == 32) & bf2jgqu2qq_lbyd[2];

	for (pa3ohjp_zdvw6w = 0; pa3ohjp_zdvw6w<vmw6vavuv7md5; pa3ohjp_zdvw6w=pa3ohjp_zdvw6w+32) begin: n4hjx3i2sc2r9o7o6vb31
		if (pa3ohjp_zdvw6w == 32) begin: w9atag6bcur3xgztz805bo0bq
			assign f4jcdkmf2du_knygwtq08v[(pa3ohjp_zdvw6w+31):pa3ohjp_zdvw6w] = vq_q6kxvnkkqf2[(pa3ohjp_zdvw6w+31):pa3ohjp_zdvw6w];
		end
		else begin: u5cnv54tg6toie36e1ly
			assign f4jcdkmf2du_knygwtq08v[(pa3ohjp_zdvw6w+31):pa3ohjp_zdvw6w] = pkxkm53fkzwapatf0zsb_qhni ? vq_q6kxvnkkqf2[63:32] : vq_q6kxvnkkqf2[31:0];
		end
	end

	assign xjstumkuxktuwybrt70f09d = t2xogqackphhs2nom6 & !ohod7vxvej8qwj; 




	assign uqi13ctmbgrce5j9 = ury740k32four[8:2];
	assign yygzyugpvajoy2ito  = ury740k32four[2:0];
	assign qvpivcc8d7j57jlwl[63:32] = fa9ntbvuu_3cuqr5[(vmw6vavuv7md5-1):(vmw6vavuv7md5-32)];
	assign qvpivcc8d7j57jlwl[31:0]  = fa9ntbvuu_3cuqr5[31:0];
	assign bf2jgqu2qq_lbyd = evqksuwcgvwotl[8:2];

	assign coiuburq3cf  = a04o140evqlw3mw;
	assign lzl17_6p6y91nh = g9rl8dm8yn;

end
endgenerate

generate
if (s_hrmp88w3m_7k29y != "uci2r") begin : fffsg0y3i9lkmt83lceang4zc8r36
	assign coiuburq3cf    = {vmw6vavuv7md5{1'b0}};
	assign v5jhtjwnqklb6oje85 = 1'b1;
	assign lzl17_6p6y91nh     = 2'd0;
end
endgenerate




























































































































































































































generate
if (vmw6vavuv7md5 == 64) begin: yzxke6lq129prnqog4xmrb2ujh76iqu
	assign jqecsbcna9xks4236v7y = d65omgobthbz58hr4v6c8vye & ( uqi13ctmbgrce5j9             == gixg8zsazjmz1x_brls) &  rgr3u9u7smu2_9zb3od6u4;
	assign bg6j3mh0cbpsnjsw8 = d65omgobthbz58hr4v6c8vye & ({uqi13ctmbgrce5j9[8:3], 1'b0} == gixg8zsazjmz1x_brls) & (uqi13ctmbgrce5j9[2] | oq56n5j5gd3i2trf1n23);
	assign g3ss6oez6hga6h4sc = d65omgobthbz58hr4v6c8vye & ( uqi13ctmbgrce5j9             == hzzi56ur3pc3ozd55y9) &  rgr3u9u7smu2_9zb3od6u4;
	assign bpf8y70t6yfklo_g8w2vz = d65omgobthbz58hr4v6c8vye & ({uqi13ctmbgrce5j9[8:3], 1'b0} == hzzi56ur3pc3ozd55y9) & (uqi13ctmbgrce5j9[2] | oq56n5j5gd3i2trf1n23);
	assign wmao806lq98cxpivg = d65omgobthbz58hr4v6c8vye & ( uqi13ctmbgrce5j9             == zvqpf_dzodsppyt2sy_) &  rgr3u9u7smu2_9zb3od6u4;
	assign d65wnf88ntcgv6j5aqzdd = d65omgobthbz58hr4v6c8vye & ({uqi13ctmbgrce5j9[8:3], 1'b0} == zvqpf_dzodsppyt2sy_) & (uqi13ctmbgrce5j9[2] | oq56n5j5gd3i2trf1n23);
	assign zyrzsibwzfi9i9wbbf = d65omgobthbz58hr4v6c8vye & ( uqi13ctmbgrce5j9             == t9kao6jz00ceq9met6r) &  rgr3u9u7smu2_9zb3od6u4;
	assign lu303j9kh0__1tuhdc3wn1 = d65omgobthbz58hr4v6c8vye & ({uqi13ctmbgrce5j9[8:3], 1'b0} == t9kao6jz00ceq9met6r) & (uqi13ctmbgrce5j9[2] | oq56n5j5gd3i2trf1n23);
	assign meq51ng31supqk_vkxuh = d65omgobthbz58hr4v6c8vye & ( uqi13ctmbgrce5j9             == vdoigs60y4azen6d3tcs) &  rgr3u9u7smu2_9zb3od6u4;
	assign vhake2p_2q859v6b79w9bt = d65omgobthbz58hr4v6c8vye & ({uqi13ctmbgrce5j9[8:3], 1'b0} == vdoigs60y4azen6d3tcs) & (uqi13ctmbgrce5j9[2] | oq56n5j5gd3i2trf1n23);
	assign nimnckhhiicxl3my3yxx = d65omgobthbz58hr4v6c8vye & ( uqi13ctmbgrce5j9             == ytd01d3exnn7ehvy8m4gi) &  rgr3u9u7smu2_9zb3od6u4;
	assign yi1sq51qvk1rehte9p8_ = d65omgobthbz58hr4v6c8vye & ({uqi13ctmbgrce5j9[8:3], 1'b0} == ytd01d3exnn7ehvy8m4gi) & (uqi13ctmbgrce5j9[2] | oq56n5j5gd3i2trf1n23);
	assign lapvh12sh70dkfu0lnktk5 = d65omgobthbz58hr4v6c8vye & ( uqi13ctmbgrce5j9             == fpg_uog8qlop0ciegpq) &  rgr3u9u7smu2_9zb3od6u4;
	assign ts8jeswko5lfbpmtqe = d65omgobthbz58hr4v6c8vye & ({uqi13ctmbgrce5j9[8:3], 1'b0} == fpg_uog8qlop0ciegpq) & (uqi13ctmbgrce5j9[2] | oq56n5j5gd3i2trf1n23);
	assign yjole_26w_x6maqonk = d65omgobthbz58hr4v6c8vye & ( uqi13ctmbgrce5j9             == xvf_oe_m8metbe7ln0og8m7x) &  rgr3u9u7smu2_9zb3od6u4;
	assign oj1yq4vf080z10xcce = d65omgobthbz58hr4v6c8vye & ({uqi13ctmbgrce5j9[8:3], 1'b0} == xvf_oe_m8metbe7ln0og8m7x) & (uqi13ctmbgrce5j9[2] | oq56n5j5gd3i2trf1n23);

	assign tf1byd_17w8d_ypae4v      = d65omgobthbz58hr4v6c8vye & ( uqi13ctmbgrce5j9             == qj3a7cq7w0bujncuh) &  rgr3u9u7smu2_9zb3od6u4;
	assign p1yn5zqqxm8yw8ox      = d65omgobthbz58hr4v6c8vye & ({uqi13ctmbgrce5j9[8:3], 1'b0} == qj3a7cq7w0bujncuh) & (uqi13ctmbgrce5j9[2] | oq56n5j5gd3i2trf1n23);
	assign h3e4drj186x9hakap0e      = d65omgobthbz58hr4v6c8vye & ( uqi13ctmbgrce5j9             == uqw9t32734czfnllj) &  rgr3u9u7smu2_9zb3od6u4;
	assign uev0sc6o93o2rcvvy3p      = d65omgobthbz58hr4v6c8vye & ({uqi13ctmbgrce5j9[8:3], 1'b0} == uqw9t32734czfnllj) & (uqi13ctmbgrce5j9[2] | oq56n5j5gd3i2trf1n23);

	assign lxnlpqnqclk48r5        = d65omgobthbz58hr4v6c8vye & ( uqi13ctmbgrce5j9             == yhf4gk3fjs1g0c7vmxpfv) &  rgr3u9u7smu2_9zb3od6u4;
	assign w6r9d62ex8olvrj0zfd7     = d65omgobthbz58hr4v6c8vye & ({uqi13ctmbgrce5j9[8:3], 1'b0} == yhf4gk3fjs1g0c7vmxpfv) & (uqi13ctmbgrce5j9[2] | oq56n5j5gd3i2trf1n23);
	assign qcv2n1t0m8gvo5cto     = d65omgobthbz58hr4v6c8vye & ( uqi13ctmbgrce5j9             == km0i5rel2kki7saovbnju)  &  rgr3u9u7smu2_9zb3od6u4;
	assign w3f078jh09ukd9z_24  = d65omgobthbz58hr4v6c8vye & ({uqi13ctmbgrce5j9[8:3], 1'b0} == km0i5rel2kki7saovbnju)  & (uqi13ctmbgrce5j9[2] | oq56n5j5gd3i2trf1n23);
end
else begin: zb7_oq7lgaq9wofvdznuz_cwj5v1bi
	assign jqecsbcna9xks4236v7y = d65omgobthbz58hr4v6c8vye & (uqi13ctmbgrce5j9 == gixg8zsazjmz1x_brls);
	assign bg6j3mh0cbpsnjsw8 = d65omgobthbz58hr4v6c8vye & (uqi13ctmbgrce5j9 == ufd6dm208s7jyarlo651ta);
	assign g3ss6oez6hga6h4sc = d65omgobthbz58hr4v6c8vye & (uqi13ctmbgrce5j9 == hzzi56ur3pc3ozd55y9);
	assign bpf8y70t6yfklo_g8w2vz = d65omgobthbz58hr4v6c8vye & (uqi13ctmbgrce5j9 == grybk8armp6w_25n2athlf);
	assign wmao806lq98cxpivg = d65omgobthbz58hr4v6c8vye & (uqi13ctmbgrce5j9 == zvqpf_dzodsppyt2sy_);
	assign d65wnf88ntcgv6j5aqzdd = d65omgobthbz58hr4v6c8vye & (uqi13ctmbgrce5j9 == kknbs_o3gqn0uzb6uxydb);
	assign zyrzsibwzfi9i9wbbf = d65omgobthbz58hr4v6c8vye & (uqi13ctmbgrce5j9 == t9kao6jz00ceq9met6r);
	assign lu303j9kh0__1tuhdc3wn1 = d65omgobthbz58hr4v6c8vye & (uqi13ctmbgrce5j9 == bk1_dfc2yewnml9b67xq);
	assign meq51ng31supqk_vkxuh = d65omgobthbz58hr4v6c8vye & (uqi13ctmbgrce5j9 == vdoigs60y4azen6d3tcs);
	assign vhake2p_2q859v6b79w9bt = d65omgobthbz58hr4v6c8vye & (uqi13ctmbgrce5j9 == ui48c9q5f2turr4gak47g);
	assign nimnckhhiicxl3my3yxx = d65omgobthbz58hr4v6c8vye & (uqi13ctmbgrce5j9 == ytd01d3exnn7ehvy8m4gi);
	assign yi1sq51qvk1rehte9p8_ = d65omgobthbz58hr4v6c8vye & (uqi13ctmbgrce5j9 == ohbi7syrfghop_1ei_7_v);
	assign lapvh12sh70dkfu0lnktk5 = d65omgobthbz58hr4v6c8vye & (uqi13ctmbgrce5j9 == fpg_uog8qlop0ciegpq);
	assign ts8jeswko5lfbpmtqe = d65omgobthbz58hr4v6c8vye & (uqi13ctmbgrce5j9 == c1lm4w95w1htl5nau42b);
	assign yjole_26w_x6maqonk = d65omgobthbz58hr4v6c8vye & (uqi13ctmbgrce5j9 == xvf_oe_m8metbe7ln0og8m7x);
	assign oj1yq4vf080z10xcce = d65omgobthbz58hr4v6c8vye & (uqi13ctmbgrce5j9 == ougtjwdhlld141546ol2ns);
	assign tf1byd_17w8d_ypae4v      = d65omgobthbz58hr4v6c8vye & (uqi13ctmbgrce5j9 == qj3a7cq7w0bujncuh);
	assign p1yn5zqqxm8yw8ox      = d65omgobthbz58hr4v6c8vye & (uqi13ctmbgrce5j9 == mt_9sbagghbuv5a);
	assign h3e4drj186x9hakap0e      = d65omgobthbz58hr4v6c8vye & (uqi13ctmbgrce5j9 == uqw9t32734czfnllj);
	assign uev0sc6o93o2rcvvy3p      = d65omgobthbz58hr4v6c8vye & (uqi13ctmbgrce5j9 == uvrkvxlxjv2ua24u);

	assign lxnlpqnqclk48r5        = d65omgobthbz58hr4v6c8vye & (uqi13ctmbgrce5j9 == yhf4gk3fjs1g0c7vmxpfv);
	assign w6r9d62ex8olvrj0zfd7     = d65omgobthbz58hr4v6c8vye & (uqi13ctmbgrce5j9 == mjsby4jqzutfz8ukh);
	assign qcv2n1t0m8gvo5cto     = d65omgobthbz58hr4v6c8vye & (uqi13ctmbgrce5j9 == km0i5rel2kki7saovbnju);
	assign w3f078jh09ukd9z_24  = d65omgobthbz58hr4v6c8vye & (uqi13ctmbgrce5j9 == yupij6i5uojje3u3bdgiy5);
end
endgenerate

wire [8:2] one397_ei0wvyl7e_5g = {bf2jgqu2qq_lbyd[8:3], 1'b0};

wire bb4evvtg5eod3fkgigx = (one397_ei0wvyl7e_5g == 7'h00);
wire xfh7zgd9w_ez4m7up = (one397_ei0wvyl7e_5g == 7'h02);
wire nm8bss06ohbt8qpok = (one397_ei0wvyl7e_5g == 7'h04);
wire l8rkjonggse89vris = (one397_ei0wvyl7e_5g == 7'h06);
wire ifh76_omx3yzqvqv_j = (one397_ei0wvyl7e_5g == 7'h08);
wire we7a_th88lk00j217 = (one397_ei0wvyl7e_5g == 7'h0a);
wire toooc9o5colgs1cnsqi = (one397_ei0wvyl7e_5g == 7'h0c);
wire nfe4x8_fatbsb522h = (one397_ei0wvyl7e_5g == 7'h0e);
wire zsd21fkw32zihz2xarc = (one397_ei0wvyl7e_5g == 7'h10);
wire jshcvmq4i2twqdie3ok2f = (one397_ei0wvyl7e_5g == 7'h12);
wire r663njeuww2be0tt = (one397_ei0wvyl7e_5g == 7'h14);
wire qhj4d758djx251ihkm = (one397_ei0wvyl7e_5g == 7'h16);
wire qw_eo0l6gnm8gpk94fwo = (one397_ei0wvyl7e_5g == 7'h18);
wire lk408jz062l1e2ie1lt = (one397_ei0wvyl7e_5g == gixg8zsazjmz1x_brls);
wire rtsnojpnpehvr61v07_d = (one397_ei0wvyl7e_5g == hzzi56ur3pc3ozd55y9);
wire fkqijso58i8nrdjr5kcly2 = (one397_ei0wvyl7e_5g == zvqpf_dzodsppyt2sy_);
wire axuore29wnf_udfwp = (one397_ei0wvyl7e_5g == t9kao6jz00ceq9met6r);
wire tijjwwswb9jyn3wq46ij = (one397_ei0wvyl7e_5g == vdoigs60y4azen6d3tcs);
wire oae86p6pcj7nv_53y3ue5z = (one397_ei0wvyl7e_5g == ytd01d3exnn7ehvy8m4gi);
wire zasnxkh7t801ov3lin = (one397_ei0wvyl7e_5g == fpg_uog8qlop0ciegpq);
wire x6h02b98rq3k7924u81qjp = (one397_ei0wvyl7e_5g == xvf_oe_m8metbe7ln0og8m7x);
wire xoi_kj5168_egj = (one397_ei0wvyl7e_5g == qj3a7cq7w0bujncuh);
wire b4rc33kqy5mijs8p1v = (one397_ei0wvyl7e_5g == uqw9t32734czfnllj);
wire j387i87httbd98jnq = (one397_ei0wvyl7e_5g == u62d_7aeq5rs779p);
wire u3rudfcix48n7apz = (one397_ei0wvyl7e_5g == qrwi8l03c71sin9ruze);
wire tqzsu534uj856bij_f = (one397_ei0wvyl7e_5g == h7qm4gdchgihbuedfbw);
wire e_8734x9adxf7j5o = (one397_ei0wvyl7e_5g == df826w0tr0ujt7no0z_0);
wire bizbwc363x3xq2xt5qhc = (one397_ei0wvyl7e_5g == o0b3kayk7gpelof4ct);
wire xmb04mdkvnstbd24w1 = (one397_ei0wvyl7e_5g == e5e_dbyenxum0n6fkma5);
wire zgrtnewjdxmg8h9wej = (one397_ei0wvyl7e_5g == yhf4gk3fjs1g0c7vmxpfv);
wire y97uguuo2l560m4_ha  = (one397_ei0wvyl7e_5g == km0i5rel2kki7saovbnju);

assign vq_q6kxvnkkqf2 =   ({64{bb4evvtg5eod3fkgigx  }} & {32'h10802223, 32'h0140006f})
                    | ({64{xfh7zgd9w_ez4m7up  }} & {32'h10801483, 32'h0ff0000f})
                    | ({64{nm8bss06ohbt8qpok  }} & {32'h7b241073, 32'h00c0006f})
                    | ({64{l8rkjonggse89vris  }} & {32'h10801483, 32'h7b349073})
                    | ({64{ifh76_omx3yzqvqv_j  }} & {32'h10802623, 32'hf1402473})
                    | ({64{we7a_th88lk00j217  }} & {32'h4004c493, 32'h00848a63})
                    | ({64{toooc9o5colgs1cnsqi  }} & {32'h10801483, 32'h02940463})
                    | ({64{nfe4x8_fatbsb522h  }} & {32'h10802423, 32'hff1ff06f})
                    | ({64{zsd21fkw32zihz2xarc  }} & {32'h7b202473, 32'h7b3024f3})
                    | ({64{jshcvmq4i2twqdie3ok2f  }} & {32'h7b3024f3, 32'h08000067})
                    | ({64{r663njeuww2be0tt  }} & {32'h00100073, 32'h7b202473})
                    | ({64{qhj4d758djx251ihkm  }} & {32'h7b3024f3, 32'h10802023})
                    | ({64{qw_eo0l6gnm8gpk94fwo  }} & {32'h7b200073, 32'h7b202473})
                    | ({64{lk408jz062l1e2ie1lt }} & {i053jzqawhse, dmi_progbuf0})
                    | ({64{rtsnojpnpehvr61v07_d }} & {g30pvzblnaf83zh, tg3msrog_0bv})
                    | ({64{fkqijso58i8nrdjr5kcly2 }} & {watz9oqgogsyjeo, j2juyav34kkmuqd})
                    | ({64{axuore29wnf_udfwp }} & {l97zx3ot2wagshr9, kriizvysvcfvd})
                    | ({64{tijjwwswb9jyn3wq46ij }} & {etxdm_c986j2h, heiy5swkajxipcai})
                    | ({64{oae86p6pcj7nv_53y3ue5z}} & {hwwlvkrpw_rd1, iw9ukx193kjidkn})
                    | ({64{zasnxkh7t801ov3lin}} & {rj3ujsskxnsw3, b81eb_9kn7xgu725})
                    | ({64{x6h02b98rq3k7924u81qjp}} & {dde_945nq4horxo, fp511hjp_uccxk4})
                    | ({64{xoi_kj5168_egj    }} & {mlyn8clead, ajymk4x2v3})
                    | ({64{b4rc33kqy5mijs8p1v    }} & {rw_eqfvro8, g2544euz9jpuu9})
                    | ({64{j387i87httbd98jnq    }} & 64'h0)
                    | ({64{u3rudfcix48n7apz    }} & 64'h0)
                    | ({64{tqzsu534uj856bij_f  }} & {mrse_xs0n5gn, jdv2ldkc9_q})
                    | ({64{e_8734x9adxf7j5o  }} & {tp7gcrgcgawl, qqgwfuykbb})
                    | ({64{bizbwc363x3xq2xt5qhc  }} & {xwh383jprd, atyzruk57fe})
                    | ({64{xmb04mdkvnstbd24w1  }} & {swxb1euiqwukq, fsq3dvu1_f7r})
                    | ({64{zgrtnewjdxmg8h9wej  }} & {hn_zgnzhnj4hl,    c3b14wbbm2jilagqe})
                    | ({64{y97uguuo2l560m4_ha   }} & {us8z6yxgvplahq18t, l5hh1f8jbhu6})
                    ;





















































endmodule














module ncec8v13ika897y(
input         qzy,
input         pg862o7b3cdc,
input         um8zsjyxn_4p,
input         joqaqv6v,
output        xu5bs,
output [31:0] cuf0p,
output        qhme7drv,
input         phl7z55l1,
input  [31:0] difhtk01a    
);

wire		jn738r_c;
wire		hi8t5vgnna3na;
wire		tz94thcv;

wire		pq1s3od1sc;
wire		vhig79ew7;
wire		dib6tggz;

wire	[31:0]	ap6cjp481mtgeyt_9p;

ux607_gnrl_dffr #(1) tfwrp3895o3ot (jn738r_c , xu5bs, qzy, pg862o7b3cdc);








ux607_gnrl_dffr #(1) js21q1cflrs5wh (pq1s3od1sc , qhme7drv, qzy, pg862o7b3cdc);









assign jn738r_c = ~tz94thcv & (xu5bs | hi8t5vgnna3na);
assign pq1s3od1sc = ~dib6tggz & (qhme7drv | vhig79ew7);

assign hi8t5vgnna3na = joqaqv6v & (um8zsjyxn_4p | phl7z55l1);
assign tz94thcv = ~joqaqv6v;

assign vhig79ew7 = joqaqv6v & (~um8zsjyxn_4p);
assign dib6tggz = um8zsjyxn_4p | phl7z55l1;

assign ap6cjp481mtgeyt_9p[31:27] = 5'd0;
assign ap6cjp481mtgeyt_9p[26:24] = 3'd0;	
assign ap6cjp481mtgeyt_9p[23]    = 1'd0;
assign ap6cjp481mtgeyt_9p[22]    = 1'b1;	
assign ap6cjp481mtgeyt_9p[21:20] = 2'd0;
assign ap6cjp481mtgeyt_9p[19]    = 1'b0;
assign ap6cjp481mtgeyt_9p[18]    = 1'b0;
assign ap6cjp481mtgeyt_9p[17]    = 1'b0;
assign ap6cjp481mtgeyt_9p[16]    = 1'b0;
assign ap6cjp481mtgeyt_9p[15]    = 1'b0;
assign ap6cjp481mtgeyt_9p[14]    = 1'b0;
assign ap6cjp481mtgeyt_9p[13]    = 1'b1;
assign ap6cjp481mtgeyt_9p[12]    = 1'b1;
assign ap6cjp481mtgeyt_9p[11]    = 1'b0;
assign ap6cjp481mtgeyt_9p[10]    = 1'b0;
assign ap6cjp481mtgeyt_9p[9]     = 1'b0;
assign ap6cjp481mtgeyt_9p[8]     = 1'b0;
assign ap6cjp481mtgeyt_9p[7]     = 1'b1;
assign ap6cjp481mtgeyt_9p[6]     = 1'b0;
assign ap6cjp481mtgeyt_9p[5]     = 1'b1;
assign ap6cjp481mtgeyt_9p[4]     = 1'b0;
assign ap6cjp481mtgeyt_9p[3:0]   = 4'd2;

assign cuf0p = um8zsjyxn_4p ? ap6cjp481mtgeyt_9p : difhtk01a;

endmodule

module q33ia3_pmvsc # (
  parameter  y76n53l844691b1v  = 41
) (
input			            yez0ldac23i95,

output			            qfuuzymrquo,
input			            jfyllx,
input			            a9c,
output			            hmb,
input			            qzy,
input			            pg862o7b3cdc, 
input	[31:0]			    nfgz90l9a50bvdr,
input			            eb1xb06elqtqv245,
output			            dz84q2c8wa_v,
output  [y76n53l844691b1v-1:0]  r6zq8pddzmjao10p,
output			            cnaq1epzg8_uh2_y

);







localparam n9yhq4z46fy7_o491 = 3'd7;






   

localparam k5v5zz_p2b48hhtfsr = 4'b0000;
localparam q7bqbah2usdmzt0v    = 4'b1000;
localparam m9_idq9vt6ir3j_ucem   = 4'b1001;
localparam deoi3trzar	    = 4'b1010;
localparam pggc0cu5	    = 4'b1011;
localparam k0y9xo3k	    = 4'b1100;
localparam k_ebupxqey9g	    = 4'b1101;
localparam g9g2m13jkgu	    = 4'b1110;
localparam j8_6nemvrado	    = 4'b1111;
localparam ldn1j7ttrydiakuf   = 4'b0001;
localparam rp8uncbkv39o_u	    = 4'b0010;
localparam rvsgjp6cm7d2p	    = 4'b0011;
localparam hkiu05mm	    = 4'b0100;
localparam hih_rr5jye5	    = 4'b0101;
localparam jk7ki709pean7	    = 4'b0110;
localparam du7oerk3swn0s	    = 4'b0111;


localparam p5f71s           = 5'b00001;
localparam p_kv_y71a1x      = 5'b10000;
localparam iv7cfne_mkoxqz       = 5'b10001;


localparam   ao_qx1lk8t0mh5c          = 2'b00;
localparam   y2w_s42cf6_94         = 2'b01;
localparam   ie_kg74b_wufbrz        = 2'b10;
localparam   yz80u836w74tl          = 2'b11;

localparam of7vq7lffln = 5;




wire		qx3du41e;
wire		d31sibjyhx;


wire	jiltdny0au7_4ma0a14n88;


wire		ouf9n20noqrgw0cl;
wire		hy3ssb0zcsakb9h9s;
wire		aqfm0yxtra_9qki;
wire		w2uioxuq9kxu4;
wire		wf57r5hv9zgqc505l9;
wire		q204koub4syelcu;
wire		gbu2s3m4x_4bbs;
wire		iyyavdsatgkm21;
wire		q1e810vt89gzw0x;
wire		a0s5ia70wr9st4ruflr;
wire		pd1xdq251ywp0kojb;
wire		xfuzomljx1xp6f0xb4v0;
wire		s5oumjp58ndkgo2z7;
wire		t6m113r1yr3tc_6;
wire		oigzvnd1fxm5xb9a3sa;
wire		icfxza6_s0kgnn23;
wire		nwi13ynijsfyitdvvrfq;
wire		zdp0xepiesnd;
wire		b67j8wcwc26z_;
wire		x3pffrhwfg281_iw;
wire		kgd3r_wvdl4fywjsz;
wire	[3:0]	ijtg0efa_3w7;
wire	[3:0]	jhrrb5snx_zr1lj;


wire	[of7vq7lffln-1:0]	g_7eo3;


wire	[y76n53l844691b1v-1:0]	nyrdflhfrhp9fdx;
wire	[y76n53l844691b1v-1:0]	ngqu4v_2wegw16sjfhvl8u16;
wire	[y76n53l844691b1v-1:0] 	k2nifhq80zylhc613z9;


wire [32-1:0] q0obiasp6da3z_e = 32'h0420122a;
wire [32-1:0] vbp39vpr6b_tjkwt = 32'h14202111;
wire [32-1:0] m_bbjo_s8fpy = 32'h04204732;
wire [32-1:0] cvumdg7g9d63o4z = (q0obiasp6da3z_e + vbp39vpr6b_tjkwt + m_bbjo_s8fpy);



wire	[1:0]	an70chyimnkpc_ycsv;
wire	[31:0]	hg2_y;
wire	[3:0]	jyyerz8ufyhz10bo6;
wire	[5:0]	zvgwfsmq_elob;
wire	[2:0]	xw9dw8yuofq_;
wire		adj3mps_9e9vv70bpkt;
wire		mlvg73lh2lunbboj;


wire	[y76n53l844691b1v-1:0]	bdo;
wire				r3we6y3bdqf4x8f;







wire	ss5woob0z0u;
wire	zs6djxr1;


wire	m0u036ta1g6rm;

wire	ud59eel;
wire	d0eh90t;


assign	ud59eel           = jfyllx; 
assign	d0eh90t           = a9c;
assign	m0u036ta1g6rm    = ouf9n20noqrgw0cl;



assign jiltdny0au7_4ma0a14n88 = d31sibjyhx | ~adj3mps_9e9vv70bpkt;

ux607_gnrl_dffr #(1) vnxpcbb8hhjztzgjf477 (jiltdny0au7_4ma0a14n88 , cnaq1epzg8_uh2_y, qzy, pg862o7b3cdc);













assign	d31sibjyhx = (ijtg0efa_3w7 == k5v5zz_p2b48hhtfsr);
ux607_gnrl_dffr #(1) iuxw4pvt696cfjknv (d31sibjyhx , qx3du41e, qzy, pg862o7b3cdc);













wire	p2_6ejdc_qawt = 1'b1;



ux607_gnrl_dfflr #(4)    qtcmiqx9l1mepp9psze  (p2_6ejdc_qawt, ijtg0efa_3w7, jhrrb5snx_zr1lj, qzy, pg862o7b3cdc);










wire bzmsmzc40xrurpnkifimn921 = hy3ssb0zcsakb9h9s;
wire [3:0] ujl72zvct4m2af2dlz = d0eh90t ? k5v5zz_p2b48hhtfsr : q7bqbah2usdmzt0v;

wire xprjy_e24o5n0zcfpcab1p4g = aqfm0yxtra_9qki;
wire [3:0] px6si32877tixdxz = d0eh90t ? m9_idq9vt6ir3j_ucem : q7bqbah2usdmzt0v; 

wire d2wn1xhq44jcdlmrg1d7 = w2uioxuq9kxu4;
wire [3:0] qyzck31yt1us32nk8ib = d0eh90t ? ldn1j7ttrydiakuf : deoi3trzar;

wire dkjrfbjo6r1zxe236kjru8 = wf57r5hv9zgqc505l9; 
wire [3:0] z__1boafts5pehkv_39va = d0eh90t ? k0y9xo3k : pggc0cu5; 

wire omdiml50jg8k9y2xeypshc = q204koub4syelcu;
wire [3:0] gg9sku7hdv_ht445wwet = d0eh90t ? k0y9xo3k : pggc0cu5;

wire d35a3ragdhx517vaeqsez = gbu2s3m4x_4bbs;
wire [3:0] kl4mked9y1w6b505eu = d0eh90t ? j8_6nemvrado : k_ebupxqey9g;

wire ar03m56wiq89td0dgj8kxr = iyyavdsatgkm21;
wire [3:0] siiabq74px_m0u_gn = d0eh90t ? g9g2m13jkgu : k_ebupxqey9g;

wire ssuanuhh73z01n36r8dxvb5 = q1e810vt89gzw0x;
wire [3:0] mk_hdyhc9u97tae3n = d0eh90t ? j8_6nemvrado : pggc0cu5;

wire yv5ywwk6v9__ri7w1bn0v4 = a0s5ia70wr9st4ruflr;
wire [3:0] wzj0zqv6izuhyltlpt = d0eh90t ? m9_idq9vt6ir3j_ucem : q7bqbah2usdmzt0v;

wire w8dg_yh9gz71_vslexw__6s = pd1xdq251ywp0kojb;
wire [3:0] t7iytxkd4eu5i9glng = d0eh90t ? k5v5zz_p2b48hhtfsr : rp8uncbkv39o_u;

wire emqfqtshmgj68j4bgyurd5r = xfuzomljx1xp6f0xb4v0;
wire [3:0] w3l5ft83z_gf53z80ou = d0eh90t ? hkiu05mm : rvsgjp6cm7d2p;

wire kz7oj7s16osk0e2mw_r1l = s5oumjp58ndkgo2z7;
wire [3:0] juo6_0pc7sds477xk4cw = d0eh90t ? hkiu05mm : rvsgjp6cm7d2p;

wire pvapzco3ytmy6la9px1y0oj1 = t6m113r1yr3tc_6;
wire [3:0] w4glerywys9wrtz = d0eh90t ? du7oerk3swn0s : hih_rr5jye5;

wire n7oxbq162fw64v0uhhuy3 = oigzvnd1fxm5xb9a3sa;
wire [3:0] b6ranqf911o_dpje = d0eh90t ? jk7ki709pean7 : hih_rr5jye5;

wire gw1wvk9xes0_gg9u4vqw = icfxza6_s0kgnn23;
wire [3:0] xptnajk36gzykajb3x4 = d0eh90t ? du7oerk3swn0s : rvsgjp6cm7d2p;

wire z2k_vvjg6e5hgmlygsao0x1w4w = nwi13ynijsfyitdvvrfq;
wire [3:0] gco1088cc7vo7x64_sl_ = d0eh90t ? m9_idq9vt6ir3j_ucem : q7bqbah2usdmzt0v;

assign ijtg0efa_3w7 =   ({4{bzmsmzc40xrurpnkifimn921   }} & ujl72zvct4m2af2dlz  )
                    | ({4{xprjy_e24o5n0zcfpcab1p4g  }} & px6si32877tixdxz )
                    | ({4{d2wn1xhq44jcdlmrg1d7    }} & qyzck31yt1us32nk8ib )
                    | ({4{dkjrfbjo6r1zxe236kjru8 }} & z__1boafts5pehkv_39va)
                    | ({4{omdiml50jg8k9y2xeypshc   }} & gg9sku7hdv_ht445wwet  )
                    | ({4{d35a3ragdhx517vaeqsez   }} & kl4mked9y1w6b505eu  )
                    | ({4{ar03m56wiq89td0dgj8kxr   }} & siiabq74px_m0u_gn  )
                    | ({4{ssuanuhh73z01n36r8dxvb5   }} & mk_hdyhc9u97tae3n  )
                    | ({4{yv5ywwk6v9__ri7w1bn0v4  }} & wzj0zqv6izuhyltlpt )
                    | ({4{w8dg_yh9gz71_vslexw__6s    }} & t7iytxkd4eu5i9glng   )
                    | ({4{emqfqtshmgj68j4bgyurd5r }} & w3l5ft83z_gf53z80ou)
                    | ({4{kz7oj7s16osk0e2mw_r1l   }} & juo6_0pc7sds477xk4cw  )
                    | ({4{pvapzco3ytmy6la9px1y0oj1   }} & w4glerywys9wrtz  )
                    | ({4{n7oxbq162fw64v0uhhuy3   }} & b6ranqf911o_dpje  )
                    | ({4{gw1wvk9xes0_gg9u4vqw   }} & xptnajk36gzykajb3x4  )
                    | ({4{z2k_vvjg6e5hgmlygsao0x1w4w  }} & gco1088cc7vo7x64_sl_ )
                    ;


















































































































assign	hy3ssb0zcsakb9h9s   = (jhrrb5snx_zr1lj == k5v5zz_p2b48hhtfsr);
assign	aqfm0yxtra_9qki  = (jhrrb5snx_zr1lj == q7bqbah2usdmzt0v);
assign	w2uioxuq9kxu4    = (jhrrb5snx_zr1lj == m9_idq9vt6ir3j_ucem);
assign	wf57r5hv9zgqc505l9 = (jhrrb5snx_zr1lj == deoi3trzar);
assign	q204koub4syelcu   = (jhrrb5snx_zr1lj == pggc0cu5);
assign	gbu2s3m4x_4bbs   = (jhrrb5snx_zr1lj == k0y9xo3k);
assign	iyyavdsatgkm21   = (jhrrb5snx_zr1lj == k_ebupxqey9g);
assign	q1e810vt89gzw0x   = (jhrrb5snx_zr1lj == g9g2m13jkgu);
assign	a0s5ia70wr9st4ruflr  = (jhrrb5snx_zr1lj == j8_6nemvrado);
assign	pd1xdq251ywp0kojb    = (jhrrb5snx_zr1lj == ldn1j7ttrydiakuf);
assign	xfuzomljx1xp6f0xb4v0 = (jhrrb5snx_zr1lj == rp8uncbkv39o_u);
assign	s5oumjp58ndkgo2z7   = (jhrrb5snx_zr1lj == rvsgjp6cm7d2p);
assign	t6m113r1yr3tc_6   = (jhrrb5snx_zr1lj == hkiu05mm);
assign	oigzvnd1fxm5xb9a3sa   = (jhrrb5snx_zr1lj == hih_rr5jye5);
assign	icfxza6_s0kgnn23   = (jhrrb5snx_zr1lj == jk7ki709pean7);
assign	nwi13ynijsfyitdvvrfq  = (jhrrb5snx_zr1lj == du7oerk3swn0s);
assign	ouf9n20noqrgw0cl = s5oumjp58ndkgo2z7 | q204koub4syelcu;


assign	zdp0xepiesnd      = ~b67j8wcwc26z_ & ~x3pffrhwfg281_iw & ~kgd3r_wvdl4fywjsz;
assign	b67j8wcwc26z_      = (g_7eo3 == p5f71s);
assign	x3pffrhwfg281_iw = (g_7eo3 == p_kv_y71a1x);
assign	kgd3r_wvdl4fywjsz  = (g_7eo3 == iv7cfne_mkoxqz);




wire	th101msyhr;
wire	ldzsjja7fyfsy0;
wire	lo33ttlpctxw0a;
wire	t7ed0l1xd_drpr1;
wire	jo5pvzs7on7djkpi6;

assign	ldzsjja7fyfsy0 = adj3mps_9e9vv70bpkt & (dz84q2c8wa_v | eb1xb06elqtqv245);
assign	lo33ttlpctxw0a = dz84q2c8wa_v & ~eb1xb06elqtqv245;
assign	t7ed0l1xd_drpr1 = ldzsjja7fyfsy0 | lo33ttlpctxw0a;
assign	jo5pvzs7on7djkpi6 = ldzsjja7fyfsy0 | ~lo33ttlpctxw0a;

ux607_gnrl_dfflr #(1)    hgmp7oei9zzkg4l  (t7ed0l1xd_drpr1, jo5pvzs7on7djkpi6, th101msyhr, qzy, pg862o7b3cdc);

















wire			    eat208xsui1ex1qb4nk2;
wire	[y76n53l844691b1v-1:0]  z0rfk3n9yggh6;

wire			    ah88342gb82;
wire			    li9_0v4r1roodxg;
wire			    sdpph5f6eyty;
wire			    lmk6qw86c_trtqtn;

assign	lmk6qw86c_trtqtn	    = ~(dz84q2c8wa_v | (eb1xb06elqtqv245 & ~th101msyhr));
assign	ah88342gb82	    = lmk6qw86c_trtqtn & kgd3r_wvdl4fywjsz & (bdo[1:0] == y2w_s42cf6_94) & ~r3we6y3bdqf4x8f;
assign	li9_0v4r1roodxg	    = lmk6qw86c_trtqtn & kgd3r_wvdl4fywjsz & (bdo[1:0] == ie_kg74b_wufbrz) & ~r3we6y3bdqf4x8f;
assign	sdpph5f6eyty		    = (~lmk6qw86c_trtqtn | r3we6y3bdqf4x8f) & kgd3r_wvdl4fywjsz;

assign	z0rfk3n9yggh6           = xfuzomljx1xp6f0xb4v0 ? {{(y76n53l844691b1v-of7vq7lffln){1'b0}}, g_7eo3} : 
			      ({{(y76n53l844691b1v-32){1'b0}}, ({32{b67j8wcwc26z_}} & cvumdg7g9d63o4z)} |
			      {{(y76n53l844691b1v-32){1'b0}}, ({32{x3pffrhwfg281_iw}} & hg2_y)} |
			      ({bdo[y76n53l844691b1v-1:2], 2'd0} & {y76n53l844691b1v{li9_0v4r1roodxg}}) |			
			      ({bdo[y76n53l844691b1v-1:34], nfgz90l9a50bvdr, 2'd0} & {y76n53l844691b1v{ah88342gb82}}) |	
			      ({bdo[y76n53l844691b1v-1:34], 32'd0, 2'd3} & {y76n53l844691b1v{sdpph5f6eyty}}));		
assign	eat208xsui1ex1qb4nk2 = (wf57r5hv9zgqc505l9 & (b67j8wcwc26z_ | x3pffrhwfg281_iw | kgd3r_wvdl4fywjsz)) | 
			      (xfuzomljx1xp6f0xb4v0);
assign	ngqu4v_2wegw16sjfhvl8u16 = s5oumjp58ndkgo2z7 ? {{(y76n53l844691b1v-of7vq7lffln){1'b0}}, ud59eel, nyrdflhfrhp9fdx[of7vq7lffln-1:1]} :
			      kgd3r_wvdl4fywjsz  ? {ud59eel, nyrdflhfrhp9fdx[y76n53l844691b1v-1:1]} : {{(y76n53l844691b1v-32){1'b0}}, ud59eel, nyrdflhfrhp9fdx[31:1]};


wire			    seu7vveakh79_3d2s9;
wire			    xw2cia3gyj30jny6vux;
wire			    g2u91orsoykttd5i7be;
wire	[y76n53l844691b1v-1:0]  u1m9njupmdjbo7u1nn2;

assign 	k2nifhq80zylhc613z9    = eat208xsui1ex1qb4nk2 ? z0rfk3n9yggh6 : ngqu4v_2wegw16sjfhvl8u16;

assign	xw2cia3gyj30jny6vux   = m0u036ta1g6rm | wf57r5hv9zgqc505l9 | xfuzomljx1xp6f0xb4v0;
assign	g2u91orsoykttd5i7be   = qx3du41e;
assign	seu7vveakh79_3d2s9   = xw2cia3gyj30jny6vux | g2u91orsoykttd5i7be;
assign	u1m9njupmdjbo7u1nn2   = g2u91orsoykttd5i7be ? {(y76n53l844691b1v){1'b0}} : k2nifhq80zylhc613z9;

ux607_gnrl_dfflr #(y76n53l844691b1v)    aw3nv3m2k50wwbr53sn83  (seu7vveakh79_3d2s9, u1m9njupmdjbo7u1nn2, nyrdflhfrhp9fdx, qzy, pg862o7b3cdc);
















wire			    a9hfqa1as24qh5;
wire			    dylpfh33_6mn6c;
wire			    t37rnx7dfpy1zb;
wire	[of7vq7lffln-1:0]       gmrtsran3wkg;

assign	t37rnx7dfpy1zb          = qx3du41e;
assign	dylpfh33_6mn6c          = nwi13ynijsfyitdvvrfq;
assign	a9hfqa1as24qh5          = t37rnx7dfpy1zb | dylpfh33_6mn6c;
assign	gmrtsran3wkg          = t37rnx7dfpy1zb ? p5f71s : nyrdflhfrhp9fdx[of7vq7lffln-1:0];

ux607_gnrl_dfflrs #(1)          kjo9p9xtccxrq6y0ccj_6ob  (a9hfqa1as24qh5, gmrtsran3wkg[0], g_7eo3[0], qzy, pg862o7b3cdc);
ux607_gnrl_dfflr #(of7vq7lffln-1)  sz8sr1_ajhe8bc8_h36nl  (a9hfqa1as24qh5, gmrtsran3wkg[of7vq7lffln-1:1], g_7eo3[of7vq7lffln-1:1], qzy, pg862o7b3cdc);
















wire       zz4mpum5bmdhwt5y8;
wire       jv6ihvjdc9gwi15d_by;
wire       l5mgrwufzhk6xo1fa_;
wire [1:0] ivkgly9zoa6f7apmxx8;

assign	adj3mps_9e9vv70bpkt = x3pffrhwfg281_iw & a0s5ia70wr9st4ruflr & nyrdflhfrhp9fdx[17];
assign	mlvg73lh2lunbboj     = x3pffrhwfg281_iw & a0s5ia70wr9st4ruflr & nyrdflhfrhp9fdx[16];
assign	xw9dw8yuofq_	   = n9yhq4z46fy7_o491; 
assign	zvgwfsmq_elob	   = 6'd7; 	 
assign	jyyerz8ufyhz10bo6	   = 4'd1; 	 

assign	jv6ihvjdc9gwi15d_by  = wf57r5hv9zgqc505l9 & kgd3r_wvdl4fywjsz & ~lmk6qw86c_trtqtn;
assign	zz4mpum5bmdhwt5y8  = mlvg73lh2lunbboj | qx3du41e | adj3mps_9e9vv70bpkt;
assign	l5mgrwufzhk6xo1fa_  = zz4mpum5bmdhwt5y8 | jv6ihvjdc9gwi15d_by;
assign	ivkgly9zoa6f7apmxx8  = zz4mpum5bmdhwt5y8 ? 2'd0 : 2'd3;

ux607_gnrl_dfflr #(2)    ihappz7fuqgp6sw3kgclp7k  (l5mgrwufzhk6xo1fa_, ivkgly9zoa6f7apmxx8, an70chyimnkpc_ycsv, qzy, pg862o7b3cdc);















assign	hg2_y   	   = {14'b0,         1'b0,     1'b0, 1'b0, xw9dw8yuofq_, an70chyimnkpc_ycsv, zvgwfsmq_elob, jyyerz8ufyhz10bo6};




wire	r208ti6km3izaay;
wire	kruczij_kjpfkhpv;
wire	abllynrv084744fo;
wire	w638h4o265g3xnltts1;
wire	m77yzqe;

assign	r3we6y3bdqf4x8f  = (an70chyimnkpc_ycsv == 2'd3);
assign	m77yzqe 	        = ^nyrdflhfrhp9fdx[1:0];
assign	r208ti6km3izaay = a0s5ia70wr9st4ruflr & kgd3r_wvdl4fywjsz & m77yzqe & ~r3we6y3bdqf4x8f;
assign	kruczij_kjpfkhpv = (eb1xb06elqtqv245 & ~th101msyhr) | qx3du41e | adj3mps_9e9vv70bpkt;
assign	abllynrv084744fo = r208ti6km3izaay | kruczij_kjpfkhpv;
assign	w638h4o265g3xnltts1 = r208ti6km3izaay & ~kruczij_kjpfkhpv;

ux607_gnrl_dfflr #(1)    kj6wrffgpvah2juf8xvq  (abllynrv084744fo, w638h4o265g3xnltts1, dz84q2c8wa_v, qzy, pg862o7b3cdc);



















wire                    vg61w67yle;
wire                    sthjqdv6;
wire                    o17mbenhrh;
wire [y76n53l844691b1v-1:0] ze_bmycz30r;


assign	vg61w67yle  = a0s5ia70wr9st4ruflr & kgd3r_wvdl4fywjsz & ~r3we6y3bdqf4x8f;
assign	sthjqdv6  = qx3du41e;
assign	o17mbenhrh  = vg61w67yle | sthjqdv6;
assign	ze_bmycz30r  = sthjqdv6 ? {(y76n53l844691b1v){1'b0}} : nyrdflhfrhp9fdx;

ux607_gnrl_dfflr #(y76n53l844691b1v)    uomi9ff2j_dwk  (o17mbenhrh, ze_bmycz30r, bdo, qzy, pg862o7b3cdc);

assign	r6zq8pddzmjao10p   = bdo;
















wire	zp182g43v2qfa;
wire	z846jnlyhsxivt;
wire	nbpz9svc6xx;
wire	h8lm37rc3x3ulm;

assign	zs6djxr1     = (q204koub4syelcu & (zdp0xepiesnd ? ss5woob0z0u : nyrdflhfrhp9fdx[0])) |
		     (s5oumjp58ndkgo2z7 & nyrdflhfrhp9fdx[0]);
assign	zp182g43v2qfa = wf57r5hv9zgqc505l9 | qx3du41e;
assign	z846jnlyhsxivt = q204koub4syelcu & m0u036ta1g6rm;
assign	nbpz9svc6xx = zp182g43v2qfa | z846jnlyhsxivt;
assign	h8lm37rc3x3ulm = zp182g43v2qfa ? 1'b0 : ud59eel;

ux607_gnrl_dfflr #(1)    x7z87ig6j8ktc7rj  (nbpz9svc6xx, h8lm37rc3x3ulm, ss5woob0z0u, qzy, pg862o7b3cdc);













wire b9t1k = yez0ldac23i95 ? qzy : ~qzy;

wire	i5rm_q4wsax;
wire	m9tn_yqgft;
wire	ok4a_dz;
wire	acg8gzrvvs;

assign	i5rm_q4wsax = m0u036ta1g6rm;
assign	m9tn_yqgft = qx3du41e;
assign	ok4a_dz = i5rm_q4wsax | m9tn_yqgft;
assign	acg8gzrvvs = m9tn_yqgft ? 1'b0 : zs6djxr1;

ux607_gnrl_dfflr #(1)    pycv3eusvuho  (ok4a_dz, acg8gzrvvs, hmb, b9t1k, pg862o7b3cdc);

wire	il8i63py563r2krvq = i5rm_q4wsax;
wire	c14x9l0rt72yr9l = m9tn_yqgft;
wire	w15waqniluhh1gn9 = ok4a_dz;
wire	dke45gymk_y1r8sbr = il8i63py563r2krvq & ~c14x9l0rt72yr9l;

ux607_gnrl_dfflr #(1)    oqaayi70y_agzdv5x  (w15waqniluhh1gn9, dke45gymk_y1r8sbr, qfuuzymrquo, b9t1k, pg862o7b3cdc);



















endmodule



module d6pt7ab0 (
input              um8zsjyxn_4p,
input              sqvy97shfxgalqcq,

output             qfuuzymrquo,    
input              uecloq2rb,    
input              dfnv8e05y_xxox4kof,
input              na29rv9xyz_vn,
input              yez0ldac23i95 ,
input              qzy,           
input              a9c,           
input              jfyllx,          
output             hmb,         
output             a02zzbowpjn06h, 
output             lr4pmtw0e3sm7,   
input              bmm03who3rv,            
input              obvunz7,
input              d5gddvhozc,      
output             gtvu1jhq,      
output       [1:0] lpv3w7_jux0x5,    
output      [31:0] v0ppt_lszz,     
output       [2:0] naonfp5kwul39,     
output       [2:0] tfljpdijxf,    
output       [3:0] c98a8jw632g1,     
output      [31:0] j8tyg8pg_v_hj12,    
output             iw4viufqn3,    
input       [31:0] eplm38kc000z,    
input              m82k9gnjrw,    
output             hj3v8ja2n1snk, 
input              liu_rgb4nf      
);

localparam vv3o1dwe8bt1m3k = 32;
localparam b4ff6gp7ae52l = 7;
localparam opmj43kpf6ptzium   = 2;
localparam y76n53l844691b1v = vv3o1dwe8bt1m3k + b4ff6gp7ae52l + opmj43kpf6ptzium;

wire                           hhflrj5pivf;

wire                           pqoqazegmgqaxyrvv;
wire                    [31:0] w4l6em1v0os9uky;
wire                           cnaq1epzg8_uh2_y;
wire        [y76n53l844691b1v-1:0] nmmjpe9w4mnr;
wire                           vhi8lz75vjbjjyjdn5ee;
wire                           m13tjzrbil5w1qrfszwu;
wire                           sxlpd0g_kavoy2igabp;

wire                           z89ho_0fnb0d857lwtdrl5e;
wire                           e7b6a043i5yg2edz5v_j8;
wire                    [31:0] amrnb4vy1vg9zdg6va1gy;


assign a02zzbowpjn06h = ( sxlpd0g_kavoy2igabp | pqoqazegmgqaxyrvv);
















wire anf7yeobyty6du66cjemb = yez0ldac23i95 ? na29rv9xyz_vn : cnaq1epzg8_uh2_y;

ux607_gnrl_dffr #(1) fazreuhl4pcgo73t77 (1'b1 , hhflrj5pivf, obvunz7, anf7yeobyty6du66cjemb);








wire hqmnbsdg9xwl1sq6grx8;

ncec8v13ika897y ncec8v13ika897y(
         .qzy          (qzy                    ),
         .pg862o7b3cdc    (dfnv8e05y_xxox4kof          ),
         .um8zsjyxn_4p    (hqmnbsdg9xwl1sq6grx8      ),
         .joqaqv6v         (z89ho_0fnb0d857lwtdrl5e    ),
         .xu5bs         (e7b6a043i5yg2edz5v_j8    ),
         .cuf0p        (amrnb4vy1vg9zdg6va1gy     ),
         .qhme7drv         (vhi8lz75vjbjjyjdn5ee        ),
         .phl7z55l1         (m13tjzrbil5w1qrfszwu        ),
         .difhtk01a        (w4l6em1v0os9uky         )
);

q33ia3_pmvsc q33ia3_pmvsc (
    .yez0ldac23i95(yez0ldac23i95),

	.qfuuzymrquo    (qfuuzymrquo     ), 
	.jfyllx           (jfyllx            ), 
	.a9c           (a9c            ), 
	.hmb           (hmb            ), 
	.qzy           (qzy            ), 
	.pg862o7b3cdc     (dfnv8e05y_xxox4kof  ),
    .nfgz90l9a50bvdr(amrnb4vy1vg9zdg6va1gy ), 
    .eb1xb06elqtqv245   (e7b6a043i5yg2edz5v_j8),
    .dz84q2c8wa_v   (z89ho_0fnb0d857lwtdrl5e),
	.r6zq8pddzmjao10p  (nmmjpe9w4mnr   ), 
	.cnaq1epzg8_uh2_y(cnaq1epzg8_uh2_y ) 
); 

wire c5ihnefsy8pg2r5q8cvmfk = sxlpd0g_kavoy2igabp & (~um8zsjyxn_4p);

u_j2imkw7hy7 u_j2imkw7hy7 (
    
	.yg8hetdkahah       (sqvy97shfxgalqcq ), 
	.w4l6em1v0os9uky(w4l6em1v0os9uky  ), 
	.lb2ioj3kfjgks   (pqoqazegmgqaxyrvv), 
	.kvdg06d7vo7wv_n   (c5ihnefsy8pg2r5q8cvmfk), 
	.nmmjpe9w4mnr  (nmmjpe9w4mnr    ), 
	.wivo          (d5gddvhozc        ), 
	.zy4t8o4ibj         (liu_rgb4nf       ), 
	.oyn5mkpu        (m82k9gnjrw      ), 
	.y7ftxl        (eplm38kc000z      ), 
	.n1xcixngo_e     (hj3v8ja2n1snk   ), 
	.rw9vqyx         (v0ppt_lszz       ), 
	.mhayix        (lpv3w7_jux0x5      ), 
	.ad5i86r        (iw4viufqn3      ), 
	.tihusk1         (naonfp5kwul39       ), 
	.abdy0h        (tfljpdijxf      ), 
	.awm5ntb_         (c98a8jw632g1       ), 
	.t6tpgz13_m        (j8tyg8pg_v_hj12      ), 
	.l4pt3          (gtvu1jhq        )  
); 

u7uyomlq26a_3s81cs bsyhozfdzho1zycgnhwn0uc6 (
	.j0ln_h     (dfnv8e05y_xxox4kof       ), 
	.p2fq1i8       (qzy                 ), 
	.pg17e0     (pqoqazegmgqaxyrvv    ), 
	.qqk5yk     (m13tjzrbil5w1qrfszwu     ), 
	.khfri3vm7  (                    ), 
	.x7bl2zxqiftsf  (                    ), 
	.kgg1udim46o  (                    )  
);

u7uyomlq26a_3s81cs rvpvlj2mh5rc2esrssk5w25pxse1qs8wus (
	.j0ln_h     (dfnv8e05y_xxox4kof       ), 
	.p2fq1i8       (qzy                 ),
	.pg17e0     (um8zsjyxn_4p           ),
	.qqk5yk     (hqmnbsdg9xwl1sq6grx8   ),
	.khfri3vm7  (                    ),
	.x7bl2zxqiftsf  (                    ),
	.kgg1udim46o  (                    ) 
); 

u7uyomlq26a_3s81cs x3u6nf50yxkyvadpx7ryo47 (
	.j0ln_h     (na29rv9xyz_vn       ), 

	.p2fq1i8       (bmm03who3rv            ), 
	.pg17e0     (vhi8lz75vjbjjyjdn5ee     ), 
	.qqk5yk     (sxlpd0g_kavoy2igabp    ), 
	.khfri3vm7  (                    ), 
	.x7bl2zxqiftsf  (                    ), 
	.kgg1udim46o  (                    ) 
);

u7uyomlq26a_3s81cs qfij8isizuzcud2mhh515t1cluyq (
	.j0ln_h     (na29rv9xyz_vn       ), 
	.p2fq1i8       (obvunz7             ), 
	.pg17e0     (hhflrj5pivf         ), 
	.qqk5yk     (lr4pmtw0e3sm7         ), 
	.khfri3vm7  (                    ), 
	.x7bl2zxqiftsf  (                    ), 
	.kgg1udim46o  (                    )  
);

endmodule




















module qlm10lcv_tyz847h7k(
  input  [32-1:0]   wz0wek1lz0   ,
  output [6-1:0]    i8vml4gn      
);


wire [6-1:0] go6xtazzkuo27;

genvar i;

assign go6xtazzkuo27[0] = wz0wek1lz0[1] | wz0wek1lz0[3] | wz0wek1lz0[5] | wz0wek1lz0[7] | wz0wek1lz0[9] |
                         wz0wek1lz0[11] | wz0wek1lz0[13] | wz0wek1lz0[15] | wz0wek1lz0[17] | wz0wek1lz0[19] |
                         wz0wek1lz0[21] | wz0wek1lz0[23] | wz0wek1lz0[25] | wz0wek1lz0[27] | wz0wek1lz0[29] |
                         wz0wek1lz0[31];

assign go6xtazzkuo27[1] = wz0wek1lz0[1] | wz0wek1lz0[2] | wz0wek1lz0[5] | wz0wek1lz0[6] | wz0wek1lz0[9] |
                         wz0wek1lz0[10] | wz0wek1lz0[13] | wz0wek1lz0[14] | wz0wek1lz0[17] | wz0wek1lz0[18] |
                         wz0wek1lz0[21] | wz0wek1lz0[22] | wz0wek1lz0[25] | wz0wek1lz0[26] | wz0wek1lz0[29] |
                         wz0wek1lz0[30];

assign go6xtazzkuo27[2] = wz0wek1lz0[1] | wz0wek1lz0[2] | wz0wek1lz0[3] | wz0wek1lz0[4] |
                         wz0wek1lz0[9] | wz0wek1lz0[10] | wz0wek1lz0[11] | wz0wek1lz0[12] | 
                         wz0wek1lz0[17] | wz0wek1lz0[18] | wz0wek1lz0[19] | wz0wek1lz0[20] |
                         wz0wek1lz0[25] | wz0wek1lz0[26] | wz0wek1lz0[27] | wz0wek1lz0[28];

assign go6xtazzkuo27[3] = wz0wek1lz0[1] | wz0wek1lz0[2] | wz0wek1lz0[3] | wz0wek1lz0[4] |
                         wz0wek1lz0[5] | wz0wek1lz0[6] | wz0wek1lz0[7] | wz0wek1lz0[8] | 
                         wz0wek1lz0[17] | wz0wek1lz0[18] | wz0wek1lz0[19] | wz0wek1lz0[20] |
                         wz0wek1lz0[21] | wz0wek1lz0[22] | wz0wek1lz0[23] | wz0wek1lz0[24];

assign go6xtazzkuo27[4] = wz0wek1lz0[1] | wz0wek1lz0[2] | wz0wek1lz0[3] | wz0wek1lz0[4] |
                         wz0wek1lz0[5] | wz0wek1lz0[6] | wz0wek1lz0[7] | wz0wek1lz0[8] | 
                         wz0wek1lz0[9] | wz0wek1lz0[10] | wz0wek1lz0[11] | wz0wek1lz0[12] |
                         wz0wek1lz0[13] | wz0wek1lz0[14] | wz0wek1lz0[15] | wz0wek1lz0[16];

assign go6xtazzkuo27[5] = wz0wek1lz0[0];

assign i8vml4gn = go6xtazzkuo27;

endmodule

module h09sftk403rm5tnmsmed(
  input  [16-1:0]   wz0wek1lz0   ,
  output [5-1:0]    i8vml4gn      
);



wire [5-1:0] go6xtazzkuo27;

assign go6xtazzkuo27[0] = wz0wek1lz0[1] | wz0wek1lz0[3] | wz0wek1lz0[5] | wz0wek1lz0[7] | wz0wek1lz0[9] |
                         wz0wek1lz0[11] | wz0wek1lz0[13] | wz0wek1lz0[15];

assign go6xtazzkuo27[1] = wz0wek1lz0[1] | wz0wek1lz0[2] | wz0wek1lz0[5] | wz0wek1lz0[6] | wz0wek1lz0[9] |
                         wz0wek1lz0[10] | wz0wek1lz0[13] | wz0wek1lz0[14];

assign go6xtazzkuo27[2] = wz0wek1lz0[1] | wz0wek1lz0[2] | wz0wek1lz0[3] | wz0wek1lz0[4] |
                         wz0wek1lz0[9] | wz0wek1lz0[10] | wz0wek1lz0[11] | wz0wek1lz0[12];

assign go6xtazzkuo27[3] = wz0wek1lz0[1] | wz0wek1lz0[2] | wz0wek1lz0[3] | wz0wek1lz0[4] |
                         wz0wek1lz0[5] | wz0wek1lz0[6] | wz0wek1lz0[7] | wz0wek1lz0[8] ;

assign go6xtazzkuo27[4] = wz0wek1lz0[0];

assign i8vml4gn = go6xtazzkuo27;

endmodule

module sqkb0d8aic395m2pbugz(
  input  [8-1:0]   wz0wek1lz0   ,
  output [4-1:0]    i8vml4gn      
);



wire [4-1:0] go6xtazzkuo27;

assign go6xtazzkuo27[0] = wz0wek1lz0[1] | wz0wek1lz0[3] | wz0wek1lz0[5] | wz0wek1lz0[7];

assign go6xtazzkuo27[1] = wz0wek1lz0[1] | wz0wek1lz0[2] | wz0wek1lz0[5] | wz0wek1lz0[6];

assign go6xtazzkuo27[2] = wz0wek1lz0[1] | wz0wek1lz0[2] | wz0wek1lz0[3] | wz0wek1lz0[4];

assign go6xtazzkuo27[3] = wz0wek1lz0[0];

assign i8vml4gn = go6xtazzkuo27;

endmodule
























module gr40tady98ryto733e# (
  parameter yk7 = 1,  
  parameter m0qq = 2,  
  parameter dk34z = 4   
) (
  input  [64-1:0]    c5qrwj5sm0vc      ,     
  input  [64-1:0]    of4kpekzgop8    ,     
  input  [64-1:0]    l59fhx3o23g9ig ,     
  input  [64-1:0]    p2v9igi9t66348 ,     
  input  [31:0]              utwav9is_83yd6ng0 ,     
  input  [31:0]              sdmfqus_d4n5v3k ,     
  input  [15:0]              ghpvhjxwavld6r6r0w2 ,     
  input  [15:0]              berx62p9_hc2bfcnyn0 ,     
  input  [ 7:0]              ky3ucnc3e8n4c_iz  ,     
  input  [ 7:0]              v98eqhdqs8d1wk_qf2  ,     
  output                     p2tb25qpyet2a_c    ,     
  output                     wms1mxki5gyfyc    ,     
  output [yk7-1:0]            tkuhwm5tyjr    ,     
  output [yk7-1:0]            rg1trb_7w92    ,     
  output [m0qq-1:0]            a1bp0x22t5vu4q    ,     
  output [m0qq-1:0]            rgxbhxlvt61yfzn    ,     
  output [m0qq-1:0]            jpltrmmj8jw4lh_  ,     
  output [m0qq-1:0]            gs2s9lvzd_phhnv  ,     
  output [dk34z-1:0]            j694o6frj_680_g     ,     
  output [dk34z-1:0]            n2nedhasxux7buh     ,     
  output [dk34z-1:0]            fnv_7okzmo6y4ne85   ,     
  output [dk34z-1:0]            u_frczxmkmo88ujnp         
);


wire [64-1:0] vj13j6dx   = c5qrwj5sm0vc;
wire [64-1:0] o1nf132fggoqq = of4kpekzgop8;




wire [64-1:0] qkd3zrjfs6hqvtnl6t = p2v9igi9t66348;
wire [64-1:0] x9yoezqjjeerpzs023x = l59fhx3o23g9ig;
wire [64-1:0] mfezwn0l0a9xv8mb0f   = qkd3zrjfs6hqvtnl6t & vj13j6dx[64-1:0];
wire [64-1:0] pwys10lsmgmqlit_6nv   = (p2v9igi9t66348 & vj13j6dx[64-1:0]) | x9yoezqjjeerpzs023x;
assign p2tb25qpyet2a_c = (|mfezwn0l0a9xv8mb0f) & ~vj13j6dx[64-1];
assign wms1mxki5gyfyc = ~(&pwys10lsmgmqlit_6nv) & vj13j6dx[64-1];




wire [31:0] d9efhzvdbkejhrwier3 = sdmfqus_d4n5v3k;
wire [31:0] h7k91xg3de1zj2qvs1m1 = utwav9is_83yd6ng0;

wire [31:0] velblczas_2jbddkbnko_   [yk7-1:0];

wire [31:0] vtczb42p35qo4o51i   [yk7-1:0];


genvar i;
generate 

for(i=0;i<yk7;i=i+1) begin: fy2dpxp4t3rrne18
    assign velblczas_2jbddkbnko_[i]   = d9efhzvdbkejhrwier3 & vj13j6dx[i*32+31:i*32];
    
    assign vtczb42p35qo4o51i[i]   = (sdmfqus_d4n5v3k & vj13j6dx[i*32+31:i*32])   | h7k91xg3de1zj2qvs1m1;
    
    assign tkuhwm5tyjr[i]    = (|velblczas_2jbddkbnko_[i])  & ~vj13j6dx[i*32+31];  
    assign rg1trb_7w92[i]    = ~(&vtczb42p35qo4o51i[i]) & vj13j6dx[i*32+31];   
    
    
end

endgenerate





wire [15:0] o0s58vb_bij2l_tn = berx62p9_hc2bfcnyn0;
wire [15:0] ee1yq2r73cowetom = ghpvhjxwavld6r6r0w2;

wire [15:0] ez9j64e6lmt8cy3y23q   [m0qq-1:0];
wire [15:0] n3umto7lg8gduqjcjxycb [m0qq-1:0];
wire [15:0] fj4b8srq6ddbrlh   [m0qq-1:0];
wire [15:0] n2ysllysvvgcp8r59i [m0qq-1:0];

generate 

for(i=0;i<m0qq;i=i+1) begin: f84hlxqog_5e
    assign ez9j64e6lmt8cy3y23q[i]   = o0s58vb_bij2l_tn & vj13j6dx[i*16+15:i*16];
    assign n3umto7lg8gduqjcjxycb[i] = o0s58vb_bij2l_tn & o1nf132fggoqq[i*16+15:i*16];
    assign fj4b8srq6ddbrlh[i]   = (berx62p9_hc2bfcnyn0 & vj13j6dx[i*16+15:i*16])   | ee1yq2r73cowetom;
    assign n2ysllysvvgcp8r59i[i] = (berx62p9_hc2bfcnyn0 & o1nf132fggoqq[i*16+15:i*16]) | ee1yq2r73cowetom;
    assign a1bp0x22t5vu4q[i]    = (|ez9j64e6lmt8cy3y23q[i])  & ~vj13j6dx[i*16+15];  
    assign rgxbhxlvt61yfzn[i]    = ~(&fj4b8srq6ddbrlh[i]) & vj13j6dx[i*16+15];   
    assign jpltrmmj8jw4lh_[i]  = (|n3umto7lg8gduqjcjxycb[i])  & ~o1nf132fggoqq[i*16+15];
    assign gs2s9lvzd_phhnv[i]  = ~(&n2ysllysvvgcp8r59i[i]) & o1nf132fggoqq[i*16+15]; 
end

endgenerate





wire [7:0] dcyaauth9qlxj39f9m = v98eqhdqs8d1wk_qf2;
wire [7:0] lf38o8thk7u2fzwbfddo = ky3ucnc3e8n4c_iz;

wire [7:0] yjx1b8mgu49i_g1bgz   [dk34z-1:0];
wire [7:0] zemurk6gd_jud5jmmbhz_ [dk34z-1:0];
wire [7:0] zx5k6q6x4s_a64mx10w   [dk34z-1:0];
wire [7:0] ew7m6fdfep2vqvd5c0cxsm [dk34z-1:0];

generate 

for(i=0;i<dk34z;i=i+1) begin: q0wo53h6xzu
    assign yjx1b8mgu49i_g1bgz[i]   = dcyaauth9qlxj39f9m & vj13j6dx[i*8+7:i*8];
    assign zemurk6gd_jud5jmmbhz_[i] = dcyaauth9qlxj39f9m & o1nf132fggoqq[i*8+7:i*8];
    assign zx5k6q6x4s_a64mx10w[i]   = (v98eqhdqs8d1wk_qf2 & vj13j6dx[i*8+7:i*8])   | lf38o8thk7u2fzwbfddo;
    assign ew7m6fdfep2vqvd5c0cxsm[i] = (v98eqhdqs8d1wk_qf2 & o1nf132fggoqq[i*8+7:i*8]) | lf38o8thk7u2fzwbfddo;
    assign j694o6frj_680_g[i]    = (|yjx1b8mgu49i_g1bgz[i])  & ~vj13j6dx[i*8+7];  
    assign n2nedhasxux7buh[i]    = ~(&zx5k6q6x4s_a64mx10w[i]) & vj13j6dx[i*8+7];   
    assign fnv_7okzmo6y4ne85[i]  = (|zemurk6gd_jud5jmmbhz_[i])  & ~o1nf132fggoqq[i*8+7];
    assign u_frczxmkmo88ujnp[i]  = ~(&ew7m6fdfep2vqvd5c0cxsm[i]) & o1nf132fggoqq[i*8+7]; 
end

endgenerate

endmodule























module rkhmkn86ap95zo99(

  
  
  
  
  input  [64-1:0] artnbioj,
  input  [64-1:0] emfjxicm,
  input  [64-1:0] ehzolf0,
  input  [5-1:0] fhhe7189lmum,
  input  [5-1:0] cpt0qfwiz, 
  input  [4-1:0] ker4nfxz2b_p53w,  

  
  
  
  
  output vjkz8n6i44pc7o,                     
  
  output cwmxezrc3jv6hzxcfc,   
  input  uig3ujuyq0_61kqb,   
  output [64-1:0] nb3w1rq_ny95rvrt,
  output xc2becmsn4fcniw6ks,

  
  
  
  output [4-1:0] p_yx415so7q1vohijb,
  
  input  j_rvclhfbeig5cqeb3_,

  
  
  
  input  [105-1:0] e19iv2rqeu5,
  input  [50-1:0] m4y6v4ncsg,

  
  
  
  output wkzq9xwwp9c3wcf3616c,
  output juy4d3jn2_92c7jefm1i6,
  output [64-1:0] qebmlqd6ka70065zibcx,
  output [64-1:0] hftmbp4yfjjsgcltu,
  input  [64-1:0] iont49tufvh5v7eetbw0m,
  input  [64-1:0] u2yurbi1gylta0pv_xpnz8ppo,

  
  
  
  input  ictx5fosbsup6y,         
  output s66_nzq5i23lbo,         

  output v51v27wp_7tuha,         
  input  isrgf76t7pxi,         



  
  
  
  input  gf33atgy,
  input  ru_wi

  );

  localparam ctu6y0yy1_ = 6;






  wire [64-1:0]              amgi_rqhtd007    = artnbioj;
  wire [64-1:0]              g7tawq8tp6    = emfjxicm;
  wire [64-1:0]              xo5bwsw4j8a     = ehzolf0;
  wire [64-1:0]              jmf1rwo8     = ehzolf0;
  wire  [5-1:0]      bj9det3k1xe2rn  = fhhe7189lmum;
  wire  [5-1:0]      cvhwe_6rucj7 = cpt0qfwiz; 
  wire [105-1:0] xlkm1ikvsatc2   = e19iv2rqeu5;
  wire [50-1:0] n6izg3jvgts   = m4y6v4ncsg;


  wire [105-1:0] nhqiwwnz4lmleg;
  wire [105-1:0] w98a0gvni829u3;
  wire [105-1:0] p8svuggnu7zvtlojt;
  wire [105-1:0] ykn2abyw7s2voefu;
  wire [105-1:0] wazt073vrvkujb_lpjze6;
  wire [105-1:0] azvwipii1valwcdp80j3_oq;
  wire [105-1:0] no56h0p6kag9edi57joc3m;

  wire ln4s1h4obzzo         = w98a0gvni829u3[95   ]
                          | w98a0gvni829u3[96  ]
                          ;

  wire ba2tpl29cmvgrvl1qqqz_qp = n6izg3jvgts[18];
  wire sr2ad0lhuts5ctwnepl5 = n6izg3jvgts[19];
  wire n5_0tyghia5to9pq5a2 = n6izg3jvgts[20];
  wire vu8cn0tjzmmmjqj_9 = ba2tpl29cmvgrvl1qqqz_qp | sr2ad0lhuts5ctwnepl5 | n5_0tyghia5to9pq5a2;
  wire y_0id5h2cb8ukkao        = n6izg3jvgts[22];
  wire yg_3i0cfu6iwmj       = n6izg3jvgts[23];
  wire hxv8akm9tnbagx         = n6izg3jvgts[14];
  wire qhmdzlcppcq8       = n6izg3jvgts[15];

  wire t_998ilixet4pdvdkju = y_0id5h2cb8ukkao | vu8cn0tjzmmmjqj_9 | yg_3i0cfu6iwmj; 


  assign wazt073vrvkujb_lpjze6 = {105{ba2tpl29cmvgrvl1qqqz_qp}} & xlkm1ikvsatc2;
  assign azvwipii1valwcdp80j3_oq = {105{sr2ad0lhuts5ctwnepl5}} & xlkm1ikvsatc2;
  assign no56h0p6kag9edi57joc3m = {105{n5_0tyghia5to9pq5a2}} & xlkm1ikvsatc2;
  assign nhqiwwnz4lmleg         = {105{hxv8akm9tnbagx}}         & xlkm1ikvsatc2;
  assign p8svuggnu7zvtlojt        = {105{y_0id5h2cb8ukkao}}        & xlkm1ikvsatc2;
  assign w98a0gvni829u3       = {105{qhmdzlcppcq8}}       & xlkm1ikvsatc2;
  assign ykn2abyw7s2voefu       = {105{yg_3i0cfu6iwmj}}       & xlkm1ikvsatc2;


  wire [64-1:0] aiiy8pexinn1bnd0jyoy6;
  wire z1hnaq01roqg6md1i028mg;
 
  





  
  
  wire [64-1:0] adydub7ly8l0x30v1_ivlfc;
  wire pqzn02_fhxv85bpjep7;


  wire [64-1:0] ya1whb4lzd9i6g2qr2yu5enshd   ;
  wire kxetexnh8sgpjk6cvyf4;







  wire [80-1:0] ray06eatktnsi4mn5w   ;
  wire [80-1:0] ixi02l50nmppg67yeekep   ; 
  wire [80-1:0] hqcobkfvvt1l5b4u9ke3jl0x8;
  wire [80-1:0] obkn6tbb4pes5xvb82ypx8ng2;
  wire [80-1:0] cl0tcivvt46muh82na        ; 
  wire [80-1:0] tktysetch337p4xj     ;
  wire [64+3:0] xcp0v_slt0baqx9h6px    ;
  wire                                mmdmrxttxmiz27        ;
  wire                                dso4rrx46c88           ;
  wire ae_pf3b_6qfu__950y636t = vu8cn0tjzmmmjqj_9 | ln4s1h4obzzo; 

  wire [64-1:0]               mnqd528vibxlk8k   = {64{ae_pf3b_6qfu__950y636t}} & amgi_rqhtd007;
  wire [64-1:0]               oaor6bvy1fu7flvavd   = {64{ae_pf3b_6qfu__950y636t}} & g7tawq8tp6;

  g_fo67k2g__407yyem_ bq1se8yvkdtiaq2fskck55(

      .m35ros_bzlaqo8y319z           ( mnqd528vibxlk8k         ),
      .uq5g_s44gt3h0fbg4zzv           ( oaor6bvy1fu7flvavd         ),
      .i8whgk1t5jsbvv8u3ojllu7         (64'b0),
      .c7cw30bh940izgc1knsjmx         (64'b0),
      .f63_o3d0oy82l6owdiogb9dqm     ( wazt073vrvkujb_lpjze6   ), 
      .uew_1l_6faqgtso37h_zds7     ( azvwipii1valwcdp80j3_oq   ), 
      .qtiogf3y1fz2gfxknzswuj     ( no56h0p6kag9edi57joc3m   ), 
      .vqnbcwzo10cg732u0           ( w98a0gvni829u3         ),

      .lbo2x74bznoaaigmxjenghis       ( cl0tcivvt46muh82na          ),
      .lm4nz97neurpj88xyqm7n8hi_c37    (),

      .s6tonq08_ria84ebdjlir           ( xcp0v_slt0baqx9h6px      ),
      .ya1whb4lzd9i6g2qr2yu5enshd     ( ya1whb4lzd9i6g2qr2yu5enshd ),
      .fl1olcli4mhazuy960y16sqh63s5   (),
      .gm0zk3gsgqtkn9_jovpqw3       ( ray06eatktnsi4mn5w     ),
      .yzauwl2y3mmfl_dtz0c89ze2       ( ixi02l50nmppg67yeekep     ),
      .p_q6uot8vlny0p1532oethvbx67    ( hqcobkfvvt1l5b4u9ke3jl0x8  ),
      .e9_hqyec0sd5hbt8qhk_tt_7mhn    ( obkn6tbb4pes5xvb82ypx8ng2  ),
      .cxxjqchsz57vq2dff3d0j       ( kxetexnh8sgpjk6cvyf4     ),

      .ymi25pa6qmirfeb9            ( mmdmrxttxmiz27          ),
      .iz4sa6lcipb1cjsz_               ( dso4rrx46c88             )
  );





  wire jjct59z68fasiq3hkv;
  wire iza744k4kjssx = mmdmrxttxmiz27 | jjct59z68fasiq3hkv;
  wire v47mqk8gjeayfhjz = n6izg3jvgts[21];

  wire [80-1:0] k7kw5knwr6540jutk5rnw;
  wire [80-1:0] r5zcjbkhohovwi9u0omvr;

  wire gq8y1doymz9nz247a7 = (mmdmrxttxmiz27 & dso4rrx46c88);

  wire [80-1:0] k9wo3uwsknspc4mtccve0  = ({80{mmdmrxttxmiz27}} & hqcobkfvvt1l5b4u9ke3jl0x8) ;

  wire [80-1:0] mu9og1s6qa3g3z_on7a8_awx  = ({80{mmdmrxttxmiz27}} & obkn6tbb4pes5xvb82ypx8ng2);

  wire [80-1:0] nw8l2uwwk8eun92i2d = ({80{mmdmrxttxmiz27}} & ray06eatktnsi4mn5w);

  wire [80-1:0] azcrrtpprsyrifk44 = ({80{mmdmrxttxmiz27}} & ixi02l50nmppg67yeekep);

  wire [321-1:0] yxz7x3t8z5j2cc0 =  {
                                                             gq8y1doymz9nz247a7     ,
                                                             k9wo3uwsknspc4mtccve0 ,
                                                             mu9og1s6qa3g3z_on7a8_awx ,
                                                             nw8l2uwwk8eun92i2d    ,
                                                             azcrrtpprsyrifk44    
                                                           };

  wire [321-1:0] v6wp4yeifqw_49xe  =  {
                                                             1'b0                        ,
                                                             80'b0 ,
                                                             80'b0 ,
                                                             k7kw5knwr6540jutk5rnw           ,
                                                             r5zcjbkhohovwi9u0omvr            
                                                           };


  wire [321-1:0] xe3uwuwthp      =  
                                                             ({321{mmdmrxttxmiz27}}     & yxz7x3t8z5j2cc0)
                                                           | ({321{jjct59z68fasiq3hkv}}     & v6wp4yeifqw_49xe)
                                                           ; 

  wire qp5zhaxmki = xe3uwuwthp[321-1];
  wire [80-1:0] ebyjq8t8vcorpng_5    = xe3uwuwthp[(80*2)-1:80];
  wire [80-1:0] np2skrwpa7s8vyu5_    = xe3uwuwthp[80-1:0];
  wire [80-1:0] wdi7t_m7a3uueuy4h = xe3uwuwthp[(80*2)+80-1:80*2];
  wire [80-1:0] q32shhpbei8myfzfayq = xe3uwuwthp[(80*2)+(80*2)-1:(80*2)+80];

  otwg2iaolmlgo34d69 wwr8d0r7r0ir0ej_3wq31cl(

      .cattuehkeqxtxg_y           ( iza744k4kjssx              ),
      .pw_vsq5tj5cykojr9ce4i         ( v47mqk8gjeayfhjz           ),      
      .owwzmmptdds6_we3no8q5           ( qp5zhaxmki                 ),

      .j3998mrey0wg8bqs4j9         (80'b0),
      .r92fvyocvp3upr8yj2g_         (80'b0),
      .kcc7r7vj7sjmae15bm_lvgt         (),

      .tjzp46d5wrtx640f            ( ebyjq8t8vcorpng_5          ),
      .q_wbix0_hlxllb5l10k            ( np2skrwpa7s8vyu5_          ), 
      .c1chm8mj_hlw8ru4c            ( cl0tcivvt46muh82na          ) 
  );









  wire sa51f1uubzvo0drqlo5;
  wire kmwyjy2334kq0grn1tg = 1'b0;
  wire [64-1:0] item2h0zpygqk9zeo;
  wire [ctu6y0yy1_-1:0] ya8hvm7f9s08f3d6;

  wire elzi9vcfgv5dfbn = sa51f1uubzvo0drqlo5 | kmwyjy2334kq0grn1tg;



  wire dxenquvmssguef0xhphhd_5m34;
  wire vj822xzl2px_z9xo3p28x59sizh = 1'b0;
  wire [64-1:0] nilxioo2gee_2g7dp;
  wire [ctu6y0yy1_-1:0] wlzbrha6e20dndaxd;

  wire z__fluu2ul_ds1yckdmjt = dxenquvmssguef0xhphhd_5m34 | vj822xzl2px_z9xo3p28x59sizh;



  wire b4_p52l0f5v37nqqq;
  wire sll0_4d8ngfpyh8lw4i;
  wire [64-1:0] zrjp4odho_;
  
  wire [ctu6y0yy1_-1:0]      by2bmev01awcb;
  
  wire t_dpnebd3dc = b4_p52l0f5v37nqqq | sll0_4d8ngfpyh8lw4i;




  
  wire ixilll769h9ctg4mrz  = ykn2abyw7s2voefu[24];
  wire opp55w_ujnk6ukodr1 = ykn2abyw7s2voefu[39];
  wire jfdp5zy_q2woeffi = ixilll769h9ctg4mrz | opp55w_ujnk6ukodr1; 
  wire h5jozrobnaxu2nqwmzv5ur;

  wire [64-1:0] r6coxdlvt72jfaw2ix_5x;
  wire [64-1:0] nab43_gl6qeifr516shtri;
  wire [64-1:0] haryili5jw0sv_jegpnpcq;

  wire rdum446o_8f6mp1iuf83ghngwk  = jfdp5zy_q2woeffi & sll0_4d8ngfpyh8lw4i;
  wire qixww3rvwwddqzrbt2ov5qindlh_ = jfdp5zy_q2woeffi & b4_p52l0f5v37nqqq;

  wire [64-1:0]  vurcuwbrjgbzpgtreom_du0 = 64'b0;
  wire [64-1:0]  wyi9ffifr4fwp310f5s9o = 64'b0;
  

  assign wkzq9xwwp9c3wcf3616c =  h5jozrobnaxu2nqwmzv5ur | rdum446o_8f6mp1iuf83ghngwk;
  assign juy4d3jn2_92c7jefm1i6 =  qixww3rvwwddqzrbt2ov5qindlh_;
  assign qebmlqd6ka70065zibcx =  h5jozrobnaxu2nqwmzv5ur ? r6coxdlvt72jfaw2ix_5x
                                                     : vurcuwbrjgbzpgtreom_du0;

  assign hftmbp4yfjjsgcltu =  h5jozrobnaxu2nqwmzv5ur ? nab43_gl6qeifr516shtri
                                                     : wyi9ffifr4fwp310f5s9o;

  wire v6y4aokp2429rlzqtj;
  wire vhph5rtzyw47zuy3s;
  wire dx2o2oi401iz;
  wire [64-1:0] fshrsdciyi905ku7;
  wire [ctu6y0yy1_-1:0]      wlxoir8fm329rj;
  wire [64-1:0] lh7ry3p923qgxhqegq;
  wire [64-1:0] bt1lqldb4uavr0gx47htp;
  wire [64-1:0] rd5gqwxxtmt2puus6k5a;
  wire [64-1:0] y_6lwsra9xergl478k2fh;


  assign haryili5jw0sv_jegpnpcq   = iont49tufvh5v7eetbw0m;
  assign bt1lqldb4uavr0gx47htp = u2yurbi1gylta0pv_xpnz8ppo; 
  assign y_6lwsra9xergl478k2fh  = iont49tufvh5v7eetbw0m; 
  assign v6y4aokp2429rlzqtj = sa51f1uubzvo0drqlo5 | dxenquvmssguef0xhphhd_5m34 | b4_p52l0f5v37nqqq;
  assign vhph5rtzyw47zuy3s  = kmwyjy2334kq0grn1tg  | vj822xzl2px_z9xo3p28x59sizh  | sll0_4d8ngfpyh8lw4i;
  assign dx2o2oi401iz       = v6y4aokp2429rlzqtj | vhph5rtzyw47zuy3s;

  assign fshrsdciyi905ku7 =  
                          ({64{elzi9vcfgv5dfbn      }} & item2h0zpygqk9zeo     )
						| ({64{z__fluu2ul_ds1yckdmjt }} & nilxioo2gee_2g7dp)
						| ({64{t_dpnebd3dc         }} & zrjp4odho_        )
						;

  assign wlxoir8fm329rj =  
                          ({ctu6y0yy1_{elzi9vcfgv5dfbn      }} & ya8hvm7f9s08f3d6     )
						| ({ctu6y0yy1_{z__fluu2ul_ds1yckdmjt }} & wlzbrha6e20dndaxd)
						| ({ctu6y0yy1_{t_dpnebd3dc         }} & by2bmev01awcb        )
						;



  uq9oowb3c0mb0eda15rcw5 # (
  	.ctu6y0yy1_ (ctu6y0yy1_)  
  )
  j5vqtsg_rmno7uu_4fikzn6u(
  	.f218verzay1lfg_t73r7h         ( v6y4aokp2429rlzqtj     ),
  	.wvyn3jdt7m5qk570c1zta          ( vhph5rtzyw47zuy3s      ),
  	.v2k5ixyb1cco74jghjt               ( fshrsdciyi905ku7           ),
  	.mhres_bf8ykyi80s               ( wlxoir8fm329rj           ),
  	.jhqv9u46f4ilao8a7rqc         ( lh7ry3p923qgxhqegq     ),
  	.en2fwj8b2lksbcaz8_f          ( rd5gqwxxtmt2puus6k5a      )
  );




  
  wire [64-1:0] g4ucoelbw2f13   = ({64{yg_3i0cfu6iwmj}} & amgi_rqhtd007);
  wire [64-1:0] t55mrbjc_fc_1v   = ({64{yg_3i0cfu6iwmj}} & g7tawq8tp6);

  aiw2b4qk64vf3344ezyf # (
  	.ctu6y0yy1_(ctu6y0yy1_)  
  )
  muge_4qe49s4rqnguzdr(
  	.amgi_rqhtd007                    ( g4ucoelbw2f13          ),
  	.otn5ycgat1c9s1a                  (64'b0),
  	.g7tawq8tp6                    ( t55mrbjc_fc_1v          ),  
  	.xlkm1ikvsatc2                   ( ykn2abyw7s2voefu         ),
  	.g36_kozc0w4bjtnf                  ( jjct59z68fasiq3hkv          ),
  	.ileuocpyluq                  ( k7kw5knwr6540jutk5rnw      ),
  	.yiexcriz0ufmy                  ( r5zcjbkhohovwi9u0omvr      ),
  	.e231c11ou7ube_b                  ( cl0tcivvt46muh82na          ),
  	.tppbcuxfcn35ghrqja5            ( b4_p52l0f5v37nqqq        ),
  	.iv4pxzd85kko8e8twyro             ( sll0_4d8ngfpyh8lw4i         ),
  	.ixlv8n_7cgrz2                  ( zrjp4odho_              ),
  	.gxtsmhtras93dt4g11                (),
  	.i8fcutzmv9eer                  ( by2bmev01awcb              ),
  	.kth4tafeif3978quzt            ( lh7ry3p923qgxhqegq     ),
  	.eltrj3g68c3h11e7zli4x0t9          (64'b0),
  	.u9d99u2san4lbuhbb             ( rd5gqwxxtmt2puus6k5a      ),
  	.xlxi2zedzir0xwdjxt           (64'b0),
  	.nb3w1rq_ny95rvrt              ( aiiy8pexinn1bnd0jyoy6  ),
  	.dkojj6fim0nxg4jvyafk            (),
  	.vjkz8n6i44pc7o                ( z1hnaq01roqg6md1i028mg    )
  );




  
  
  wire [64-1:0] ky4112jmao_ii = ({64{y_0id5h2cb8ukkao}} & amgi_rqhtd007);
  wire [64-1:0] w2jwy3yhck4bvr = ({64{y_0id5h2cb8ukkao}} & g7tawq8tp6);

  i6tr_dyutx06rp9skham4 # (
  	.ctu6y0yy1_(ctu6y0yy1_)  
  )
  qbwaik87a4x2whuuuu1_mc (
  	.amgi_rqhtd007                    ( ky4112jmao_ii             ),
  	.h33_crpt0l75o                 (64'b0), 
  	.g7tawq8tp6                    ( w2jwy3yhck4bvr             ),
  	.jmf1rwo8                     ( jmf1rwo8                 ), 
  	.xo5bwsw4j8a                     ( xo5bwsw4j8a                 ), 
  	.xlkm1ikvsatc2                   ( p8svuggnu7zvtlojt            ),
  	.lzal8kswefl9gv4kqdclkfx23         ( sa51f1uubzvo0drqlo5       ),
  	.udhgtu0ck3hr1aj               ( item2h0zpygqk9zeo             ),
  	.so4zxlxtb1t9lx               ( ya8hvm7f9s08f3d6             ),
  	.q7c4bjf1j8kujxtvei               ( lh7ry3p923qgxhqegq       ),
  	.bdd_smghkpbtvkxlxpdyq2perm    ( dxenquvmssguef0xhphhd_5m34  ),
  	.sznwd73uhzrymh69lt9dcfpa          ( nilxioo2gee_2g7dp        ),
  	.l4ik_e9aa1bhu66b138          ( wlzbrha6e20dndaxd        ),
  	.zvnjpa2uy_h98fk1u8zei9w          ( lh7ry3p923qgxhqegq       ),
  	.sazh4of6fhumdu0qyo1yjk2u00eee     ( h5jozrobnaxu2nqwmzv5ur   ),
  	.m9e0b_s90djin0iqc0ts9v          ( r6coxdlvt72jfaw2ix_5x        ),
  	.yqf19lhru49yxe2r5x0diu          ( nab43_gl6qeifr516shtri        ),
  	.yhru2nhdb63arfxbb25pgcp          ( haryili5jw0sv_jegpnpcq        ),  
  	.nb3w1rq_ny95rvrt              ( adydub7ly8l0x30v1_ivlfc     ),
  	.vjkz8n6i44pc7o                ( pqzn02_fhxv85bpjep7       ),
  	.m6ouh9hkcy63fxj02                ( y_0id5h2cb8ukkao              ),
  	.gf33atgy                          ( gf33atgy                      ),
  	.ru_wi                        ( ru_wi                    )
  );




  
  wire  w363n7ci30h3kw2g1oktlj1puysbju;    
  wire  lygqe2977b3fd_0eit3wg_nnfirn;    
  wire th583ebkp2cj56crsivefzygk81o65_h2;
  wire  vz2rm7lc9ctulrdhe1kv8wdmobft;    
  wire hlmhgsbtxsmi7y1a7oshnntydp27pj;
  wire dshcfm3k8zhyftxq_xw9j106j59z7notf;
  wire  gdebc5b6o6bv57ax1bw;
  
  
  wire [64-1:0] nx4gyto1vnfvb7wx   = amgi_rqhtd007;
  wire [64-1:0] n9r03am0pez   = g7tawq8tp6;
  wire [63:0] usrh37qm6nz8yamj6_h_pmbv5;
  wire [63:0] mipc_c8bfwk8khoqgtsj65f1f;
  wire [63:0] pm3m6aucefl9oas0vqgwfm;
  wire [63:0] yc5f_bw94gu1iari4qpmo269z;

  qhqypfyt2lgewc2ne9xw pvyf6sg7jq3de18vn_1pigf(
   .a4p3huz_qaf92as          (nhqiwwnz4lmleg),
   .e4_5otstd9ttd5eebgmf        (w98a0gvni829u3),
   .n6izg3jvgts              (n6izg3jvgts),
   .amgi_rqhtd007               (nx4gyto1vnfvb7wx),
   .g7tawq8tp6               (n9r03am0pez),
   .w363n7ci30h3kw2g1oktlj1puysbju    (w363n7ci30h3kw2g1oktlj1puysbju),
   .lygqe2977b3fd_0eit3wg_nnfirn      (lygqe2977b3fd_0eit3wg_nnfirn),
  .th583ebkp2cj56crsivefzygk81o65_h2(th583ebkp2cj56crsivefzygk81o65_h2),
  .vz2rm7lc9ctulrdhe1kv8wdmobft  (vz2rm7lc9ctulrdhe1kv8wdmobft),
  .hlmhgsbtxsmi7y1a7oshnntydp27pj  (hlmhgsbtxsmi7y1a7oshnntydp27pj),
  .dshcfm3k8zhyftxq_xw9j106j59z7notf(dshcfm3k8zhyftxq_xw9j106j59z7notf),
  
   
   .usrh37qm6nz8yamj6_h_pmbv5    (usrh37qm6nz8yamj6_h_pmbv5),
   .mipc_c8bfwk8khoqgtsj65f1f    (mipc_c8bfwk8khoqgtsj65f1f),
   .pm3m6aucefl9oas0vqgwfm    (pm3m6aucefl9oas0vqgwfm),
   .yc5f_bw94gu1iari4qpmo269z    (yc5f_bw94gu1iari4qpmo269z),
   .gdebc5b6o6bv57ax1bw      (gdebc5b6o6bv57ax1bw)
  );

  wire [64-1:0] azehbzuwas1onyt65   = {64{qhmdzlcppcq8}} & amgi_rqhtd007;
  wire [64-1:0] pcko5kg7h0yh1z    = {64{qhmdzlcppcq8}} & xo5bwsw4j8a;
  wire [64-1:0] l7mctsr6ttfp83pl8jo7;
  wire a2o96wlgs_5sqzm2a7ba_;

  a37xq53sqhw4q7cxzwmz  g336vkeo9czv_mcd57bxpyj2s(
  .tvdvyldvwqhx7g8r9di         (ictx5fosbsup6y),
  .izj2me9tmzxitrpzl1tr         (s66_nzq5i23lbo),
  .rgcs7q5ke7h8fte8jecm         (v51v27wp_7tuha),
  .pzhh8hyzbdb80ac8sdd_49         (isrgf76t7pxi),
  .t_998ilixet4pdvdkju          (t_998ilixet4pdvdkju),
  .l7mctsr6ttfp83pl8jo7      (l7mctsr6ttfp83pl8jo7),
  .a2o96wlgs_5sqzm2a7ba_          (a2o96wlgs_5sqzm2a7ba_),
  .cwmxezrc3jv6hzxcfc    (cwmxezrc3jv6hzxcfc),
  .uig3ujuyq0_61kqb    (uig3ujuyq0_61kqb),
  .j_rvclhfbeig5cqeb3_         (j_rvclhfbeig5cqeb3_),
  .gdebc5b6o6bv57ax1bw          (gdebc5b6o6bv57ax1bw),
  .w363n7ci30h3kw2g1oktlj1puysbju(w363n7ci30h3kw2g1oktlj1puysbju),
  .lygqe2977b3fd_0eit3wg_nnfirn  (lygqe2977b3fd_0eit3wg_nnfirn),
  .th583ebkp2cj56crsivefzygk81o65_h2(th583ebkp2cj56crsivefzygk81o65_h2),
  .vz2rm7lc9ctulrdhe1kv8wdmobft  (vz2rm7lc9ctulrdhe1kv8wdmobft),
  .hlmhgsbtxsmi7y1a7oshnntydp27pj  (hlmhgsbtxsmi7y1a7oshnntydp27pj),
  .dshcfm3k8zhyftxq_xw9j106j59z7notf(dshcfm3k8zhyftxq_xw9j106j59z7notf),
  .bj9det3k1xe2rn               (bj9det3k1xe2rn),
  .cvhwe_6rucj7              (cvhwe_6rucj7),
  .amgi_rqhtd007                 (azehbzuwas1onyt65),
  .xo5bwsw4j8a                  (pcko5kg7h0yh1z),
  .usrh37qm6nz8yamj6_h_pmbv5      (usrh37qm6nz8yamj6_h_pmbv5),
  .mipc_c8bfwk8khoqgtsj65f1f      (mipc_c8bfwk8khoqgtsj65f1f),
  .pm3m6aucefl9oas0vqgwfm      (pm3m6aucefl9oas0vqgwfm),
  .yc5f_bw94gu1iari4qpmo269z      (yc5f_bw94gu1iari4qpmo269z),
  .xcp0v_slt0baqx9h6px         (xcp0v_slt0baqx9h6px),
  .a4p3huz_qaf92as            (nhqiwwnz4lmleg),
  .e4_5otstd9ttd5eebgmf          (w98a0gvni829u3),
  .n6izg3jvgts                (n6izg3jvgts),
  .jsz4fvx2s3ijb5            (ker4nfxz2b_p53w),
  .vjkz8n6i44pc7o             (vjkz8n6i44pc7o),
  .nb3w1rq_ny95rvrt           (nb3w1rq_ny95rvrt),        
  .xc2becmsn4fcniw6ks            (xc2becmsn4fcniw6ks),        
  .p_yx415so7q1vohijb           (p_yx415so7q1vohijb),
  .gf33atgy                       (gf33atgy),
  .ru_wi                     (ru_wi)
  );





  assign l7mctsr6ttfp83pl8jo7 =  
                             ({64{yg_3i0cfu6iwmj}} & aiiy8pexinn1bnd0jyoy6)       
                           | ({64{y_0id5h2cb8ukkao}} & adydub7ly8l0x30v1_ivlfc)
                           | ({64{vu8cn0tjzmmmjqj_9}} & ya1whb4lzd9i6g2qr2yu5enshd)
                           
                           ;


  assign a2o96wlgs_5sqzm2a7ba_   = 
                             (yg_3i0cfu6iwmj  & z1hnaq01roqg6md1i028mg)       
                           | (y_0id5h2cb8ukkao   & pqzn02_fhxv85bpjep7)
                           | (vu8cn0tjzmmmjqj_9 & kxetexnh8sgpjk6cvyf4)
                           
                           ;
  

endmodule




















module otwg2iaolmlgo34d69 (

  input  cattuehkeqxtxg_y,
  input  pw_vsq5tj5cykojr9ce4i,
  input  owwzmmptdds6_we3no8q5,

  input  [80-1:0] j3998mrey0wg8bqs4j9,
  input  [80-1:0] r92fvyocvp3upr8yj2g_,
  output [80-1:0] kcc7r7vj7sjmae15bm_lvgt, 

  input  [80-1:0] tjzp46d5wrtx640f   ,
  input  [80-1:0] q_wbix0_hlxllb5l10k   , 
  output [80-1:0] c1chm8mj_hlw8ru4c
  );











  
  
  
  

  localparam h8hbjimfai3byrx8du67czk7ob5 = ((80*2)+(80*2)+1); 

  wire mm3q580thw0s;
  wire [80-1:0] az6qlcqsx_0  ;
  wire [80-1:0] cqqzeukmh  ; 
  wire [80-1:0] s72up0gw70;
  wire [80-1:0] r1065fzikc4ea;



  assign  {
    az6qlcqsx_0
   ,cqqzeukmh
   ,s72up0gw70
   ,r1065fzikc4ea
   ,mm3q580thw0s
    }
    = 
        ({h8hbjimfai3byrx8du67czk7ob5{cattuehkeqxtxg_y}} & {
             tjzp46d5wrtx640f   
            ,q_wbix0_hlxllb5l10k   
            ,j3998mrey0wg8bqs4j9
            ,r92fvyocvp3upr8yj2g_
            ,owwzmmptdds6_we3no8q5
          })
        ;

     
  wire [80-1:0] do_4d6t05wx7ap = az6qlcqsx_0;
  wire [80-1:0] gh1pq3ezuu8hf = cqqzeukmh;
  wire eaakrh1bs245q = mm3q580thw0s;
  wire [80-1:0] cl0tcivvt46muh82na = do_4d6t05wx7ap + gh1pq3ezuu8hf + eaakrh1bs245q;

  wire [80-1:0] tktysetch337p4xj = {80{1'b0}};

  assign c1chm8mj_hlw8ru4c    = cl0tcivvt46muh82na    ;
  assign kcc7r7vj7sjmae15bm_lvgt = tktysetch337p4xj ;

endmodule                                      
                                               






















module g_fo67k2g__407yyem_(

  
  
  
  input  [64-1:0] m35ros_bzlaqo8y319z  ,
  input  [64-1:0] uq5g_s44gt3h0fbg4zzv  ,
  input  [64-1:0] i8whgk1t5jsbvv8u3ojllu7,
  input  [64-1:0] c7cw30bh940izgc1knsjmx,
  input  [105-1:0] f63_o3d0oy82l6owdiogb9dqm,
  input  [105-1:0] uew_1l_6faqgtso37h_zds7,
  input  [105-1:0] qtiogf3y1fz2gfxknzswuj,
  input  [105-1:0] vqnbcwzo10cg732u0,

  
  
  


  

  output [64+3:0] s6tonq08_ria84ebdjlir,
  output [64-1:0] ya1whb4lzd9i6g2qr2yu5enshd,
  output [64-1:0] fl1olcli4mhazuy960y16sqh63s5,
  output cxxjqchsz57vq2dff3d0j, 


  
  
  
  
  
  output [80-1:0] gm0zk3gsgqtkn9_jovpqw3   ,
  output [80-1:0] yzauwl2y3mmfl_dtz0c89ze2   ,
  output [80-1:0] p_q6uot8vlny0p1532oethvbx67,
  output [80-1:0] e9_hqyec0sd5hbt8qhk_tt_7mhn,
  output ymi25pa6qmirfeb9,
  output iz4sa6lcipb1cjsz_,

  input  [80-1:0] lbo2x74bznoaaigmxjenghis   ,
  input  [80-1:0] lm4nz97neurpj88xyqm7n8hi_c37 

  );


  
  wire p4diuazqfby     = f63_o3d0oy82l6owdiogb9dqm[5   ];
  wire u1mn5wzoquj0    = f63_o3d0oy82l6owdiogb9dqm[6  ];
  wire nn8f1wf_9ovyh   = f63_o3d0oy82l6owdiogb9dqm[7 ];
  wire ye2b0mu4    = f63_o3d0oy82l6owdiogb9dqm[8  ];
  wire wsflp3hzxrkbzt   = f63_o3d0oy82l6owdiogb9dqm[9 ];
  wire i8joes9bj   = f63_o3d0oy82l6owdiogb9dqm[10 ];
  wire tguh9z4uqcbc     = f63_o3d0oy82l6owdiogb9dqm[11   ];
  wire sudgj682o    = f63_o3d0oy82l6owdiogb9dqm[12  ];
  wire goy125ul4oyvze   = f63_o3d0oy82l6owdiogb9dqm[13 ];
  wire wx_n37n3i1x    = f63_o3d0oy82l6owdiogb9dqm[14  ];
  wire rmydqk33eq   = f63_o3d0oy82l6owdiogb9dqm[15 ];
  wire a35tr1zbyo   = f63_o3d0oy82l6owdiogb9dqm[16 ];
  wire pzqv8u85il7   = f63_o3d0oy82l6owdiogb9dqm[17 ];
  wire ertz5b_giw  = f63_o3d0oy82l6owdiogb9dqm[18];
  wire cifajstnxdcka54  = f63_o3d0oy82l6owdiogb9dqm[19];
  wire yubia8yl4bb9c  = f63_o3d0oy82l6owdiogb9dqm[20];
  wire nvxuttrynz12  = f63_o3d0oy82l6owdiogb9dqm[21];
  wire c79vtanyxxram    = f63_o3d0oy82l6owdiogb9dqm[22  ];
  wire kv8kqf2jbw7    = f63_o3d0oy82l6owdiogb9dqm[23  ];
  wire rpacmi1zwp95    = f63_o3d0oy82l6owdiogb9dqm[24  ];
  wire gwqnhrtp4    = f63_o3d0oy82l6owdiogb9dqm[25  ];
  wire ypjg3i7dl0    = f63_o3d0oy82l6owdiogb9dqm[26  ];
  wire f0ohe956w   = f63_o3d0oy82l6owdiogb9dqm[27 ];
  wire sgrjfkl65o    = uew_1l_6faqgtso37h_zds7[5   ];
  wire dibsgfg5skf   = uew_1l_6faqgtso37h_zds7[6  ];
  wire c5lcbbkciw3vc6  = uew_1l_6faqgtso37h_zds7[7 ];
  wire zzgsxoa1dhkia   = uew_1l_6faqgtso37h_zds7[8  ];
  wire hj4cvyrejb  = uew_1l_6faqgtso37h_zds7[9 ];
  wire qe0l_afxffya5u7  = uew_1l_6faqgtso37h_zds7[10 ];
  wire z5yswe15v5    = uew_1l_6faqgtso37h_zds7[11   ];
  wire kbhyn5jnow32   = uew_1l_6faqgtso37h_zds7[12  ];
  wire qobqx6nyqpdj  = uew_1l_6faqgtso37h_zds7[13 ];
  wire aymsj4sczg   = uew_1l_6faqgtso37h_zds7[14  ];
  wire dow464urmsra  = uew_1l_6faqgtso37h_zds7[15 ];
  wire avyzty88svfq  = uew_1l_6faqgtso37h_zds7[16 ];
  wire jadgqd8db09k   = uew_1l_6faqgtso37h_zds7[17   ];
  wire u0_em9zn7vlcw  = uew_1l_6faqgtso37h_zds7[18  ];
  wire kdjefopml9bs5xby = uew_1l_6faqgtso37h_zds7[19 ];
  wire pfvv152dbk8llva  = uew_1l_6faqgtso37h_zds7[20  ];
  wire hev7phfsjoj2rx = uew_1l_6faqgtso37h_zds7[21];
  wire pf8w_s2ljvmav   = uew_1l_6faqgtso37h_zds7[22  ];
  wire gnqbx7qld2fa7g3  = uew_1l_6faqgtso37h_zds7[23 ];
  wire xfvbro69bv0tep = uew_1l_6faqgtso37h_zds7[24];
  wire go1xs0z8qd8zwe1  = uew_1l_6faqgtso37h_zds7[25 ];
  wire xjhmnd_xa2du_6g = uew_1l_6faqgtso37h_zds7[26];
  wire uq9_y2l5dw6q   = uew_1l_6faqgtso37h_zds7[27  ];
  wire nd0h5wrkl093u9  = uew_1l_6faqgtso37h_zds7[28 ];
  wire ixdkvwus8b28me = uew_1l_6faqgtso37h_zds7[29];
  wire a0mwf5tzfds7  = uew_1l_6faqgtso37h_zds7[30 ];
  wire hbtor719sgm6b1 = uew_1l_6faqgtso37h_zds7[31];
  wire ojuxyctz1rpf9   = uew_1l_6faqgtso37h_zds7[32  ];
  wire baz5vbi_zd  = uew_1l_6faqgtso37h_zds7[33 ];
  wire th_ekweb7vq1u = uew_1l_6faqgtso37h_zds7[34];
  wire dmvcpit4cpt  = uew_1l_6faqgtso37h_zds7[35 ];
  wire m8a77l1aday = uew_1l_6faqgtso37h_zds7[36];
  wire hmrx98l_nazsdh  = uew_1l_6faqgtso37h_zds7[37 ];
  wire s_s20wslhcr0ke = uew_1l_6faqgtso37h_zds7[38];
  wire ld80dv0dk64f7k_ = uew_1l_6faqgtso37h_zds7[39];
  wire yh6x5_h5s1677y = uew_1l_6faqgtso37h_zds7[40];
  wire ptn87uauvfy = uew_1l_6faqgtso37h_zds7[41];
  wire uo2vcr1g3uksaw   = uew_1l_6faqgtso37h_zds7[42  ];
  wire zd6qkrf4rnr   = uew_1l_6faqgtso37h_zds7[43  ];
  wire l30nioha_vjc   = uew_1l_6faqgtso37h_zds7[44  ];
  wire lcecqtg_qt8r   = uew_1l_6faqgtso37h_zds7[45  ];
  wire rpk5hmf4ck8wgf   = uew_1l_6faqgtso37h_zds7[46  ];
  wire ex4t35fb30  = uew_1l_6faqgtso37h_zds7[47 ];
  wire ngx30dib82    = f63_o3d0oy82l6owdiogb9dqm[28   ];
  wire t_ph70ukeyywgs   = f63_o3d0oy82l6owdiogb9dqm[29  ];
  wire px3mvn60rnd3    = f63_o3d0oy82l6owdiogb9dqm[30   ];
  wire qdsnvv2pfb   = f63_o3d0oy82l6owdiogb9dqm[31  ];
  wire fjs_jspf73t3    = f63_o3d0oy82l6owdiogb9dqm[32   ];
  wire cobog9zs7x   = f63_o3d0oy82l6owdiogb9dqm[33  ];
  wire bj_7u836    = f63_o3d0oy82l6owdiogb9dqm[34   ];
  wire ivgy7v_9d   = f63_o3d0oy82l6owdiogb9dqm[35  ];
  wire k8n93nsn    = f63_o3d0oy82l6owdiogb9dqm[36   ];
  wire cyen5b13oh4_xj   = f63_o3d0oy82l6owdiogb9dqm[37  ];
  wire q9fg5x53ud    = f63_o3d0oy82l6owdiogb9dqm[38   ];
  wire gami8f4x_a1qsq   = f63_o3d0oy82l6owdiogb9dqm[39  ];
  wire iemiml6mv3q     = f63_o3d0oy82l6owdiogb9dqm[40    ];
  wire y5gwqbpjit     = f63_o3d0oy82l6owdiogb9dqm[41    ];
  wire fydew0oon    = f63_o3d0oy82l6owdiogb9dqm[42   ];
  wire y25ionvuir_7h    = vqnbcwzo10cg732u0[95   ];
  wire os8t29xj34wk1p   = vqnbcwzo10cg732u0[96  ];
  wire ou7qpu3vjjk85    = f63_o3d0oy82l6owdiogb9dqm[43   ];
  wire b1g44t5xg   = f63_o3d0oy82l6owdiogb9dqm[44  ];
  wire v8zhxapoqe9pai  = f63_o3d0oy82l6owdiogb9dqm[45 ];
  wire mi03r0i3pb2   = f63_o3d0oy82l6owdiogb9dqm[46  ];
  wire oygn_r3rov  = f63_o3d0oy82l6owdiogb9dqm[47 ];
  wire m7m_joml4n    = f63_o3d0oy82l6owdiogb9dqm[48   ];
  wire xctdxcce22b2ol   = f63_o3d0oy82l6owdiogb9dqm[49  ];
  wire trkjd6mgoj41p  = f63_o3d0oy82l6owdiogb9dqm[50 ];
  wire yqm2e9l8qflhps   = f63_o3d0oy82l6owdiogb9dqm[51  ];
  wire cj6waeyow1  = f63_o3d0oy82l6owdiogb9dqm[52 ];
  wire xvhser      = f63_o3d0oy82l6owdiogb9dqm[53     ];
  wire edjqonhqt    = qtiogf3y1fz2gfxknzswuj[5   ];
  wire ztcp1s5cilmtw   = qtiogf3y1fz2gfxknzswuj[6  ];
  wire gupesgjbpwp5  = qtiogf3y1fz2gfxknzswuj[7 ];
  wire dxjvbl6h8ng   = qtiogf3y1fz2gfxknzswuj[8  ];
  wire t8eyqdo1vo1  = qtiogf3y1fz2gfxknzswuj[9 ];
  wire ni6p3ov9    = qtiogf3y1fz2gfxknzswuj[10   ];
  wire peb3kamgab6d   = qtiogf3y1fz2gfxknzswuj[11  ];
  wire i38hv8qg0tacqkm  = qtiogf3y1fz2gfxknzswuj[12 ];
  wire wfftg1tajppe   = qtiogf3y1fz2gfxknzswuj[13  ];
  wire vky13xw8f8jbgve  = qtiogf3y1fz2gfxknzswuj[14 ];
  wire v7ggem9i79klp1   = qtiogf3y1fz2gfxknzswuj[15   ];
  wire e4xu4gzspzdeoi  = qtiogf3y1fz2gfxknzswuj[16  ];
  wire a942bxg8vbx5s9 = qtiogf3y1fz2gfxknzswuj[17 ];
  wire zg4vqn28eg  = qtiogf3y1fz2gfxknzswuj[18  ];
  wire oaxsuvqvhxpls6h = qtiogf3y1fz2gfxknzswuj[19];
  wire vgumwbwo_6   = qtiogf3y1fz2gfxknzswuj[20  ];
  wire uzk425e3dzmu  = qtiogf3y1fz2gfxknzswuj[21 ];
  wire mngbcl1stzk7 = qtiogf3y1fz2gfxknzswuj[22];
  wire a42iwg_hdrm3vy  = qtiogf3y1fz2gfxknzswuj[23 ];
  wire vg2q1cvp3u8g = qtiogf3y1fz2gfxknzswuj[24];
  wire r1mu3vovzv0r   = qtiogf3y1fz2gfxknzswuj[25  ];
  wire h7fncem5z5x9  = qtiogf3y1fz2gfxknzswuj[26 ];
  wire y77krdi8tlj = qtiogf3y1fz2gfxknzswuj[27];
  wire qp2h493he29  = qtiogf3y1fz2gfxknzswuj[28 ];
  wire ryxvixwjxi_ub7ot = qtiogf3y1fz2gfxknzswuj[29];
  wire d1watr0ftji_r   = qtiogf3y1fz2gfxknzswuj[30  ];
  wire gum0xuidct  = qtiogf3y1fz2gfxknzswuj[31 ];
  wire er05uikr04d34ioh = qtiogf3y1fz2gfxknzswuj[32];
  wire tgrv6fv3nm45  = qtiogf3y1fz2gfxknzswuj[33 ];
  wire m30h0_l1chll9 = qtiogf3y1fz2gfxknzswuj[34];
  wire y5rwe1utr6   = qtiogf3y1fz2gfxknzswuj[35  ];
  wire ycwtj7_ux8co   = qtiogf3y1fz2gfxknzswuj[36  ];
  wire gzsw9ptxn8f   = qtiogf3y1fz2gfxknzswuj[37  ];
  wire lhtfca0wde   = qtiogf3y1fz2gfxknzswuj[38  ];
  wire yrqwiv8x45   = qtiogf3y1fz2gfxknzswuj[39  ];







  
  
  wire e03ora27k00u_e   = p4diuazqfby   | tguh9z4uqcbc; 
  wire umletcb8zgwqs  = u1mn5wzoquj0  | sudgj682o ; 
  wire iqxdtyt_g9dloiv = nn8f1wf_9ovyh | goy125ul4oyvze; 
  wire kdnn4d_qr2_jt4n3  = ye2b0mu4  | wx_n37n3i1x ; 
  wire au1gh_eazilnry  = wsflp3hzxrkbzt  | rmydqk33eq ; 
  wire svzbv80johvs = i8joes9bj | a35tr1zbyo; 

  wire k5tw9oeheqlih4   = sgrjfkl65o   | z5yswe15v5   | jadgqd8db09k  | pf8w_s2ljvmav   | uq9_y2l5dw6q  | ojuxyctz1rpf9  ; 
  wire imjs03vic384a18  = dibsgfg5skf  | kbhyn5jnow32  | u0_em9zn7vlcw | gnqbx7qld2fa7g3  | nd0h5wrkl093u9 | baz5vbi_zd ; 
  wire fsok4w6z0ij77ih = c5lcbbkciw3vc6 | qobqx6nyqpdj | kdjefopml9bs5xby| xfvbro69bv0tep | ixdkvwus8b28me| th_ekweb7vq1u; 
  wire ijnb_gpo7xg3r1  = zzgsxoa1dhkia  | aymsj4sczg  | pfvv152dbk8llva | go1xs0z8qd8zwe1  | a0mwf5tzfds7 | dmvcpit4cpt ; 
  wire ltcar0xe__n9nh61k = hj4cvyrejb  | dow464urmsra; 
  wire yed1aglcls65oj = qe0l_afxffya5u7 | avyzty88svfq | hev7phfsjoj2rx| xjhmnd_xa2du_6g | hbtor719sgm6b1| m8a77l1aday; 

  wire ijlmx1ho6tz   = edjqonhqt   | ni6p3ov9   | v7ggem9i79klp1  | vgumwbwo_6   | r1mu3vovzv0r  | d1watr0ftji_r  ; 
  wire x3e45geoeepfd_9pa  = ztcp1s5cilmtw  | peb3kamgab6d  | e4xu4gzspzdeoi | uzk425e3dzmu  | h7fncem5z5x9 | gum0xuidct ; 
  wire pvy_15wdbehc4s63n = gupesgjbpwp5 | i38hv8qg0tacqkm | a942bxg8vbx5s9| mngbcl1stzk7 | y77krdi8tlj| er05uikr04d34ioh; 
  wire azm_djrz3r5raujmu  = dxjvbl6h8ng  | wfftg1tajppe  | zg4vqn28eg | a42iwg_hdrm3vy  | qp2h493he29 | tgrv6fv3nm45 ; 
  wire sred4q00s3ugie6bhl = t8eyqdo1vo1 | vky13xw8f8jbgve | oaxsuvqvhxpls6h| vg2q1cvp3u8g | ryxvixwjxi_ub7ot| m30h0_l1chll9; 

  wire hlx2yqcuw7mugxd   = ngx30dib82  | px3mvn60rnd3 ;
  wire gjgqa949f4epnz  = t_ph70ukeyywgs | qdsnvv2pfb;

  wire n0uej4ag_la   = fjs_jspf73t3  | k8n93nsn ;
  wire jcv5t8qp92n4yn_  = cobog9zs7x | cyen5b13oh4_xj;
  wire u340gmafpm_q0kft   = bj_7u836  | q9fg5x53ud ;
  wire u4kt5axdfc1f  = ivgy7v_9d | gami8f4x_a1qsq;

  wire lwh7ejgwbe0y3xd6   = ou7qpu3vjjk85   | m7m_joml4n  ; 
  wire e6mszw3shdp5  = b1g44t5xg  | xctdxcce22b2ol ; 
  wire p1b08_so0a9eejxiuw = v8zhxapoqe9pai | trkjd6mgoj41p; 
  wire h_u6dnfrybg78e0tn  = mi03r0i3pb2  | yqm2e9l8qflhps ; 
  wire i7uc6ffwjktqvuq4q6 = oygn_r3rov | cj6waeyow1; 

  wire tmrmbibjnw  = yubia8yl4bb9c | nvxuttrynz12 | ertz5b_giw | cifajstnxdcka54 ;
  wire yl7v16qdbo3u7 = yh6x5_h5s1677y | ptn87uauvfy | s_s20wslhcr0ke | ld80dv0dk64f7k_;
  wire g8dm1b58pm6xt = pzqv8u85il7| nvxuttrynz12| cifajstnxdcka54 | hmrx98l_nazsdh| ptn87uauvfy| ld80dv0dk64f7k_;

  wire cr75ulfp     =  tmrmbibjnw | yl7v16qdbo3u7 | g8dm1b58pm6xt;
  wire c9hqqulyow5pvq  = rpacmi1zwp95  | gwqnhrtp4   | c79vtanyxxram   | kv8kqf2jbw7 ; 
  wire g2s8ge1hum_lb = l30nioha_vjc | lcecqtg_qt8r  | uo2vcr1g3uksaw  | zd6qkrf4rnr;
  wire brrzcx4c49ey = iemiml6mv3q | y5gwqbpjit;
  wire pmct0ov7_sv0 = gzsw9ptxn8f | lhtfca0wde  | y5rwe1utr6  | ycwtj7_ux8co;
  wire jpt8d5z4s = c9hqqulyow5pvq | g2s8ge1hum_lb | brrzcx4c49ey | pmct0ov7_sv0;

  wire gv93tjc7rha = ypjg3i7dl0 | f0ohe956w | rpk5hmf4ck8wgf | ex4t35fb30 | fydew0oon | yrqwiv8x45;
 
  wire h0xl_5 = y25ionvuir_7h | os8t29xj34wk1p;


  
  
  wire b5rzoldza22sb  = p4diuazqfby | u1mn5wzoquj0  | ye2b0mu4 |  wsflp3hzxrkbzt;
  wire lqhl5nqoq7lfmc  = nn8f1wf_9ovyh | i8joes9bj;
  wire aeaere3i7e23 = b5rzoldza22sb | lqhl5nqoq7lfmc;

  wire ry_xj_27plplx1 = sgrjfkl65o | dibsgfg5skf | zzgsxoa1dhkia | hj4cvyrejb;
  wire xaabzrcv_raxz = c5lcbbkciw3vc6 | qe0l_afxffya5u7;
  wire d5rqmmzhqlmo9g_c = ry_xj_27plplx1 | xaabzrcv_raxz;
  
  wire q1yh6x8lrrng = edjqonhqt | ztcp1s5cilmtw | dxjvbl6h8ng;
  wire tqciamxv2cnjc = gupesgjbpwp5 | t8eyqdo1vo1;
  wire ogjz62jz907v2 = q1yh6x8lrrng | tqciamxv2cnjc;

  wire puthzl6v_gagc37  = ngx30dib82 ;
  wire ndjzhv18pdknqdg  = t_ph70ukeyywgs;
  wire x06kbvmm_1ew  = puthzl6v_gagc37 | ndjzhv18pdknqdg;

  wire zopjtkfsisw  = fjs_jspf73t3 |  bj_7u836  ;
  wire gj5vh6m57syo6u  = cobog9zs7x |  ivgy7v_9d;
  wire uqc77d2rlan5  = zopjtkfsisw | gj5vh6m57syo6u;

  wire g1v10rklyrj1l81hm = ou7qpu3vjjk85   | b1g44t5xg  | mi03r0i3pb2 ;
  wire rzd2hcw89e200ggc = v8zhxapoqe9pai | oygn_r3rov ;
  wire sw42pegskxo1j = g1v10rklyrj1l81hm | rzd2hcw89e200ggc ; 

  wire ehxjmrr4a83haci0 = jadgqd8db09k | u0_em9zn7vlcw | pfvv152dbk8llva ;
  wire uiuqumf3h3juzv_rner = kdjefopml9bs5xby | hev7phfsjoj2rx;
  wire a6bi_6k_4l8jx17e5 = ehxjmrr4a83haci0 | uiuqumf3h3juzv_rner;

  wire p5bi0utoyxujnli = pf8w_s2ljvmav | gnqbx7qld2fa7g3 | go1xs0z8qd8zwe1 ;
  wire j7pgmypqwndz232ey3 = xfvbro69bv0tep | xjhmnd_xa2du_6g;
  wire z42jii1vw3c1ys2x = p5bi0utoyxujnli | j7pgmypqwndz232ey3;

  wire fu3jigjcdxom_x  = uq9_y2l5dw6q | nd0h5wrkl093u9| a0mwf5tzfds7;
  wire aiphwaji28ool7  = ixdkvwus8b28me | hbtor719sgm6b1;
  wire roujn5dz1r9vfxa2  = fu3jigjcdxom_x | aiphwaji28ool7;

  wire p8hb0e1kz7_wj0  = ojuxyctz1rpf9 | baz5vbi_zd | dmvcpit4cpt;
  wire evgs_c8j8lssbfa1  = th_ekweb7vq1u | m8a77l1aday;
  wire t03c5iq5nxjj17dgf  = p8hb0e1kz7_wj0 | evgs_c8j8lssbfa1;
  
  wire mid3yvd1dc5p_3 = v7ggem9i79klp1 | e4xu4gzspzdeoi | zg4vqn28eg ;
  wire d33k1t15iao77sn8eq = a942bxg8vbx5s9 | oaxsuvqvhxpls6h;
  wire mr6gygq2r8eshp2cj = mid3yvd1dc5p_3 | d33k1t15iao77sn8eq;

  wire nhk0haqb79ub07mq2b = vgumwbwo_6 | uzk425e3dzmu | a42iwg_hdrm3vy ;
  wire ghwvor5rmxzau7tznu = mngbcl1stzk7 | vg2q1cvp3u8g;
  wire insn017okyfbloukc = nhk0haqb79ub07mq2b | ghwvor5rmxzau7tznu;

  wire ocl0e6_c3wncrmc6  = r1mu3vovzv0r | h7fncem5z5x9| qp2h493he29;
  wire qtw5zaawn8u4jd9dy  = y77krdi8tlj | ryxvixwjxi_ub7ot;
  wire oo3l5yfmx2itl  = ocl0e6_c3wncrmc6 | qtw5zaawn8u4jd9dy;

  wire bsi917d7yfryhti9  = d1watr0ftji_r | gum0xuidct | tgrv6fv3nm45;
  wire egbv5yccd8p4nkls  = er05uikr04d34ioh | m30h0_l1chll9;
  wire ilh98i86sgjp7  = bsi917d7yfryhti9 | egbv5yccd8p4nkls;

  wire y5fcft2979miyo = tguh9z4uqcbc   | sudgj682o  | wx_n37n3i1x | rmydqk33eq | ertz5b_giw | cifajstnxdcka54 | kv8kqf2jbw7 | c79vtanyxxram;
  wire ovpxn8hcr5sg7gu = goy125ul4oyvze | a35tr1zbyo | yubia8yl4bb9c | nvxuttrynz12 | gwqnhrtp4 | rpacmi1zwp95 | h0xl_5;
  wire dpfu5qbd2ew5mxu = y5fcft2979miyo | ovpxn8hcr5sg7gu ;
  
  wire e10mbsw7wquig = z5yswe15v5 | kbhyn5jnow32 |  aymsj4sczg | dow464urmsra | s_s20wslhcr0ke | ld80dv0dk64f7k_ | zd6qkrf4rnr | uo2vcr1g3uksaw;
  wire mmo5t4gqbmx0 = qobqx6nyqpdj | avyzty88svfq | yh6x5_h5s1677y | ptn87uauvfy | lcecqtg_qt8r | l30nioha_vjc ;
  wire fs5ihva8cewrcc5j = e10mbsw7wquig | mmo5t4gqbmx0;
  
  wire h2ip0rex3tgx3 = ni6p3ov9 | peb3kamgab6d |  wfftg1tajppe |  ycwtj7_ux8co | y5rwe1utr6;
  wire ik95b3bzb6651bvr = i38hv8qg0tacqkm | vky13xw8f8jbgve |  lhtfca0wde | gzsw9ptxn8f ;
  wire da00qq0n3p6f35f = h2ip0rex3tgx3 | ik95b3bzb6651bvr;

  wire lmqvm9loqx5tiub =  px3mvn60rnd3  ;
  wire arkju513nouw =  qdsnvv2pfb ;
  wire cxmega4p8g =  lmqvm9loqx5tiub | arkju513nouw ;

  wire gm1n06hqq92sw4_ = q9fg5x53ud  | k8n93nsn | brrzcx4c49ey;
  wire zzh_n0oxtxd6zi = gami8f4x_a1qsq | cyen5b13oh4_xj;
  wire exl_abiv15e = gm1n06hqq92sw4_ | zzh_n0oxtxd6zi;

  wire dfcpt8muurpn6 = m7m_joml4n   | xctdxcce22b2ol  | yqm2e9l8qflhps ;
  wire lzu7zvw68i3ihdsw = trkjd6mgoj41p | cj6waeyow1 ;
  wire gtp49bjcaikct_5 = dfcpt8muurpn6 | lzu7zvw68i3ihdsw ;
  wire a4398r0pvs = sw42pegskxo1j | gtp49bjcaikct_5; 

  
  
  wire mf5fcnu2azr = aeaere3i7e23 | d5rqmmzhqlmo9g_c | z42jii1vw3c1ys2x | t03c5iq5nxjj17dgf |
                x06kbvmm_1ew | uqc77d2rlan5 | gv93tjc7rha | sw42pegskxo1j | xvhser | ogjz62jz907v2
                | insn017okyfbloukc | ilh98i86sgjp7;

  wire m0mq6jm4ys = dpfu5qbd2ew5mxu | fs5ihva8cewrcc5j | a6bi_6k_4l8jx17e5 | roujn5dz1r9vfxa2 |
                cxmega4p8g | exl_abiv15e | gtp49bjcaikct_5 | da00qq0n3p6f35f 
                | mr6gygq2r8eshp2cj | oo3l5yfmx2itl;

  wire [64-1:0] yxz3vex1f   = m35ros_bzlaqo8y319z  ;
  wire [64-1:0] afthitl2   = uq5g_s44gt3h0fbg4zzv  ;
  wire [64-1:0] tz6u29u8fwu9n_i = i8whgk1t5jsbvv8u3ojllu7;
  wire [64-1:0] s_0mxmrxstpu = c7cw30bh940izgc1knsjmx;

  
  

  wire[7:0] mfqlkqsfqqtr7aq3 = yxz3vex1f[63:56];  
  wire[7:0] c855qo4w5w6shr01k = yxz3vex1f[55:48];
  wire[7:0] tlqrl7o_ea5f7jvuz = yxz3vex1f[47:40];
  wire[7:0] za_gepbwiydx41hlau = yxz3vex1f[39:32];
  wire[7:0] bdaw595w6ylh6t3 = yxz3vex1f[31:24];  
  wire[7:0] kmxpyw7wqu2t_gzzj = yxz3vex1f[23:16];
  wire[7:0] io2x7wr4ojvgigpt = yxz3vex1f[15:8 ];
  wire[7:0] l0vwpa90rm8y_ronbdy = yxz3vex1f[7 :0 ];
  wire[7:0] qea_ieqiyamdyl4a_r = ~mfqlkqsfqqtr7aq3;  
  wire[7:0] m5mvfvapj5hwubsq24t32h9 = ~c855qo4w5w6shr01k;
  wire[7:0] qy46f8x2_p9_avu_yxk = ~tlqrl7o_ea5f7jvuz;
  wire[7:0] k6a5b9u9o5e5e2zt_p = ~za_gepbwiydx41hlau;
  wire[7:0] xgevy4awjdswvvqc1g9ie2 = ~bdaw595w6ylh6t3;  
  wire[7:0] n8kxu2euntozsbkacz = ~kmxpyw7wqu2t_gzzj;
  wire[7:0] tp2kk00j9852eqxln2 = ~io2x7wr4ojvgigpt;
  wire[7:0] i9yvzlsza1100l33ahy2 = ~l0vwpa90rm8y_ronbdy;
  wire u67ocgqs0ji6 = mfqlkqsfqqtr7aq3[7];
  wire fytthe9rcpw = c855qo4w5w6shr01k[7];
  wire hfuuhnhjjbzyhr = tlqrl7o_ea5f7jvuz[7];
  wire rhmxsn4ow99l3 = za_gepbwiydx41hlau[7];
  wire tj0mpvq6bvwu = bdaw595w6ylh6t3[7];
  wire s28zkzzcmxybp8mt = kmxpyw7wqu2t_gzzj[7];
  wire jxmxj59r3yqcgf5z = io2x7wr4ojvgigpt[7];
  wire apwk5icq9cv = l0vwpa90rm8y_ronbdy[7];
  wire ypuadjidxyfdybfwgl9 = qea_ieqiyamdyl4a_r[7];
  wire h36daabl2rsl0tsr43y = m5mvfvapj5hwubsq24t32h9[7];
  wire t1e0bugyoi597hx24 = qy46f8x2_p9_avu_yxk[7];
  wire zy9qt1dks5iib9vehzdf = k6a5b9u9o5e5e2zt_p[7];
  wire vli_9lhakwcu7im3ji6l = xgevy4awjdswvvqc1g9ie2[7];
  wire f4zi2kui0ji6s9fv = n8kxu2euntozsbkacz[7];
  wire fppmy95e8mpnbiby8 = tp2kk00j9852eqxln2[7];
  wire efn1_uky5_l91c_62t = i9yvzlsza1100l33ahy2[7];
  wire[15:0] ug44br6vqgrl = {mfqlkqsfqqtr7aq3,c855qo4w5w6shr01k};  
  wire[15:0] z9tavnbfnm_4 = {tlqrl7o_ea5f7jvuz,za_gepbwiydx41hlau};
  wire[15:0] qurlzg4fi3qln = {bdaw595w6ylh6t3,kmxpyw7wqu2t_gzzj};
  wire[15:0] uydrrfewr6ksaehu = {io2x7wr4ojvgigpt,l0vwpa90rm8y_ronbdy};
  wire[15:0] nvlpyddg1wr2om4m12i = {qea_ieqiyamdyl4a_r,m5mvfvapj5hwubsq24t32h9};  
  wire[15:0] pg762iiol2fljfgvqmzs = {qy46f8x2_p9_avu_yxk,k6a5b9u9o5e5e2zt_p};
  wire[15:0] zk_53533f4oe6mmptg = {xgevy4awjdswvvqc1g9ie2,n8kxu2euntozsbkacz};
  wire[15:0] wwx8k3mblud3m1eg_y = {tp2kk00j9852eqxln2,i9yvzlsza1100l33ahy2};
  
  wire[31:0] b_xqc3mgz11e = {ug44br6vqgrl,z9tavnbfnm_4};
  wire[31:0] x4vwdbhy47grdx6 = {qurlzg4fi3qln,uydrrfewr6ksaehu};
  wire[31:0] y7rms3iwbod90teylc90 = {nvlpyddg1wr2om4m12i,pg762iiol2fljfgvqmzs};
  wire[31:0] dlq8_mc8wk9ae8tp = {zk_53533f4oe6mmptg,wwx8k3mblud3m1eg_y};

    wire [80-1:0] g0aqd08ou7rfnv3ndp =
      ({80{b5rzoldza22sb}} & {1'b0,u67ocgqs0ji6,mfqlkqsfqqtr7aq3,1'b0,fytthe9rcpw,c855qo4w5w6shr01k,
                                               1'b0,hfuuhnhjjbzyhr,tlqrl7o_ea5f7jvuz,1'b0,rhmxsn4ow99l3,za_gepbwiydx41hlau,   
                                               1'b0,tj0mpvq6bvwu,bdaw595w6ylh6t3,1'b0,s28zkzzcmxybp8mt,kmxpyw7wqu2t_gzzj,  
                                               1'b0,jxmxj59r3yqcgf5z,io2x7wr4ojvgigpt,1'b0,apwk5icq9cv,l0vwpa90rm8y_ronbdy})  
    | ({80{lqhl5nqoq7lfmc}} & {2'b00,mfqlkqsfqqtr7aq3, 2'b00,c855qo4w5w6shr01k, 2'b00,tlqrl7o_ea5f7jvuz, 2'b00,za_gepbwiydx41hlau,  
                                               2'b00,bdaw595w6ylh6t3, 2'b00,kmxpyw7wqu2t_gzzj, 2'b00,io2x7wr4ojvgigpt, 2'b00,l0vwpa90rm8y_ronbdy})  
    | ({80{y5fcft2979miyo}} & {1'b0,u67ocgqs0ji6,mfqlkqsfqqtr7aq3,1'b1,fytthe9rcpw,c855qo4w5w6shr01k,
                                               1'b1,hfuuhnhjjbzyhr,tlqrl7o_ea5f7jvuz,1'b1,rhmxsn4ow99l3,za_gepbwiydx41hlau,
                                               1'b1,tj0mpvq6bvwu,bdaw595w6ylh6t3,1'b1,s28zkzzcmxybp8mt,kmxpyw7wqu2t_gzzj,
                                               1'b1,jxmxj59r3yqcgf5z,io2x7wr4ojvgigpt,1'b1,apwk5icq9cv,l0vwpa90rm8y_ronbdy}) 
    | ({80{ovpxn8hcr5sg7gu }} & {2'b00,mfqlkqsfqqtr7aq3, 2'b10,c855qo4w5w6shr01k, 2'b10,tlqrl7o_ea5f7jvuz, 2'b10,za_gepbwiydx41hlau,
                                                2'b10,bdaw595w6ylh6t3, 2'b10,kmxpyw7wqu2t_gzzj, 2'b10,io2x7wr4ojvgigpt, 2'b10,l0vwpa90rm8y_ronbdy}) 
    | ({80{ypjg3i7dl0 | f0ohe956w}} 
                                                 & {2'b00,mfqlkqsfqqtr7aq3, 2'b00,c855qo4w5w6shr01k, 2'b00,tlqrl7o_ea5f7jvuz, 2'b00,za_gepbwiydx41hlau,
                                                    2'b00,bdaw595w6ylh6t3, 2'b00,kmxpyw7wqu2t_gzzj, 2'b00,io2x7wr4ojvgigpt, 2'b00,l0vwpa90rm8y_ronbdy}) 
    | ({80{ry_xj_27plplx1 }}
                                            & {3'b000, u67ocgqs0ji6, ug44br6vqgrl,  3'b000, hfuuhnhjjbzyhr, z9tavnbfnm_4,   
                                              3'b000, tj0mpvq6bvwu, qurlzg4fi3qln,  3'b000, jxmxj59r3yqcgf5z, uydrrfewr6ksaehu})  
    | ({80{ehxjmrr4a83haci0 | fu3jigjcdxom_x}}
                                            & {3'b000, u67ocgqs0ji6, ug44br6vqgrl,  3'b000, hfuuhnhjjbzyhr, z9tavnbfnm_4,   
                                               3'b100, tj0mpvq6bvwu, qurlzg4fi3qln,  3'b000, jxmxj59r3yqcgf5z, uydrrfewr6ksaehu})  
    | ({80{xaabzrcv_raxz }}
                                            & {4'h0,ug44br6vqgrl, 4'h0,z9tavnbfnm_4, 4'h0,qurlzg4fi3qln, 4'h0,uydrrfewr6ksaehu})  
    | ({80{uiuqumf3h3juzv_rner | aiphwaji28ool7}}
                                            & {4'b0000,ug44br6vqgrl, 4'b0000,z9tavnbfnm_4, 4'b1000,qurlzg4fi3qln, 4'b0000,uydrrfewr6ksaehu})  
    | ({80{rpk5hmf4ck8wgf | ex4t35fb30}}
                                            & {4'h0,ug44br6vqgrl, 4'h0,z9tavnbfnm_4, 4'h0,qurlzg4fi3qln, 4'h0,uydrrfewr6ksaehu})  
    | ({80{e10mbsw7wquig}}
                                            & {3'b000,u67ocgqs0ji6, ug44br6vqgrl, 3'b100,hfuuhnhjjbzyhr, z9tavnbfnm_4, 
                                               3'b100,tj0mpvq6bvwu, qurlzg4fi3qln, 3'b100,jxmxj59r3yqcgf5z, uydrrfewr6ksaehu}) 
    | ({80{p5bi0utoyxujnli | p8hb0e1kz7_wj0}}
                                            & {3'b000,u67ocgqs0ji6, ug44br6vqgrl, 3'b100,hfuuhnhjjbzyhr, z9tavnbfnm_4, 
                                               3'b000,tj0mpvq6bvwu, qurlzg4fi3qln, 3'b100,jxmxj59r3yqcgf5z, uydrrfewr6ksaehu}) 
    | ({80{mmo5t4gqbmx0 }}
                                            & {4'b0000,ug44br6vqgrl, 4'b1000,z9tavnbfnm_4, 4'b1000,qurlzg4fi3qln, 4'b1000,uydrrfewr6ksaehu}) 
    | ({80{j7pgmypqwndz232ey3 | evgs_c8j8lssbfa1}}
                                            & {4'b0000,ug44br6vqgrl, 4'b1000,z9tavnbfnm_4, 4'b0000,qurlzg4fi3qln, 4'b1000,uydrrfewr6ksaehu}) 
    | ({80{(puthzl6v_gagc37 | zopjtkfsisw | lmqvm9loqx5tiub | gm1n06hqq92sw4_ )}} 
                                                 & {47'b0,tj0mpvq6bvwu, qurlzg4fi3qln, uydrrfewr6ksaehu}) 
    | ({80{(ndjzhv18pdknqdg | gj5vh6m57syo6u | arkju513nouw | zzh_n0oxtxd6zi | fydew0oon)}}
                                                 & {48'b0,qurlzg4fi3qln, uydrrfewr6ksaehu})  
    | ({80{(g1v10rklyrj1l81hm | dfcpt8muurpn6 | xvhser)}} 
                                                 & {15'b0,u67ocgqs0ji6,yxz3vex1f})
    | ({80{(rzd2hcw89e200ggc | lzu7zvw68i3ihdsw)}} 
                                                 & {16'b0,yxz3vex1f})
    
    | ({80{q1yh6x8lrrng }} & {7'b000, u67ocgqs0ji6, b_xqc3mgz11e,  7'h00, tj0mpvq6bvwu, x4vwdbhy47grdx6})  
    | ({80{mid3yvd1dc5p_3 | ocl0e6_c3wncrmc6}}
                                              & {7'b000, u67ocgqs0ji6, b_xqc3mgz11e,  7'h00, tj0mpvq6bvwu, x4vwdbhy47grdx6})  
    | ({80{tqciamxv2cnjc }} & {8'h00,b_xqc3mgz11e, 8'h00,x4vwdbhy47grdx6})  
    | ({80{d33k1t15iao77sn8eq | qtw5zaawn8u4jd9dy}}
                                              & {8'h00, b_xqc3mgz11e, 8'h00, x4vwdbhy47grdx6})  
    | ({80{yrqwiv8x45}}  & {8'h00, b_xqc3mgz11e, 8'h00, x4vwdbhy47grdx6})  
    | ({80{h2ip0rex3tgx3}}
                                            & {7'h00, u67ocgqs0ji6, b_xqc3mgz11e, 7'h40, tj0mpvq6bvwu, x4vwdbhy47grdx6}) 
    | ({80{nhk0haqb79ub07mq2b | bsi917d7yfryhti9}}
                                            & {7'h00, u67ocgqs0ji6, b_xqc3mgz11e, 7'h40, tj0mpvq6bvwu, x4vwdbhy47grdx6}) 
    | ({80{ik95b3bzb6651bvr }}
                                            & {8'h00, b_xqc3mgz11e, 8'h80, x4vwdbhy47grdx6}) 
    | ({80{ghwvor5rmxzau7tznu | egbv5yccd8p4nkls}}
                                            & {8'h00, b_xqc3mgz11e, 8'h80, x4vwdbhy47grdx6}) 
    ;
  wire[7:0] tw9ki934xehoq8 = afthitl2[63:56];  
  wire[7:0] q9cii0knfkzpzmo = afthitl2[55:48];
  wire[7:0] s8amssre_wgztttyk = afthitl2[47:40];
  wire[7:0] oip62i3gqus90p3_ = afthitl2[39:32];
  wire[7:0] mkdo3k6oahvj1wx = afthitl2[31:24];  
  wire[7:0] f6kvbyx3whxntsm = afthitl2[23:16];
  wire[7:0] oavwfeahe75zx1l = afthitl2[15:8 ];
  wire[7:0] p0uj0k3yvjy98a28 = afthitl2[7 :0 ];
  wire[7:0] w20x495cbb7i388wgks = ~tw9ki934xehoq8;  
  wire[7:0] kr_yb61rfnwwd4151olf = ~q9cii0knfkzpzmo;
  wire[7:0] mrq19_szsu3twjbvdxybs = ~s8amssre_wgztttyk;
  wire[7:0] spntsnggyob6ibh46b = ~oip62i3gqus90p3_;
  wire[7:0] a28dfvr46yscpsxxrqas = ~mkdo3k6oahvj1wx;  
  wire[7:0] frfa1tkv3o5jto1_rx = ~f6kvbyx3whxntsm;
  wire[7:0] nstrhjdlr5f4u5l6j98e = ~oavwfeahe75zx1l;
  wire[7:0] e4e1zt1mv_7awhuytdi51fg = ~p0uj0k3yvjy98a28;
  wire cbzbmu27xirmn = tw9ki934xehoq8[7];
  wire dyw_n7no3f2_x = q9cii0knfkzpzmo[7];
  wire ldm4_5itwcwe_bp = s8amssre_wgztttyk[7];
  wire l3p4ad20uuokz = oip62i3gqus90p3_[7];
  wire dbezizgky8oe_1s = mkdo3k6oahvj1wx[7];
  wire hx5mapiqg5pmw = f6kvbyx3whxntsm[7];
  wire pn8lwvdt87m = oavwfeahe75zx1l[7];
  wire ppmpgu269l3ge4_e = p0uj0k3yvjy98a28[7];
  wire qy4465l158u4avl1st = w20x495cbb7i388wgks[7];
  wire akl056wm04gojrqnu = kr_yb61rfnwwd4151olf[7];
  wire gb3vkwmv5r_y65x7u = mrq19_szsu3twjbvdxybs[7];
  wire tpfl0ae8soivk66ff6 = spntsnggyob6ibh46b[7];
  wire zlhgyh5dfmt_aom = a28dfvr46yscpsxxrqas[7];
  wire qw4mdq7ebl14308ui = frfa1tkv3o5jto1_rx[7];
  wire s0kk19tok_qxdimmy = nstrhjdlr5f4u5l6j98e[7];
  wire jj9veqnp7ig8m6_4uk1 = e4e1zt1mv_7awhuytdi51fg[7];
  wire[15:0] jq5vss15lef0fq = {tw9ki934xehoq8,q9cii0knfkzpzmo};  
  wire[15:0] vi_9c4xfw3laf = {s8amssre_wgztttyk,oip62i3gqus90p3_};
  wire[15:0] s_jnoaq4rvg2k5qk = {mkdo3k6oahvj1wx,f6kvbyx3whxntsm};
  wire[15:0] ighridqr233htz = {oavwfeahe75zx1l,p0uj0k3yvjy98a28};
  wire[15:0] d19dz7sd0y4n14u7q2iiu = {w20x495cbb7i388wgks,kr_yb61rfnwwd4151olf};  
  wire[15:0] o3odbzchqomo1ykxtvrfo = {mrq19_szsu3twjbvdxybs,spntsnggyob6ibh46b};
  wire[15:0] xb9ns8h_licc_3r22el = {a28dfvr46yscpsxxrqas,frfa1tkv3o5jto1_rx};
  wire[15:0] zmuacjwbp82p1iy9_f = {nstrhjdlr5f4u5l6j98e,e4e1zt1mv_7awhuytdi51fg};

  wire[31:0] bw3242dwyw8g = {jq5vss15lef0fq,vi_9c4xfw3laf};
  wire[31:0] is0m6qik1xe3onr0 = {s_jnoaq4rvg2k5qk,ighridqr233htz};
  wire[31:0] jsfb7rigmw_f0kn1qye3 = {d19dz7sd0y4n14u7q2iiu,o3odbzchqomo1ykxtvrfo};
  wire[31:0] jm_j4gy26gvwm99in = {xb9ns8h_licc_3r22el,zmuacjwbp82p1iy9_f};



    wire [80-1:0] ccbzdmuytukdpcsy26d =
        ({80{b5rzoldza22sb}} & {1'b0,cbzbmu27xirmn,tw9ki934xehoq8,  1'b0,dyw_n7no3f2_x,q9cii0knfkzpzmo,
                                                 1'b0,ldm4_5itwcwe_bp,s8amssre_wgztttyk,  1'b0,l3p4ad20uuokz,oip62i3gqus90p3_, 
                                                 1'b0,dbezizgky8oe_1s,mkdo3k6oahvj1wx,  1'b0,hx5mapiqg5pmw,f6kvbyx3whxntsm,
                                                 1'b0,pn8lwvdt87m,oavwfeahe75zx1l,  1'b0,ppmpgu269l3ge4_e,p0uj0k3yvjy98a28}) 
      | ({80{lqhl5nqoq7lfmc}} & {2'b00,tw9ki934xehoq8, 2'b00,q9cii0knfkzpzmo, 2'b00,s8amssre_wgztttyk, 2'b00,oip62i3gqus90p3_,  
                                                 2'b00,mkdo3k6oahvj1wx, 2'b00,f6kvbyx3whxntsm, 2'b00,oavwfeahe75zx1l, 2'b00,p0uj0k3yvjy98a28})  
      | ({80{y5fcft2979miyo}} & {1'b0,qy4465l158u4avl1st,w20x495cbb7i388wgks,  1'b1,akl056wm04gojrqnu,kr_yb61rfnwwd4151olf,
                                                 1'b1,gb3vkwmv5r_y65x7u,mrq19_szsu3twjbvdxybs,  1'b1,tpfl0ae8soivk66ff6,spntsnggyob6ibh46b,   
                                                 1'b1,zlhgyh5dfmt_aom,a28dfvr46yscpsxxrqas,  1'b1,qw4mdq7ebl14308ui,frfa1tkv3o5jto1_rx,
                                                 1'b1,s0kk19tok_qxdimmy,nstrhjdlr5f4u5l6j98e,  1'b1,jj9veqnp7ig8m6_4uk1,e4e1zt1mv_7awhuytdi51fg})  
      | ({80{ovpxn8hcr5sg7gu}} & {2'b01,w20x495cbb7i388wgks,2'b11,kr_yb61rfnwwd4151olf,2'b11,mrq19_szsu3twjbvdxybs,2'b11,spntsnggyob6ibh46b,  
                                                 2'b11,a28dfvr46yscpsxxrqas,2'b11,frfa1tkv3o5jto1_rx,2'b11,nstrhjdlr5f4u5l6j98e,2'b11,e4e1zt1mv_7awhuytdi51fg}) 
      | ({80{ry_xj_27plplx1  }} & {3'b000 , cbzbmu27xirmn,jq5vss15lef0fq, 3'b000 , ldm4_5itwcwe_bp,vi_9c4xfw3laf, 
                                                    3'b000 , dbezizgky8oe_1s,s_jnoaq4rvg2k5qk, 3'b000 , pn8lwvdt87m,ighridqr233htz}) 
      | ({80{xaabzrcv_raxz  }} & {4'b0000,jq5vss15lef0fq,4'b0000, vi_9c4xfw3laf, 4'b0000, s_jnoaq4rvg2k5qk,4'b0000, ighridqr233htz})
      | ({80{e10mbsw7wquig  }} & {3'b000 ,qy4465l158u4avl1st,d19dz7sd0y4n14u7q2iiu, 3'b100 ,gb3vkwmv5r_y65x7u,o3odbzchqomo1ykxtvrfo, 
                                                    3'b100 ,zlhgyh5dfmt_aom,xb9ns8h_licc_3r22el, 3'b100 ,s0kk19tok_qxdimmy,zmuacjwbp82p1iy9_f}) 
      | ({80{mmo5t4gqbmx0  }} & {4'b0001,d19dz7sd0y4n14u7q2iiu, 4'b1001,o3odbzchqomo1ykxtvrfo, 4'b1001,xb9ns8h_licc_3r22el, 4'b1001,zmuacjwbp82p1iy9_f})
      | ({80{ehxjmrr4a83haci0}} & {3'b000 ,ldm4_5itwcwe_bp, vi_9c4xfw3laf, 3'b000 ,qy4465l158u4avl1st, d19dz7sd0y4n14u7q2iiu,  
                                                    3'b100 ,pn8lwvdt87m, ighridqr233htz, 3'b000 ,zlhgyh5dfmt_aom, xb9ns8h_licc_3r22el}) 
      | ({80{uiuqumf3h3juzv_rner}} & {4'b0000,vi_9c4xfw3laf, 4'b0001,d19dz7sd0y4n14u7q2iiu, 4'b1000,ighridqr233htz, 4'b0001,xb9ns8h_licc_3r22el}) 
      | ({80{p5bi0utoyxujnli}} & {3'b000 ,gb3vkwmv5r_y65x7u, o3odbzchqomo1ykxtvrfo, 3'b100 , cbzbmu27xirmn,jq5vss15lef0fq,   
                                                    3'b000 ,s0kk19tok_qxdimmy, zmuacjwbp82p1iy9_f, 3'b100 , dbezizgky8oe_1s,s_jnoaq4rvg2k5qk}) 
      | ({80{j7pgmypqwndz232ey3}} & {4'b0001,o3odbzchqomo1ykxtvrfo,4'b1000, jq5vss15lef0fq, 4'b0001,zmuacjwbp82p1iy9_f,4'b1000, s_jnoaq4rvg2k5qk}) 
      | ({80{fu3jigjcdxom_x }} & {3'b000 ,cbzbmu27xirmn,jq5vss15lef0fq, 3'b000, gb3vkwmv5r_y65x7u, o3odbzchqomo1ykxtvrfo,
                                                    3'b100 ,dbezizgky8oe_1s,s_jnoaq4rvg2k5qk, 3'b000, s0kk19tok_qxdimmy, zmuacjwbp82p1iy9_f}) 
      | ({80{aiphwaji28ool7 }} & {4'b0000,jq5vss15lef0fq,  4'b0001,o3odbzchqomo1ykxtvrfo, 4'b1000,s_jnoaq4rvg2k5qk,  4'b0001,zmuacjwbp82p1iy9_f}) 
      | ({80{p8hb0e1kz7_wj0 }} & {3'b000 ,qy4465l158u4avl1st, d19dz7sd0y4n14u7q2iiu,  3'b100 ,  ldm4_5itwcwe_bp,vi_9c4xfw3laf, 
                                                    3'b000 ,zlhgyh5dfmt_aom, xb9ns8h_licc_3r22el,  3'b100 ,  pn8lwvdt87m,ighridqr233htz}) 
      | ({80{evgs_c8j8lssbfa1 }} & {4'b0001,d19dz7sd0y4n14u7q2iiu, 4'b1000,vi_9c4xfw3laf,  4'b0001,xb9ns8h_licc_3r22el, 4'b1000,ighridqr233htz}) 
      | ({80{(puthzl6v_gagc37 | zopjtkfsisw)}} & {47'b0,dbezizgky8oe_1s,s_jnoaq4rvg2k5qk,ighridqr233htz}) 
      | ({80{(ndjzhv18pdknqdg | gj5vh6m57syo6u)}} & {48'b0,s_jnoaq4rvg2k5qk,ighridqr233htz})
      | ({80{(lmqvm9loqx5tiub | gm1n06hqq92sw4_)}} & {47'b0,zlhgyh5dfmt_aom,xb9ns8h_licc_3r22el,zmuacjwbp82p1iy9_f}) 
      | ({80{(arkju513nouw | zzh_n0oxtxd6zi)}} & {48'h1,xb9ns8h_licc_3r22el,zmuacjwbp82p1iy9_f}) 
         
      | ({80{ypjg3i7dl0 | f0ohe956w}}   & {2'b0,{8{u67ocgqs0ji6}},2'b0,{8{fytthe9rcpw}},2'b0,{8{hfuuhnhjjbzyhr}},2'b0,{8{rhmxsn4ow99l3}}, 
                                                            2'b0,{8{tj0mpvq6bvwu}},2'b0,{8{s28zkzzcmxybp8mt}},2'b0,{8{jxmxj59r3yqcgf5z}},2'b0,{8{apwk5icq9cv}}}) 
      | ({80{rpk5hmf4ck8wgf | ex4t35fb30}} & {4'b000,{16{u67ocgqs0ji6}},4'b0000,{16{hfuuhnhjjbzyhr}},  
                                                            4'b000,{16{tj0mpvq6bvwu}},4'b0000,{16{jxmxj59r3yqcgf5z}}}) 
      | ({80{fydew0oon}}  & {48'b0,{32{yxz3vex1f[31]}}}) 
      | ({80{(g1v10rklyrj1l81hm | xvhser )}} & {15'b0,cbzbmu27xirmn,afthitl2})
      | ({80{(rzd2hcw89e200ggc )}} & {16'b0,afthitl2})
      | ({80{(dfcpt8muurpn6 )}} & {15'b0,qy4465l158u4avl1st,d19dz7sd0y4n14u7q2iiu,o3odbzchqomo1ykxtvrfo,xb9ns8h_licc_3r22el,zmuacjwbp82p1iy9_f})
      | ({80{(lzu7zvw68i3ihdsw)}} & {16'b1,d19dz7sd0y4n14u7q2iiu,o3odbzchqomo1ykxtvrfo,xb9ns8h_licc_3r22el,zmuacjwbp82p1iy9_f})
    
      | ({80{q1yh6x8lrrng  }} & {7'h00 , cbzbmu27xirmn,bw3242dwyw8g, 7'h00 , dbezizgky8oe_1s,is0m6qik1xe3onr0}) 
      | ({80{tqciamxv2cnjc  }} & {8'h00 ,bw3242dwyw8g,8'h00, is0m6qik1xe3onr0})
      | ({80{h2ip0rex3tgx3  }} & {7'h00 ,qy4465l158u4avl1st,jsfb7rigmw_f0kn1qye3, 7'h40 ,zlhgyh5dfmt_aom,jm_j4gy26gvwm99in}) 
      | ({80{ik95b3bzb6651bvr  }} & {8'h01 ,jsfb7rigmw_f0kn1qye3, 8'h81,jm_j4gy26gvwm99in})
      | ({80{mid3yvd1dc5p_3}} & {7'h00 ,dbezizgky8oe_1s, is0m6qik1xe3onr0, 7'h00,qy4465l158u4avl1st, jsfb7rigmw_f0kn1qye3}) 
      | ({80{d33k1t15iao77sn8eq}} & {8'h00 ,is0m6qik1xe3onr0, 8'h01,jsfb7rigmw_f0kn1qye3}) 
      | ({80{nhk0haqb79ub07mq2b}} & {7'h00 ,zlhgyh5dfmt_aom, jm_j4gy26gvwm99in, 7'h40 , cbzbmu27xirmn,bw3242dwyw8g}) 
      | ({80{ghwvor5rmxzau7tznu}} & {8'h01 ,jm_j4gy26gvwm99in,8'h80, bw3242dwyw8g}) 
      | ({80{ocl0e6_c3wncrmc6 }} & {7'h00 ,cbzbmu27xirmn,bw3242dwyw8g, 7'h00 , zlhgyh5dfmt_aom, jm_j4gy26gvwm99in}) 
      | ({80{qtw5zaawn8u4jd9dy }} & {8'h00 ,bw3242dwyw8g,  8'h01,jm_j4gy26gvwm99in}) 
      | ({80{bsi917d7yfryhti9 }} & {7'h01 ,qy4465l158u4avl1st, jsfb7rigmw_f0kn1qye3,  7'h40 ,  dbezizgky8oe_1s,is0m6qik1xe3onr0}) 
      | ({80{egbv5yccd8p4nkls }} & {8'h01 ,jsfb7rigmw_f0kn1qye3, 8'h80,is0m6qik1xe3onr0}) 
      | ({80{yrqwiv8x45}}  & {8'b0,{32{yxz3vex1f[63]}}, 8'b0,{32{yxz3vex1f[31]}}}) 

         ;


    assign gm0zk3gsgqtkn9_jovpqw3    = g0aqd08ou7rfnv3ndp;
    assign yzauwl2y3mmfl_dtz0c89ze2    = ccbzdmuytukdpcsy26d;
    assign p_q6uot8vlny0p1532oethvbx67 = {80{1'b0}};
    assign e9_hqyec0sd5hbt8qhk_tt_7mhn = {80{1'b0}};

    wire [80-1:0] wrcjvt7pl1j_ = lbo2x74bznoaaigmxjenghis; 
    wire [80-1:0] pql_x0d2rvu = {80{1'b0}}; 
  
  
  
  
  
  wire hqnlo6e255u  = ertz5b_giw | yubia8yl4bb9c;
  wire jo7yipzy2h3jz  = cifajstnxdcka54 | nvxuttrynz12;
  wire t7axzg9ce60zd6 = s_s20wslhcr0ke | yh6x5_h5s1677y;
  wire m8hj_dc0v8ev = ld80dv0dk64f7k_ | ptn87uauvfy;
     
  wire [64-1:0] s8uaye8t3jn74 = {64{g8dm1b58pm6xt}} & yxz3vex1f;
  wire [64-1:0] hi1u2lv6_w = {64{g8dm1b58pm6xt}} & afthitl2;

  
    wire ws8yznrqgmoz33 = ~(|(s8uaye8t3jn74[63:56] ^ hi1u2lv6_w[63:56]));
    wire g3n4v542vigm64 = ~(|(s8uaye8t3jn74[55:48] ^ hi1u2lv6_w[55:48]));
    wire hp35hjpk4rg3f_ = ~(|(s8uaye8t3jn74[47:40] ^ hi1u2lv6_w[47:40]));
    wire rzq4bau1oarknz = ~(|(s8uaye8t3jn74[39:32] ^ hi1u2lv6_w[39:32]));
    wire ad9izx45ntfize = ~(|(s8uaye8t3jn74[31:24] ^ hi1u2lv6_w[31:24]));
    wire knmhuu5ssr3v7r = ~(|(s8uaye8t3jn74[23:16] ^ hi1u2lv6_w[23:16]));
    wire ou443_2_cgxkvg = ~(|(s8uaye8t3jn74[15:8 ] ^ hi1u2lv6_w[15:8 ]));
    wire c_b4_l7s6lqrbt3 = ~(|(s8uaye8t3jn74[7 :0 ] ^ hi1u2lv6_w[7 :0 ]));

  wire [64-1:0] fv68og9aqaq_eys = {
                            {8{ws8yznrqgmoz33}},
                            {8{g3n4v542vigm64}},
                            {8{hp35hjpk4rg3f_}},
                            {8{rzq4bau1oarknz}}, 
                            {8{ad9izx45ntfize}},
                            {8{knmhuu5ssr3v7r}},
                            {8{ou443_2_cgxkvg}},
                            {8{c_b4_l7s6lqrbt3}}};
  
  wire [64-1:0] ktt_uk91lm = {
                            {8{wrcjvt7pl1j_[78]}},
                            {8{wrcjvt7pl1j_[68]}},
                            {8{wrcjvt7pl1j_[58]}},
                            {8{wrcjvt7pl1j_[48]}},  
                            {8{wrcjvt7pl1j_[38]}},
                            {8{wrcjvt7pl1j_[28]}},
                            {8{wrcjvt7pl1j_[18]}},
                            {8{wrcjvt7pl1j_[8 ]}} };

  wire [64-1:0] w18m590v6_dtao = fv68og9aqaq_eys | ktt_uk91lm;

  
  wire xgt92qp6ejym7qe = ~(|(s8uaye8t3jn74[63:48] ^ hi1u2lv6_w[63:48]));
  wire nfirl25xo3pzqe4ql = ~(|(s8uaye8t3jn74[47:32] ^ hi1u2lv6_w[47:32]));
  wire wtlckwx_g1og6da = ~(|(s8uaye8t3jn74[31:16] ^ hi1u2lv6_w[31:16]));
  wire xcj7s5uevcy092w = ~(|(s8uaye8t3jn74[15:0 ] ^ hi1u2lv6_w[15:0 ]));

  wire [64-1:0] wjsbr9e4pkva = {
                             {16{xgt92qp6ejym7qe}},
                             {16{nfirl25xo3pzqe4ql}}, 
                             {16{wtlckwx_g1og6da}},
                             {16{xcj7s5uevcy092w}}};

  
  wire [64-1:0] jwzvxv6uofyke6 = {
                             {16{wrcjvt7pl1j_[76]}},
                             {16{wrcjvt7pl1j_[56]}}, 
                             {16{wrcjvt7pl1j_[36]}},
                             {16{wrcjvt7pl1j_[16]}}};

  wire [64-1:0] i1b7rm2c70dh_ak = wjsbr9e4pkva | jwzvxv6uofyke6;

  wire [64-1:0] ufa33rbvjwk = 
                        ({64{pzqv8u85il7}}  & fv68og9aqaq_eys )  
                       |({64{hqnlo6e255u}}  & ktt_uk91lm ) 
                       |({64{jo7yipzy2h3jz}}  & w18m590v6_dtao )
                       |({64{hmrx98l_nazsdh}} & wjsbr9e4pkva)  
                       |({64{t7axzg9ce60zd6}} & jwzvxv6uofyke6) 
                       |({64{m8hj_dc0v8ev}} & i1b7rm2c70dh_ak)
                       ;

  
  
  
  
  
  
  
  
  
  
  
  
  
  
  

  
  
  
  
  
  
  

  
  
  
  
  
  
  

  
  
  
  
  

  
  
  
  
  

 
  
  
  
  
  
  


  
  
  wire [64-1:0] pnoaou8emb9_b = {
                          (wrcjvt7pl1j_[78] ? afthitl2[63:56] : yxz3vex1f[63:56]),
                          (wrcjvt7pl1j_[68] ? afthitl2[55:48] : yxz3vex1f[55:48]),
                          (wrcjvt7pl1j_[58] ? afthitl2[47:40] : yxz3vex1f[47:40]),
                          (wrcjvt7pl1j_[48] ? afthitl2[39:32] : yxz3vex1f[39:32]), 
                          (wrcjvt7pl1j_[38] ? afthitl2[31:24] : yxz3vex1f[31:24]),
                          (wrcjvt7pl1j_[28] ? afthitl2[23:16] : yxz3vex1f[23:16]),
                          (wrcjvt7pl1j_[18] ? afthitl2[15:8 ] : yxz3vex1f[15:8 ]),
                          (wrcjvt7pl1j_[8 ] ? afthitl2[7 :0 ] : yxz3vex1f[7 :0 ])};

  wire [64-1:0] s9_1a5sf0e = {
                          (wrcjvt7pl1j_[78] ? yxz3vex1f[63:56] : afthitl2[63:56]),
                          (wrcjvt7pl1j_[68] ? yxz3vex1f[55:48] : afthitl2[55:48]),
                          (wrcjvt7pl1j_[58] ? yxz3vex1f[47:40] : afthitl2[47:40]),
                          (wrcjvt7pl1j_[48] ? yxz3vex1f[39:32] : afthitl2[39:32]), 
                          (wrcjvt7pl1j_[38] ? yxz3vex1f[31:24] : afthitl2[31:24]),
                          (wrcjvt7pl1j_[28] ? yxz3vex1f[23:16] : afthitl2[23:16]),
                          (wrcjvt7pl1j_[18] ? yxz3vex1f[15:8 ] : afthitl2[15:8 ]),
                          (wrcjvt7pl1j_[8 ] ? yxz3vex1f[7 :0 ] : afthitl2[7 :0 ])};

  wire [64-1:0] wokr41xa4vigqpe  =  ({64{c79vtanyxxram | rpacmi1zwp95 }} & pnoaou8emb9_b)
                                     |  ({64{kv8kqf2jbw7 | gwqnhrtp4 }} & s9_1a5sf0e);  
  
  wire [64-1:0] s0jem23hm369m_ = {
                           (wrcjvt7pl1j_[76] ? afthitl2[63:48] : yxz3vex1f[63:48]),
                           (wrcjvt7pl1j_[56] ? afthitl2[47:32] : yxz3vex1f[47:32]),
                           (wrcjvt7pl1j_[36] ? afthitl2[31:16] : yxz3vex1f[31:16]),
                           (wrcjvt7pl1j_[16] ? afthitl2[15:0 ] : yxz3vex1f[15:0 ])};

  wire [64-1:0] b4ghg6beg = {
                           (wrcjvt7pl1j_[76] ? yxz3vex1f[63:48] : afthitl2[63:48]),
                           (wrcjvt7pl1j_[56] ? yxz3vex1f[47:32] : afthitl2[47:32]),
                           (wrcjvt7pl1j_[36] ? yxz3vex1f[31:16] : afthitl2[31:16]),
                           (wrcjvt7pl1j_[16] ? yxz3vex1f[15:0 ] : afthitl2[15:0 ])};

  wire [64-1:0] ire1qcgu3cincas  =  ({64{uo2vcr1g3uksaw | l30nioha_vjc }} & s0jem23hm369m_)
                                        |({64{zd6qkrf4rnr | lcecqtg_qt8r }} & b4ghg6beg);  
  
  wire [64-1:0] t4lezi94p =  wrcjvt7pl1j_[32] ? {{64-32{afthitl2[31]}},afthitl2[31:0]} : {{64-32{yxz3vex1f[31]}},yxz3vex1f[31:0]};
  wire [64-1:0] fcnp1chzz646r =  wrcjvt7pl1j_[32] ? {{64-32{yxz3vex1f[31]}},yxz3vex1f[31:0]} : {{64-32{afthitl2[31]}},afthitl2[31:0]}; 

  wire [64-1:0] atxzdtmrjbea  =  ({64{iemiml6mv3q}} & t4lezi94p)
                                       |({64{y5gwqbpjit}} & fcnp1chzz646r);  

  wire [64-1:0] j0z_c8aj817e5q =  {
                                      (wrcjvt7pl1j_[72] ? bw3242dwyw8g : b_xqc3mgz11e),
                                      (wrcjvt7pl1j_[32] ? is0m6qik1xe3onr0 : x4vwdbhy47grdx6)
                                     };


  wire [64-1:0] p57xuv__ifghc =  {
                                      (wrcjvt7pl1j_[72] ? b_xqc3mgz11e : bw3242dwyw8g),
                                      (wrcjvt7pl1j_[32] ? x4vwdbhy47grdx6 : is0m6qik1xe3onr0)
                                     };

  wire [64-1:0] siaf_d_tl16ww6r9  =  ({64{y5rwe1utr6 | gzsw9ptxn8f}} & j0z_c8aj817e5q)
                                        |({64{ycwtj7_ux8co | lhtfca0wde}} & p57xuv__ifghc);  




  wire [64-1:0] ivcpoenlvs_zrk8 = ({64{c9hqqulyow5pvq }} & wokr41xa4vigqpe )  
                                   | ({64{g2s8ge1hum_lb}} & ire1qcgu3cincas)  
                                   | ({64{brrzcx4c49ey }} & atxzdtmrjbea )
                                   | ({64{pmct0ov7_sv0}} & siaf_d_tl16ww6r9)
                                   ;



  
  
  wire evmvst7bfbhg = kdnn4d_qr2_jt4n3 | au1gh_eazilnry  | svzbv80johvs  
                    | ijnb_gpo7xg3r1 | ltcar0xe__n9nh61k | yed1aglcls65oj
                    | hlx2yqcuw7mugxd  | gjgqa949f4epnz | n0uej4ag_la  
                    | azm_djrz3r5raujmu  | sred4q00s3ugie6bhl 
                    | jcv5t8qp92n4yn_ | h_u6dnfrybg78e0tn  | i7uc6ffwjktqvuq4q6;
  

  wire dhtimibzgwimr2  = kdnn4d_qr2_jt4n3  | svzbv80johvs | ypjg3i7dl0;
  wire k1qk74_avk = ijnb_gpo7xg3r1 | yed1aglcls65oj| rpk5hmf4ck8wgf;
  wire f0axh_3szq  = n0uej4ag_la  | jcv5t8qp92n4yn_ | hlx2yqcuw7mugxd  | gjgqa949f4epnz| fydew0oon ;
  wire zhj0mle6aadmqa = azm_djrz3r5raujmu | sred4q00s3ugie6bhl | yrqwiv8x45;
  wire nvuerngsqym = h_u6dnfrybg78e0tn | i7uc6ffwjktqvuq4q6;                
  wire wfyu80hvukirek = f0ohe956w | au1gh_eazilnry;
  wire jdi1rvyhuok3zzz = ex4t35fb30 | ltcar0xe__n9nh61k;
  wire zprrej81j8e7 = evmvst7bfbhg | gv93tjc7rha;
  
  wire[2:0] qjlacm_go = ({3{dhtimibzgwimr2 }} & 3'b000) 
                      | ({3{k1qk74_avk}} & 3'b001) 
                      | ({3{f0axh_3szq }} & 3'b010)
                      | ({3{zhj0mle6aadmqa}} & 3'b110)
                      | ({3{nvuerngsqym}} & 3'b011)
                      | ({3{wfyu80hvukirek}} & 3'b100)
                      | ({3{jdi1rvyhuok3zzz}} & 3'b101)
                         ;

  wire nvrjuq  = kdnn4d_qr2_jt4n3 | au1gh_eazilnry;
  wire s5hzzmy_  = svzbv80johvs;
  wire c1bldoa = ijnb_gpo7xg3r1 | ltcar0xe__n9nh61k | hlx2yqcuw7mugxd;
  wire wimx049 = qe0l_afxffya5u7 | avyzty88svfq | t_ph70ukeyywgs | qdsnvv2pfb;
  wire wz05g5r = n0uej4ag_la | azm_djrz3r5raujmu;
  wire kawmn4y5ol33 = jcv5t8qp92n4yn_ | t8eyqdo1vo1 | vky13xw8f8jbgve;
  wire wxg4q_ly = gv93tjc7rha;
  wire hx3hr203 = hev7phfsjoj2rx | hbtor719sgm6b1 | oaxsuvqvhxpls6h | ryxvixwjxi_ub7ot; 
  wire k99rxinyba = xjhmnd_xa2du_6g | m8a77l1aday | vg2q1cvp3u8g | m30h0_l1chll9; 
  wire qghwr_71jegd = h_u6dnfrybg78e0tn;
  wire ooams9rewa96 = i7uc6ffwjktqvuq4q6;
  wire[3:0] ck6o6flrt  = ({4{nvrjuq  }} & 4'b0000)  
                      | ({4{s5hzzmy_  }} & 4'b0001)  
                      | ({4{c1bldoa }} & 4'b0010)  
                      | ({4{wimx049 }} & 4'b0011) 
                      | ({4{wz05g5r }} & 4'b0100)  
                      | ({4{kawmn4y5ol33 }} & 4'b0101)  
                      | ({4{wxg4q_ly }} & 4'b0110) 
                      | ({4{hx3hr203}} & 4'b0111) 
                      | ({4{k99rxinyba}} & 4'b1000)  
                      | ({4{qghwr_71jegd }} & 4'b1001)  
                      | ({4{ooams9rewa96 }} & 4'b1010)  
                        ;
  
  wire k65w3sg3e = (kdnn4d_qr2_jt4n3 | au1gh_eazilnry | a35tr1zbyo  
                | ijnb_gpo7xg3r1 | ltcar0xe__n9nh61k  | avyzty88svfq 
                | pfvv152dbk8llva | hev7phfsjoj2rx |  go1xs0z8qd8zwe1 | xjhmnd_xa2du_6g   
                | a0mwf5tzfds7 | hbtor719sgm6b1 |  dmvcpit4cpt | m8a77l1aday   
                | zg4vqn28eg | oaxsuvqvhxpls6h |  a42iwg_hdrm3vy | vg2q1cvp3u8g   
                | qp2h493he29 | ryxvixwjxi_ub7ot |  tgrv6fv3nm45 | m30h0_l1chll9   
                | hlx2yqcuw7mugxd |  qdsnvv2pfb   
                | n0uej4ag_la |  cyen5b13oh4_xj   
                | azm_djrz3r5raujmu |  vky13xw8f8jbgve   
                | h_u6dnfrybg78e0tn |  cj6waeyow1   
               );
  wire r2zqwi571k5ppf;
    wire [64-1:0] wj1ukvyuohpl4xrz  ;
    wire [64-1:0] pb7kaoib_jjclvbf_r;
  s20vasmduccat9_3 pfjomapoyb6fgakd41 (
      
      .pugy9o4i2pr3ns8yo3       (wrcjvt7pl1j_),
      .qg0gj_1bem7nt1wek5w2bc     (pql_x0d2rvu),
      .wip5afkxmbs5dou       (qjlacm_go     ), 
      .dgvew5k86brk_8uip        (ck6o6flrt      ), 
      .phlh_dccd75w7xikxtg03      (k65w3sg3e        ), 
      .jqnqhlv1gjf2k3xg4      (zprrej81j8e7      ), 
      .vvoozaywykiwmels       (wj1ukvyuohpl4xrz   ),
      .m50l82p03g15y_ehxthx1     (pb7kaoib_jjclvbf_r ),
      .hsvg_y2njolj1bl          (r2zqwi571k5ppf    )
  );

  

  wire b9r3isyjg1w3h_gqmdzb9xou = f0ohe956w | ex4t35fb30 | wsflp3hzxrkbzt | hj4cvyrejb | rmydqk33eq | dow464urmsra;
  wire [64-1:0] pr7v58nej9domw9c7 =  
        ({64{e03ora27k00u_e   }} & {wrcjvt7pl1j_[77:70],wrcjvt7pl1j_[67:60],wrcjvt7pl1j_[57:50],wrcjvt7pl1j_[47:40], 
                                        wrcjvt7pl1j_[37:30],wrcjvt7pl1j_[27:20],wrcjvt7pl1j_[17:10],wrcjvt7pl1j_[ 7: 0]})
      | ({64{umletcb8zgwqs | iqxdtyt_g9dloiv }} 
                                     & {wrcjvt7pl1j_[78:71],wrcjvt7pl1j_[68:61],wrcjvt7pl1j_[58:51],wrcjvt7pl1j_[48:41], 
                                        wrcjvt7pl1j_[38:31],wrcjvt7pl1j_[28:21],wrcjvt7pl1j_[18:11],wrcjvt7pl1j_[ 8: 1]})
      | ({64{cr75ulfp       }} & ufa33rbvjwk )
      | ({64{jpt8d5z4s    }} & ivcpoenlvs_zrk8)
      | ({64{k5tw9oeheqlih4  }} & {wrcjvt7pl1j_[75:60],wrcjvt7pl1j_[55:40],wrcjvt7pl1j_[35:20],wrcjvt7pl1j_[15:0]})
      | ({64{imjs03vic384a18 | fsok4w6z0ij77ih}} 
                                     & {wrcjvt7pl1j_[76:61],wrcjvt7pl1j_[56:41],wrcjvt7pl1j_[36:21],wrcjvt7pl1j_[16:1]})
      | ({64{u340gmafpm_q0kft | gami8f4x_a1qsq }} 
                                     & {{64-32{wrcjvt7pl1j_[32]}},wrcjvt7pl1j_[32: 1]})
      | ({64{ivgy7v_9d }} 
                                     & {{64-32{1'b0}},wrcjvt7pl1j_[32: 1]})
      | ({64{xvhser}} 
                                     & {wrcjvt7pl1j_[64:1]})
      | ({64{lwh7ejgwbe0y3xd6  }} & wrcjvt7pl1j_[63: 0])
      | ({64{e6mszw3shdp5 | p1b08_so0a9eejxiuw}} & wrcjvt7pl1j_[64: 1])
      | ({64{dhtimibzgwimr2 | k1qk74_avk | f0axh_3szq | zhj0mle6aadmqa}} 
                                     & {wj1ukvyuohpl4xrz[63:56],wj1ukvyuohpl4xrz[55:48],wj1ukvyuohpl4xrz[47:40],wj1ukvyuohpl4xrz[39:32],
                                        wj1ukvyuohpl4xrz[31:24],wj1ukvyuohpl4xrz[23:16],wj1ukvyuohpl4xrz[15: 8],wj1ukvyuohpl4xrz[ 7: 0]})
      | ({64{h_u6dnfrybg78e0tn | i7uc6ffwjktqvuq4q6 | b9r3isyjg1w3h_gqmdzb9xou}} 
                                     & {wj1ukvyuohpl4xrz[64-1:0]})
      | ({64{ijlmx1ho6tz  }} & {wrcjvt7pl1j_[71:40],wrcjvt7pl1j_[31:0]})
      | ({64{x3e45geoeepfd_9pa | pvy_15wdbehc4s63n}} 
                                     & {wrcjvt7pl1j_[72:41],wrcjvt7pl1j_[32:1]})
        ;

  assign ymi25pa6qmirfeb9 = m0mq6jm4ys | mf5fcnu2azr | h0xl_5;
  assign iz4sa6lcipb1cjsz_ = m0mq6jm4ys | xvhser | h0xl_5;
  
  
  wire [7:0] txv1tfb04aa = ({8{wrcjvt7pl1j_[78]}} & (~wrcjvt7pl1j_[77:70])) | ({8{~wrcjvt7pl1j_[78]}} & wrcjvt7pl1j_[77:70]) ; 
  wire [7:0] pzzm7pbhp = ({8{wrcjvt7pl1j_[68]}} & (~wrcjvt7pl1j_[67:60])) | ({8{~wrcjvt7pl1j_[68]}} & wrcjvt7pl1j_[67:60]) ; 
  wire [7:0] gc7w3onzb = ({8{wrcjvt7pl1j_[58]}} & (~wrcjvt7pl1j_[57:50])) | ({8{~wrcjvt7pl1j_[58]}} & wrcjvt7pl1j_[57:50]) ; 
  wire [7:0] blea2gjhi = ({8{wrcjvt7pl1j_[48]}} & (~wrcjvt7pl1j_[47:40])) | ({8{~wrcjvt7pl1j_[48]}} & wrcjvt7pl1j_[47:40]) ; 
  wire [7:0] tk_l5nlhk10 = ({8{wrcjvt7pl1j_[38]}} & (~wrcjvt7pl1j_[37:30])) | ({8{~wrcjvt7pl1j_[38]}} & wrcjvt7pl1j_[37:30]) ; 
  wire [7:0] rmjiwsgg = ({8{wrcjvt7pl1j_[28]}} & (~wrcjvt7pl1j_[27:20])) | ({8{~wrcjvt7pl1j_[28]}} & wrcjvt7pl1j_[27:20]) ; 
  wire [7:0] sze9miov8 = ({8{wrcjvt7pl1j_[18]}} & (~wrcjvt7pl1j_[17:10])) | ({8{~wrcjvt7pl1j_[18]}} & wrcjvt7pl1j_[17:10]) ; 
  wire [7:0] qo3ep5rrww = ({8{wrcjvt7pl1j_[ 8]}} & (~wrcjvt7pl1j_[ 7: 0])) | ({8{~wrcjvt7pl1j_[ 8]}} & wrcjvt7pl1j_[ 7: 0]) ; 

  wire [7:0] ezeo6u2btla = {wrcjvt7pl1j_[78], wrcjvt7pl1j_[68], wrcjvt7pl1j_[58], wrcjvt7pl1j_[48],
                        wrcjvt7pl1j_[38], wrcjvt7pl1j_[28], wrcjvt7pl1j_[18], wrcjvt7pl1j_[ 8]};
  wire [1:0] wfdeqdy8dj029;
  wire [1:0] ml4qiwrdp1y953a9u;
  wire [1:0] qylju6u_ms6p;
  wire [1:0] vnahsd7ljbw5ck7z;
  wire [2:0] gd7hglmtecg;
  wire [2:0] tzwvwhlnlce;
  gg0ubjxsd5riswv #(2) zcic5uwj6hobiorywg8cw(.frgfco({1'b0,ezeo6u2btla[7]}), 
                                           .ii({1'b0,ezeo6u2btla[6]}), 
                                           .fij51v({1'b0,ezeo6u2btla[5]}), 
                                           .cuzhl9({1'b0,ezeo6u2btla[4]}), 
                                           .c (wfdeqdy8dj029), 
                                           .s (ml4qiwrdp1y953a9u));
  gg0ubjxsd5riswv #(2) fdmgfjooq1d5jx3s44qbrnk(.frgfco({1'b0,ezeo6u2btla[3]}), 
                                           .ii({1'b0,ezeo6u2btla[2]}), 
                                           .fij51v({1'b0,ezeo6u2btla[1]}), 
                                           .cuzhl9({1'b0,ezeo6u2btla[0]}), 
                                           .c (qylju6u_ms6p), 
                                           .s (vnahsd7ljbw5ck7z));
  gg0ubjxsd5riswv #(3) xlkjaigo8wrdj1gug8ir1rbu(.frgfco({1'b0,wfdeqdy8dj029}), 
                                           .ii({1'b0,ml4qiwrdp1y953a9u}), 
                                           .fij51v({1'b0,qylju6u_ms6p}), 
                                           .cuzhl9({1'b0,vnahsd7ljbw5ck7z}), 
                                           .c (gd7hglmtecg), 
                                           .s (tzwvwhlnlce));
  wire [3:0] roapbsh_saei = {1'b0,gd7hglmtecg} + {1'b0,tzwvwhlnlce};
  
  assign s6tonq08_ria84ebdjlir = ({64+4{h0xl_5}} & {roapbsh_saei,txv1tfb04aa,pzzm7pbhp,gc7w3onzb,blea2gjhi,
                                                               tk_l5nlhk10,rmjiwsgg,sze9miov8,qo3ep5rrww});

  wire [64-1:0]  ucdthfkff54i3uyept0tyx = pr7v58nej9domw9c7; 

  assign ya1whb4lzd9i6g2qr2yu5enshd   = ucdthfkff54i3uyept0tyx;
  assign fl1olcli4mhazuy960y16sqh63s5 = {64{1'b0}};
  assign cxxjqchsz57vq2dff3d0j = r2zqwi571k5ppf;



endmodule




















module cwe8y4czjwvbx6znvqv5wg09qsfw(
    input [64:0] ho7hbln__5mzkxd,
    input [64:0] e7e6yf3rwo5s,
    input [64:0] zpa9wht92mu,
    input [64:0] mx84o3rvy8,
    input [64:0] l6dri5njf3xti3j,
    input [64:0] d986vh8a8wdpib0,
    input [64:0] xfnf1gelth,
    input [64:0] n2t6qssk9yjxv,
    input [64:0] nvjphm8kit9,
    input [33:0] yj4jcdxd_qu6m3mon,
    input [34:0] af86r5akqaznjghqqft,
    output [66:0] wrcjvt7pl1j_
);



wire [66:0] lfjxb788ju8p5z56tj;
wire [66:0] pmjc2r4mlimgsd1u7;
wire [66:0] fb5kiq1vtucdrem_;
wire [66:0] g69w6k4vbwhlsgn5p6wi;
wire [66:0] mwonk7q78krtp35lt;
wire [66:0] p2d4ghaaopmvw;
wire [66:0] zp2qz4re4cl228e38rt;
wire [66:0] tp76l_5mv705xq8cgq;
wire [66:0] hufizt69101tjw4;
wire [66:0] p132_ik3uo6mxhks82;
wire [66:0] a0_j63tohthvfeu;
wire [66:0] zaghc2q5gzfv80d9kt;

wire [64:0] v4wb28582p1y13tpsm;
wire [64:0] lr88j9kepgbptohd;
wire [64:0] y1t85ych1ui_co0h_;
wire [64:0] v_2j97vhdvhg1qwa3;
wire [64:0] xe1ree9fnb0apt1kz;

assign  lfjxb788ju8p5z56tj = {{2{e7e6yf3rwo5s[64]}}, e7e6yf3rwo5s};
assign  pmjc2r4mlimgsd1u7 = {{2{zpa9wht92mu[64]}}, zpa9wht92mu};
assign  fb5kiq1vtucdrem_ = {{2{mx84o3rvy8[64]}}, mx84o3rvy8};
assign  g69w6k4vbwhlsgn5p6wi = {{2{l6dri5njf3xti3j[64]}}, l6dri5njf3xti3j};
assign  zp2qz4re4cl228e38rt = {{2{d986vh8a8wdpib0[64]}}, d986vh8a8wdpib0};
assign  tp76l_5mv705xq8cgq = {{2{xfnf1gelth[64]}}, xfnf1gelth};
assign  hufizt69101tjw4 = {{2{n2t6qssk9yjxv[64]}}, n2t6qssk9yjxv};
assign  p132_ik3uo6mxhks82 = {{2{nvjphm8kit9[64]}}, nvjphm8kit9};


assign  v4wb28582p1y13tpsm = ho7hbln__5mzkxd;
assign  lr88j9kepgbptohd = {{31{yj4jcdxd_qu6m3mon[33]}}, yj4jcdxd_qu6m3mon};
assign  y1t85ych1ui_co0h_ = {30'b0, af86r5akqaznjghqqft};

  gg0ubjxsd5riswv #(67) odlt_zna1fp0es2d(.frgfco(lfjxb788ju8p5z56tj), 
                                      .ii(pmjc2r4mlimgsd1u7), 
                                      .fij51v(fb5kiq1vtucdrem_), 
                                      .cuzhl9(g69w6k4vbwhlsgn5p6wi), 
                                      .c (mwonk7q78krtp35lt), 
                                      .s (p2d4ghaaopmvw));

  gg0ubjxsd5riswv #(67) xt4crwlv7g41l316t(.frgfco(zp2qz4re4cl228e38rt), 
                                      .ii(tp76l_5mv705xq8cgq), 
                                      .fij51v(hufizt69101tjw4), 
                                      .cuzhl9(p132_ik3uo6mxhks82), 
                                      .c (a0_j63tohthvfeu), 
                                      .s (zaghc2q5gzfv80d9kt));

  opvhnxssc7yjqmd3 #(65) e8_db00cty22_0a(.frgfco(v4wb28582p1y13tpsm), 
                                      .ii(lr88j9kepgbptohd), 
                                      .fij51v(y1t85ych1ui_co0h_), 
                                      .c (v_2j97vhdvhg1qwa3), 
                                      .s (xe1ree9fnb0apt1kz)); 


wire [68:0] ta1eiqchseappkrl;
wire [68:0] qyzgt2vysfapnj3szu;
wire [68:0] mzw2d5094vo17qupz;
wire [68:0] dj93swsd9warg;
wire [68:0] wmg0jo8v5easew;

wire [68:0] hqmry1jntyqzi4ab;
wire [68:0] i3z60qjrf5y1q693g;
wire [68:0] or5i_zgol1sux33;
wire [68:0] heyrakjwqzl27q;
wire [68:0] homl8mgryidbw_z;

assign ta1eiqchseappkrl = {{2{mwonk7q78krtp35lt[66]}},mwonk7q78krtp35lt};
assign qyzgt2vysfapnj3szu = {{2{p2d4ghaaopmvw[66]}},p2d4ghaaopmvw};
assign mzw2d5094vo17qupz = {{2{a0_j63tohthvfeu[66]}},a0_j63tohthvfeu};
assign hqmry1jntyqzi4ab = {{2{zaghc2q5gzfv80d9kt[66]}},zaghc2q5gzfv80d9kt};
assign i3z60qjrf5y1q693g = {{4{v_2j97vhdvhg1qwa3[64]}},v_2j97vhdvhg1qwa3};
assign or5i_zgol1sux33 = {{4{xe1ree9fnb0apt1kz[64]}},xe1ree9fnb0apt1kz};

  opvhnxssc7yjqmd3 #(69) uw808c6pfbjdwc(.frgfco(ta1eiqchseappkrl), 
                                      .ii(qyzgt2vysfapnj3szu), 
                                      .fij51v(mzw2d5094vo17qupz), 
                                      .c (dj93swsd9warg), 
                                      .s (wmg0jo8v5easew)); 

  opvhnxssc7yjqmd3 #(69) v4582i3ayu76xh6q(.frgfco(hqmry1jntyqzi4ab), 
                                      .ii(i3z60qjrf5y1q693g), 
                                      .fij51v(or5i_zgol1sux33), 
                                      .c (heyrakjwqzl27q), 
                                      .s (homl8mgryidbw_z)); 



wire [70:0] ig5nwoqiqun75gvb6hd;
wire [70:0] bzehn50i29cp_c3;
wire [70:0] gqy9qfc88c5nlx_sh9u8;
wire [70:0] c2qu200yhu_qkb0duc3;
wire [70:0] wgx5nl1gdrk6bnd;
wire [70:0] vyd77edvnmpus;

assign ig5nwoqiqun75gvb6hd = {{2{dj93swsd9warg[68]}}, dj93swsd9warg};
assign bzehn50i29cp_c3 = {{2{wmg0jo8v5easew[68]}}, wmg0jo8v5easew};
assign gqy9qfc88c5nlx_sh9u8 = {{2{heyrakjwqzl27q[68]}}, heyrakjwqzl27q};
assign c2qu200yhu_qkb0duc3 = {{2{homl8mgryidbw_z[68]}}, homl8mgryidbw_z};

  gg0ubjxsd5riswv #(71) z169bbuutkmguqkkoi(.frgfco(ig5nwoqiqun75gvb6hd), 
                                      .ii(bzehn50i29cp_c3), 
                                      .fij51v(gqy9qfc88c5nlx_sh9u8), 
                                      .cuzhl9(c2qu200yhu_qkb0duc3), 
                                      .c (wgx5nl1gdrk6bnd), 
                                      .s (vyd77edvnmpus));

wire [71:0] v6yt5ccneunjpdhyg2 = {wgx5nl1gdrk6bnd[70],wgx5nl1gdrk6bnd} + {vyd77edvnmpus[70],vyd77edvnmpus}; 

assign wrcjvt7pl1j_ = v6yt5ccneunjpdhyg2[66:0];

endmodule



















module a37xq53sqhw4q7cxzwmz(
  input tvdvyldvwqhx7g8r9di,
  output izj2me9tmzxitrpzl1tr,
  output rgcs7q5ke7h8fte8jecm,
  input  pzhh8hyzbdb80ac8sdd_49,
  input  t_998ilixet4pdvdkju,
  input [64-1:0] l7mctsr6ttfp83pl8jo7,
  input  a2o96wlgs_5sqzm2a7ba_,
  output cwmxezrc3jv6hzxcfc,
  input  uig3ujuyq0_61kqb,
  input j_rvclhfbeig5cqeb3_,
  input gdebc5b6o6bv57ax1bw,
  input w363n7ci30h3kw2g1oktlj1puysbju,
  input lygqe2977b3fd_0eit3wg_nnfirn,
  input th583ebkp2cj56crsivefzygk81o65_h2,
  input vz2rm7lc9ctulrdhe1kv8wdmobft,
  input hlmhgsbtxsmi7y1a7oshnntydp27pj,
  input dshcfm3k8zhyftxq_xw9j106j59z7notf,
  input [63:0] usrh37qm6nz8yamj6_h_pmbv5,
  input [63:0] mipc_c8bfwk8khoqgtsj65f1f,
  input [63:0] pm3m6aucefl9oas0vqgwfm,
  input [63:0] yc5f_bw94gu1iari4qpmo269z,
  input [5-1:0]  bj9det3k1xe2rn,
  input [5-1:0] cvhwe_6rucj7,
  input [64-1:0] amgi_rqhtd007,
  input [64-1:0] xo5bwsw4j8a,
  input [64+3:0] xcp0v_slt0baqx9h6px,
  input [105-1:0] a4p3huz_qaf92as,
  input [105-1:0] e4_5otstd9ttd5eebgmf,
  input [50-1:0] n6izg3jvgts,
  input  [4-1:0] jsz4fvx2s3ijb5,
  output [64-1:0] nb3w1rq_ny95rvrt,        
  output vjkz8n6i44pc7o,
  output xc2becmsn4fcniw6ks,        
  output [4-1:0] p_yx415so7q1vohijb,
  input gf33atgy,
  input ru_wi
);

  wire eojd5fb       = a4p3huz_qaf92as[15]; 
  wire o0snf_gso30ua      = 1'b0;
  wire xn1f1pv3xq9j     = 1'b0;
  wire ch1i9dybknbuw      = a4p3huz_qaf92as[16]; 
  wire ntp3h6qp      = a4p3huz_qaf92as[9];
  wire gqej_k2u1l4m      = a4p3huz_qaf92as[17];
  wire s7h0yqvmtsxj      = a4p3huz_qaf92as[18];
  wire wgvga5xo      = a4p3huz_qaf92as[19];
  wire fx9_o1uw35rbg      = a4p3huz_qaf92as[20];
  wire kn5fa7ovnhnx      = a4p3huz_qaf92as[21];
  wire u_k_oszo40vsx      = a4p3huz_qaf92as[22];
  wire ksqlq_qg3d     = a4p3huz_qaf92as[10];
  wire yyrimhfarrpqm     = a4p3huz_qaf92as[5];
  wire mcnxhlts_l6su5y    = a4p3huz_qaf92as[6];
  wire mfqddwpbt3pb     = a4p3huz_qaf92as[7];
  wire k0zpfgcn5bak    = a4p3huz_qaf92as[8];
  wire r_si8qamg50      = a4p3huz_qaf92as[11];
  wire vc8jimsljb     = a4p3huz_qaf92as[12];
  wire cqcm3m7k      = a4p3huz_qaf92as[13];
  wire l1fra0t6408e_6     = a4p3huz_qaf92as[14];
  wire zt47pxlvcnvwaj     = e4_5otstd9ttd5eebgmf[48];
  wire mxh5z6vyj5     = e4_5otstd9ttd5eebgmf[49];
  wire dcd8vqqpxs     = e4_5otstd9ttd5eebgmf[50];
  wire w4hjaq5ha     = e4_5otstd9ttd5eebgmf[103];
  wire gddu1322qyclw5    = e4_5otstd9ttd5eebgmf[104];
  wire uqitfc00xwe     = e4_5otstd9ttd5eebgmf[98];
  wire mtm0jygbpquyx_     = e4_5otstd9ttd5eebgmf[101];
  wire oi_q1zg22f_j     = e4_5otstd9ttd5eebgmf[102];
  wire r1h7wsdxc      = e4_5otstd9ttd5eebgmf[99];
  wire akokb5adw5      = e4_5otstd9ttd5eebgmf[100];
  wire i3t5mrrybl5      = e4_5otstd9ttd5eebgmf[97];
  wire dr32dt_a9g     = e4_5otstd9ttd5eebgmf[7];
  wire jctnij88_5a      = e4_5otstd9ttd5eebgmf[8];
  wire mydhpyzp8hjwy     = e4_5otstd9ttd5eebgmf[9];
  wire rtuq1m6b67r7u    = e4_5otstd9ttd5eebgmf[10];
  wire r_39wh4gt2t15     = e4_5otstd9ttd5eebgmf[11];
  wire nhvy44ogg7437     = e4_5otstd9ttd5eebgmf[12];
  wire lm0p0_l8v3c     = e4_5otstd9ttd5eebgmf[13];
  wire m2p4w1oz_anbe    = e4_5otstd9ttd5eebgmf[14];
  wire dc4k61sy3n_z1m     = e4_5otstd9ttd5eebgmf[15];
  wire ychqrju9d5fye7j    = e4_5otstd9ttd5eebgmf[16];
  wire d1zrh920nh    = e4_5otstd9ttd5eebgmf[17];
  wire uu7kphuq      = e4_5otstd9ttd5eebgmf[6];
  wire cnluzxjjp1rcx     = e4_5otstd9ttd5eebgmf[5];
  wire ig7u5q3yu6kicnh    = e4_5otstd9ttd5eebgmf[18];
  wire exe5zfxbfu0_8    = e4_5otstd9ttd5eebgmf[19];
  wire y7jlwr4xt5op   = e4_5otstd9ttd5eebgmf[20];
  wire tu3h2v18zj    = e4_5otstd9ttd5eebgmf[21];
  wire hc_xm8msfc3   = e4_5otstd9ttd5eebgmf[22];
  wire edwtafv6h     = e4_5otstd9ttd5eebgmf[23];
  wire fqhz535idl    = e4_5otstd9ttd5eebgmf[24];
  wire yptobqxpymp       = e4_5otstd9ttd5eebgmf[25];
  wire n64e5158axn6      = e4_5otstd9ttd5eebgmf[26];
  wire wq_as4te8v_b       = e4_5otstd9ttd5eebgmf[27];
  wire ga7v537skbsy      = e4_5otstd9ttd5eebgmf[28];
  wire sjjokf_h      = e4_5otstd9ttd5eebgmf[29];
  wire n4q1xxu4x_3hl      = e4_5otstd9ttd5eebgmf[30];
  wire hq5o156te      = e4_5otstd9ttd5eebgmf[31];
  wire tdmjh8lo4z5      = e4_5otstd9ttd5eebgmf[32];
  wire iatq6q6eq      = e4_5otstd9ttd5eebgmf[33];
  wire hqgpv7iwel4t     = e4_5otstd9ttd5eebgmf[34];
  wire rte1rpxc      = e4_5otstd9ttd5eebgmf[35];
  wire scwyr94dp     = e4_5otstd9ttd5eebgmf[36];
  wire xu4g6q5o_     = e4_5otstd9ttd5eebgmf[37];
  wire jqjgwcghbu      = e4_5otstd9ttd5eebgmf[38];
  wire xpm18ev4bbldh     = e4_5otstd9ttd5eebgmf[39];
  wire lm6sobl4jhpz      = e4_5otstd9ttd5eebgmf[40];
  wire sdiqw5ujf      = e4_5otstd9ttd5eebgmf[41];
  wire w3m1avjrhe    = e4_5otstd9ttd5eebgmf[42];
  wire b3sltjkxd     = e4_5otstd9ttd5eebgmf[43];
  wire nbcmgtqjii6     = e4_5otstd9ttd5eebgmf[44];
  wire he1npja1q     = e4_5otstd9ttd5eebgmf[45];
  wire e8kmdrlj7pv    = e4_5otstd9ttd5eebgmf[46];
  wire y44x7fnhxvoz85    = e4_5otstd9ttd5eebgmf[47];
  wire hbgz8fj2       = e4_5otstd9ttd5eebgmf[51];
  wire h80eeiznk     = e4_5otstd9ttd5eebgmf[52];
  wire e14xup9fo8q72     = e4_5otstd9ttd5eebgmf[53];
  wire qz487t2wc1     = e4_5otstd9ttd5eebgmf[54];
  wire m4ru19tg0     = e4_5otstd9ttd5eebgmf[55];
  wire b9j3bhreofzf    = e4_5otstd9ttd5eebgmf[56];
  wire uz5zh9l2ar1q    = e4_5otstd9ttd5eebgmf[57];
  wire l_rmt2esx6tvr     = e4_5otstd9ttd5eebgmf[58];
  wire mku_74ifgnfieu2    = e4_5otstd9ttd5eebgmf[59];
  wire a1q5p89kjv     = e4_5otstd9ttd5eebgmf[60];
  wire hniqik4tqx     = e4_5otstd9ttd5eebgmf[61];
  wire znkntww0_qvy0     = e4_5otstd9ttd5eebgmf[62];
  wire fj3p9vcal5     = e4_5otstd9ttd5eebgmf[63];
  wire yuimu6qrm3    = e4_5otstd9ttd5eebgmf[64];
  wire i7uhvhnm5dzd0    = e4_5otstd9ttd5eebgmf[65];
  wire o2476dr5c9g     = e4_5otstd9ttd5eebgmf[66];
  wire vmjyb2bbjdd1t4     = e4_5otstd9ttd5eebgmf[67];
  wire h_aqv6_zs     = e4_5otstd9ttd5eebgmf[96];
  wire ylft74onr      = e4_5otstd9ttd5eebgmf[95];
  wire o2nfdhz09d    = e4_5otstd9ttd5eebgmf[68];
  wire l6zlxtervy    = e4_5otstd9ttd5eebgmf[69];
  wire mcnugl6b38bsf5    = e4_5otstd9ttd5eebgmf[70];
  wire zvbl_p8a9z    = e4_5otstd9ttd5eebgmf[71];
  wire cdgcsm3vnv1    = e4_5otstd9ttd5eebgmf[72];
  wire m5iytfsnw380oj8    = e4_5otstd9ttd5eebgmf[73];
  wire e2eni70ck7d6     = e4_5otstd9ttd5eebgmf[74 ];
  wire ud802vo0svz2     = e4_5otstd9ttd5eebgmf[75 ];
  wire subovxyhs     = e4_5otstd9ttd5eebgmf[76 ];
  wire a6zk75ptahqc   = e4_5otstd9ttd5eebgmf[77];   
  wire ydcwgy1tbx4w_fb   = e4_5otstd9ttd5eebgmf[78];   
  wire yp4xcxckn5uo5   = e4_5otstd9ttd5eebgmf[79];   
  wire crm5avimdh    = e4_5otstd9ttd5eebgmf[80 ];   
  wire xtb4kjd8ti4    = e4_5otstd9ttd5eebgmf[81 ];   
  wire tvirf9_p_qjq    = e4_5otstd9ttd5eebgmf[82 ];   
  wire dni4x70aj_us6o    = e4_5otstd9ttd5eebgmf[83 ];   
  wire ocdf16j148vr5   = e4_5otstd9ttd5eebgmf[84];   
  wire d8i2e0e5umxqv     = e4_5otstd9ttd5eebgmf[85  ];   
  wire bn_3usiy5s    = e4_5otstd9ttd5eebgmf[86 ];   
  wire ll4ct_hdk57a9    = e4_5otstd9ttd5eebgmf[87 ];   
  wire ethevzph7my   = e4_5otstd9ttd5eebgmf[88];   
  wire xmoo0yw3go8i   = e4_5otstd9ttd5eebgmf[89];   
  wire i_l9_tprh9u0    = e4_5otstd9ttd5eebgmf[90 ];   
  wire hndp_kuba5nlp   = e4_5otstd9ttd5eebgmf[91];   
  wire tmcnfufl_fi42     = e4_5otstd9ttd5eebgmf[92  ];   
  wire vi1b_x4jzofb    = e4_5otstd9ttd5eebgmf[93 ];   
  wire anx2k4uqqlku    = e4_5otstd9ttd5eebgmf[94 ];   





  wire oyxjs3av0z67vqd9z93 = n6izg3jvgts[1];
  wire laksv6w2w3g85egjh = n6izg3jvgts[5];

  wire jj1e19z04mdd1903k6 = n6izg3jvgts[2]; 
  wire obyenny15k41m98a7jhajt = n6izg3jvgts[6]; 

  wire l_mrsjnfjwcw23l = n6izg3jvgts[3]; 
   wire t124x7d61613qbluy3 = n6izg3jvgts[7]; 

  wire xbbag3r7y2il4kz_fdcb =  n6izg3jvgts[4];
  wire chgsl3e3omcgzcmhcdwnd9 =  n6izg3jvgts[8];
  wire hxv8akm9tnbagx = n6izg3jvgts[14];
  wire qhmdzlcppcq8 = n6izg3jvgts[15];
  wire b43ixz6gjo_3lsem91csma = ntp3h6qp | xn1f1pv3xq9j | ksqlq_qg3d; 
  wire i23hpo2hianl9_xpewemf = gqej_k2u1l4m | s7h0yqvmtsxj | wgvga5xo;



  wire ubyk3d30hk8vuj7jjny689v146curyxy = b3sltjkxd | nbcmgtqjii6 | he1npja1q
                                   | o2nfdhz09d | l6zlxtervy | mcnugl6b38bsf5
                                   | a6zk75ptahqc | ydcwgy1tbx4w_fb | yp4xcxckn5uo5
                                   ;
  wire [64-1:0] pcko5kg7h0yh1z = j_rvclhfbeig5cqeb3_ ? nb3w1rq_ny95rvrt : xo5bwsw4j8a;

  wire [1:0]  lokgn5ampy2sq813dph9iluv99z;
  assign lokgn5ampy2sq813dph9iluv99z[0] = e8kmdrlj7pv | y44x7fnhxvoz85;
  assign lokgn5ampy2sq813dph9iluv99z[1] =r1h7wsdxc | akokb5adw5 | mtm0jygbpquyx_ | oi_q1zg22f_j | nhvy44ogg7437 | r_39wh4gt2t15;
  wire [1:0]  nsmvy4s6iv7_wyo2_otdx6ka79;
  assign nsmvy4s6iv7_wyo2_otdx6ka79[0] = e8kmdrlj7pv | y44x7fnhxvoz85;
  assign nsmvy4s6iv7_wyo2_otdx6ka79[1] =r1h7wsdxc | akokb5adw5 | mtm0jygbpquyx_ | oi_q1zg22f_j | nhvy44ogg7437 | r_39wh4gt2t15;

  wire upbbycb5makv3xss7d_ueoxns88bj = n6izg3jvgts[25];
  wire isxv0tqhyam      = n6izg3jvgts[26];
  wire a0qgw4hnfjjkdr_nhqk3i = 
                          h80eeiznk | e14xup9fo8q72 | qz487t2wc1 | edwtafv6h | fqhz535idl
                          | m4ru19tg0 | b9j3bhreofzf | l_rmt2esx6tvr | mku_74ifgnfieu2 | uz5zh9l2ar1q
                          | a1q5p89kjv | hniqik4tqx | i7uhvhnm5dzd0 | yuimu6qrm3 | fj3p9vcal5
                          | znkntww0_qvy0 | o2476dr5c9g | vmjyb2bbjdd1t4
                          | crm5avimdh | xtb4kjd8ti4 | tvirf9_p_qjq
                          | dni4x70aj_us6o | ocdf16j148vr5 | ll4ct_hdk57a9
                          | ethevzph7my | xmoo0yw3go8i | i_l9_tprh9u0
                          | hndp_kuba5nlp | h_aqv6_zs
                          ;

  wire t5r22u8u84ja1kz = e8kmdrlj7pv | y44x7fnhxvoz85 | b3sltjkxd | nbcmgtqjii6 | he1npja1q;

  wire lhe9qqf_zddxeoabsci_jsy2o = hbgz8fj2 | w4hjaq5ha | gddu1322qyclw5;
  wire gnql1wtsvs8lc_ilos7_mf2 = edwtafv6h | fqhz535idl | m4ru19tg0 | b9j3bhreofzf | l_rmt2esx6tvr | mku_74ifgnfieu2 | uz5zh9l2ar1q 
                              | wq_as4te8v_b | ga7v537skbsy | sjjokf_h | yptobqxpymp | n64e5158axn6;
  wire nvbe_d2m8frf6lhejs370g = lm6sobl4jhpz | sdiqw5ujf | w3m1avjrhe;
  wire ci22asx1f0mb9cas2qyhxdbjz7 =  iatq6q6eq | hqgpv7iwel4t | rte1rpxc | scwyr94dp | xu4g6q5o_ | jqjgwcghbu | xpm18ev4bbldh; 
  wire lq2yw3ecpj0d3nv481jxvgb8ocz = e8kmdrlj7pv | y44x7fnhxvoz85 | n4q1xxu4x_3hl | hq5o156te | tdmjh8lo4z5 ;
  wire d3mzo0dhh20fvpjk45g58qkdakf = exe5zfxbfu0_8|y7jlwr4xt5op|tu3h2v18zj|hc_xm8msfc3;
  wire gqdeg_zyb4xaw4ewd8lcc0ppphj = lm0p0_l8v3c | m2p4w1oz_anbe | dc4k61sy3n_z1m | ychqrju9d5fye7j; 
  wire mwbdq5y4q2vm_jjdra48kiwmnhgdmw2o = uu7kphuq | cnluzxjjp1rcx |  jctnij88_5a |  mydhpyzp8hjwy; 
  wire i66_7g0ft50oteolikly2sl  = lq2yw3ecpj0d3nv481jxvgb8ocz 
                               | d3mzo0dhh20fvpjk45g58qkdakf
                               | gqdeg_zyb4xaw4ewd8lcc0ppphj
                               | mwbdq5y4q2vm_jjdra48kiwmnhgdmw2o
                               ;
  wire m1srzg1de1n94hnbvq4vdq = isxv0tqhyam & (~(nvbe_d2m8frf6lhejs370g 
                                              | ci22asx1f0mb9cas2qyhxdbjz7 
                                              | i66_7g0ft50oteolikly2sl 
                                              | a0qgw4hnfjjkdr_nhqk3i 
                                              ));
  wire hf3_u19xhtm47jygm346ih5592f = n6izg3jvgts[28]; 
  wire scmnbmg4dt1z5dy2efq2oclr2rrw = r1h7wsdxc | akokb5adw5 | mtm0jygbpquyx_ | oi_q1zg22f_j
                                   | zt47pxlvcnvwaj | mxh5z6vyj5 | dcd8vqqpxs
                                   | uqitfc00xwe | i3t5mrrybl5 | yptobqxpymp | n64e5158axn6
                                   | wq_as4te8v_b | ga7v537skbsy | sjjokf_h | dr32dt_a9g
                                   | rtuq1m6b67r7u | ig7u5q3yu6kicnh | d1zrh920nh | nhvy44ogg7437
                                   | r_39wh4gt2t15 | m2p4w1oz_anbe | dc4k61sy3n_z1m | ychqrju9d5fye7j
                                   | exe5zfxbfu0_8 | y7jlwr4xt5op | tu3h2v18zj | hc_xm8msfc3
                                   | lm0p0_l8v3c | uu7kphuq | cnluzxjjp1rcx | jctnij88_5a 
                                   | mydhpyzp8hjwy | n4q1xxu4x_3hl | hq5o156te | tdmjh8lo4z5
                                   | iatq6q6eq | hqgpv7iwel4t | rte1rpxc | scwyr94dp
                                   | xu4g6q5o_ | jqjgwcghbu | xpm18ev4bbldh | lm6sobl4jhpz
                                   | sdiqw5ujf | w3m1avjrhe
                                   | zvbl_p8a9z | cdgcsm3vnv1| m5iytfsnw380oj8
                                   | o2nfdhz09d | l6zlxtervy| mcnugl6b38bsf5
                                   | a6zk75ptahqc | ydcwgy1tbx4w_fb| yp4xcxckn5uo5
                                   ;
  wire fwyll5w8ae07xgdgo39mexv4ixjyh2v6h = hf3_u19xhtm47jygm346ih5592f & (~scmnbmg4dt1z5dy2efq2oclr2rrw); 
  wire i326youmut2f1nc3n5g954hksk2i_xk8_ = hf3_u19xhtm47jygm346ih5592f & scmnbmg4dt1z5dy2efq2oclr2rrw; 
  wire l1fkxm0gnih0xhcg05fcz2g9h3q6r0wm7f = ci22asx1f0mb9cas2qyhxdbjz7 & (~scmnbmg4dt1z5dy2efq2oclr2rrw);
  wire dpr2g7tab1p_jkdlwh1uh6f0pk = ci22asx1f0mb9cas2qyhxdbjz7 & scmnbmg4dt1z5dy2efq2oclr2rrw;
  wire nqrawbn8solmf6u8m2qj256f0kiqc = nvbe_d2m8frf6lhejs370g & (~scmnbmg4dt1z5dy2efq2oclr2rrw);
  wire uph5v1440arp4wwekqz3w5epcssoq = nvbe_d2m8frf6lhejs370g & scmnbmg4dt1z5dy2efq2oclr2rrw;
  wire br30p3wqrhus0g438nkl08fe033ge = gnql1wtsvs8lc_ilos7_mf2 & (~scmnbmg4dt1z5dy2efq2oclr2rrw);
  wire ss3dr3dcf16zyxd7vzqkavqcfsg67a = gnql1wtsvs8lc_ilos7_mf2 & scmnbmg4dt1z5dy2efq2oclr2rrw;
  wire q73_mo9ywdxgnaqt5j3bkgy = yptobqxpymp | n64e5158axn6;
  wire yr49c02b6h4zwd =     
                        
                         |m2p4w1oz_anbe |dc4k61sy3n_z1m  |ychqrju9d5fye7j  |lm0p0_l8v3c |uu7kphuq
                         |cnluzxjjp1rcx  |jctnij88_5a    |mydhpyzp8hjwy
                         |iatq6q6eq   |hqgpv7iwel4t 
                         |rte1rpxc   |scwyr94dp   |xu4g6q5o_  |jqjgwcghbu |xpm18ev4bbldh
                         |n4q1xxu4x_3hl   |hq5o156te    |tdmjh8lo4z5
                        
                         |b3sltjkxd |nbcmgtqjii6  |he1npja1q |tu3h2v18zj |exe5zfxbfu0_8 | hc_xm8msfc3 | y7jlwr4xt5op  
                         |a6zk75ptahqc |ydcwgy1tbx4w_fb  |yp4xcxckn5uo5
                        ;
  wire f1fq641fouvrm9yr1i = yuimu6qrm3 | i7uhvhnm5dzd0;
  wire rkd9qofi1kl4toh4 = znkntww0_qvy0 | fj3p9vcal5
                        | crm5avimdh | xtb4kjd8ti4 | tvirf9_p_qjq
                        | d8i2e0e5umxqv  | bn_3usiy5s 
                        | dni4x70aj_us6o | ocdf16j148vr5
                        | ll4ct_hdk57a9 | ethevzph7my | xmoo0yw3go8i 
                        | i_l9_tprh9u0 | hndp_kuba5nlp
                        ;

  parameter uneg70cdsrth1_hntmv = 0;
  parameter vlce4jn2kvx35c3mp = 1;
  parameter vrk4v02ziadwgyqaph8 = 2;
  parameter kcvaxstqpset40tc9xb = 3;
  parameter w8tb5rz6h4lragd143b1 = 4; 
  wire jujbzkikqi6bkoc = d1zrh920nh | ig7u5q3yu6kicnh | y7jlwr4xt5op | hc_xm8msfc3;
  wire tatmybs7ap1zwxm = nhvy44ogg7437 | m2p4w1oz_anbe | ychqrju9d5fye7j | r_39wh4gt2t15;
  wire uwaom12cwzsp48qb4gg5 = rtuq1m6b67r7u;
  wire edgkfsbwss3jeiha5b9 = dr32dt_a9g | cnluzxjjp1rcx;
  wire [3:0] kfgyebl8h3dbx234323 = {edgkfsbwss3jeiha5b9, uwaom12cwzsp48qb4gg5, tatmybs7ap1zwxm, jujbzkikqi6bkoc};

  wire znsowcs8aawt14bwmm7pw028ej = rte1rpxc | scwyr94dp| xu4g6q5o_ | wq_as4te8v_b | ga7v537skbsy | sjjokf_h
                              ;
  wire q41nhsca9cpo8c5nxkf06aiaq9l5rtqk4ewc0 = rte1rpxc | scwyr94dp| xu4g6q5o_ | wq_as4te8v_b | ga7v537skbsy | sjjokf_h
                                        ;
  wire qm58hvuf0bd4w3wh45efr0cm3_hg =  jqjgwcghbu | xpm18ev4bbldh 
                                 | uz5zh9l2ar1q | l_rmt2esx6tvr | mku_74ifgnfieu2 
                                 ;
  wire fk79f3abowqk6mjcsntt5r2yo505028bazs =  jqjgwcghbu | xpm18ev4bbldh;
  wire sm_kcjumavrifsevqbr07v0146ebrc = y44x7fnhxvoz85 | jctnij88_5a | mydhpyzp8hjwy
                                      | edwtafv6h | fqhz535idl | ll4ct_hdk57a9 | ethevzph7my | xmoo0yw3go8i
                                      | tmcnfufl_fi42 | vi1b_x4jzofb | anx2k4uqqlku
                                      ;
  wire wj49kn8i8h4pmijeabgtzdr5_lhgmj4cuthy = jctnij88_5a | mydhpyzp8hjwy;
  wire gjexwhnf55ge45we9zlwto5i_ = yuimu6qrm3 | znkntww0_qvy0 | hniqik4tqx | vmjyb2bbjdd1t4
                                 | i_l9_tprh9u0 | hndp_kuba5nlp
                                 ;

  wire ljwz9swzfae4gwikasz9hr5vo9s_ = y44x7fnhxvoz85 | jctnij88_5a | mydhpyzp8hjwy | hniqik4tqx | znkntww0_qvy0 | yuimu6qrm3 | vmjyb2bbjdd1t4 
                                 | wq_as4te8v_b | sjjokf_h | rte1rpxc | xu4g6q5o_ | jqjgwcghbu | xpm18ev4bbldh
                                 | l_rmt2esx6tvr  | uz5zh9l2ar1q | edwtafv6h | fqhz535idl
                                 | ll4ct_hdk57a9 | tmcnfufl_fi42 | i_l9_tprh9u0 | hndp_kuba5nlp
                                 ;
  wire hsbein0es69cegvi14edf67z = y44x7fnhxvoz85 | jctnij88_5a | mydhpyzp8hjwy | hniqik4tqx | znkntww0_qvy0 | yuimu6qrm3 | vmjyb2bbjdd1t4
                                 | edwtafv6h | fqhz535idl | jqjgwcghbu | xpm18ev4bbldh | scwyr94dp | ga7v537skbsy | mku_74ifgnfieu2
                                 | ll4ct_hdk57a9 | tmcnfufl_fi42 | i_l9_tprh9u0 | hndp_kuba5nlp
                                 ;
  wire w3ac6v7xj7_3r4asx4m1qtd_49 = y44x7fnhxvoz85 | jctnij88_5a | mydhpyzp8hjwy
                                      | ll4ct_hdk57a9 | tmcnfufl_fi42 | i_l9_tprh9u0 | hndp_kuba5nlp
                                      | yuimu6qrm3 | znkntww0_qvy0 | hniqik4tqx | vmjyb2bbjdd1t4
                                      ;
  wire k4hr3kb1bde2oauuy3q90vzs9mk = y44x7fnhxvoz85 | jctnij88_5a | mydhpyzp8hjwy
                                      | ll4ct_hdk57a9 | tmcnfufl_fi42 | i_l9_tprh9u0 | hndp_kuba5nlp
                                      | yuimu6qrm3 | znkntww0_qvy0 | hniqik4tqx | vmjyb2bbjdd1t4
                                      ;
  wire rhgr1_e2xizfvqs2vj0adgzyeb5m4 = gjexwhnf55ge45we9zlwto5i_ | l_rmt2esx6tvr  | uz5zh9l2ar1q
                                | edwtafv6h | fqhz535idl 
                                | ethevzph7my | xmoo0yw3go8i | vi1b_x4jzofb | anx2k4uqqlku
                                ;
  wire h2sx13k_xe6f3u68cqn83xyod4lw6 = gjexwhnf55ge45we9zlwto5i_ | mku_74ifgnfieu2
                                | edwtafv6h | fqhz535idl 
                                | ethevzph7my | xmoo0yw3go8i | vi1b_x4jzofb | anx2k4uqqlku
                                ;
  wire mhjy407z1nazwxp6suqjikjzdvz = gjexwhnf55ge45we9zlwto5i_
                                | ethevzph7my | xmoo0yw3go8i | vi1b_x4jzofb | anx2k4uqqlku
                                ;
  wire jdja1s6u6xg80xifaosyd17it = gjexwhnf55ge45we9zlwto5i_
                                | ethevzph7my | xmoo0yw3go8i | vi1b_x4jzofb | anx2k4uqqlku
                                ;

  wire glz_okqbz0246to0645f_n8ki4m4ou4eg56 =  jctnij88_5a | mydhpyzp8hjwy | jqjgwcghbu | xpm18ev4bbldh | wq_as4te8v_b | sjjokf_h | rte1rpxc | xu4g6q5o_ ;
  wire umek5q7x_wgum07ebg811kbe48aoc0lxusp =  jctnij88_5a | mydhpyzp8hjwy | jqjgwcghbu | xpm18ev4bbldh | scwyr94dp | ga7v537skbsy;
  wire a9el8g68vlgcghrbndp03kmppzv3z2lljnqd =  jctnij88_5a | mydhpyzp8hjwy;
  wire atgnb2938zuik2yjjn0y7l2ns03ay6n326w =  jctnij88_5a | mydhpyzp8hjwy; 
  wire [7:0] l5ufd9cta9ufq6cd7a7r = {
                                     jdja1s6u6xg80xifaosyd17it, mhjy407z1nazwxp6suqjikjzdvz, h2sx13k_xe6f3u68cqn83xyod4lw6, rhgr1_e2xizfvqs2vj0adgzyeb5m4
                                    ,k4hr3kb1bde2oauuy3q90vzs9mk, w3ac6v7xj7_3r4asx4m1qtd_49, hsbein0es69cegvi14edf67z, ljwz9swzfae4gwikasz9hr5vo9s_
                                   };
  wire [3:0] kdd7zbk_2mtjb7hi2ezxsetsb11i00 = {atgnb2938zuik2yjjn0y7l2ns03ay6n326w, a9el8g68vlgcghrbndp03kmppzv3z2lljnqd, 
                                           umek5q7x_wgum07ebg811kbe48aoc0lxusp, glz_okqbz0246to0645f_n8ki4m4ou4eg56};


  wire [4:0] saq0lc9n82nipomxtf8qbwe4ppxxa;
  assign saq0lc9n82nipomxtf8qbwe4ppxxa[0] = mtm0jygbpquyx_ | oi_q1zg22f_j|d1zrh920nh|ig7u5q3yu6kicnh|tu3h2v18zj|exe5zfxbfu0_8|hc_xm8msfc3|y7jlwr4xt5op
                                        | zvbl_p8a9z | cdgcsm3vnv1 | m5iytfsnw380oj8
                                        ;
  assign saq0lc9n82nipomxtf8qbwe4ppxxa[1] = r1h7wsdxc | akokb5adw5|r_39wh4gt2t15|nhvy44ogg7437|lm0p0_l8v3c|dc4k61sy3n_z1m|m2p4w1oz_anbe|ychqrju9d5fye7j;
  assign saq0lc9n82nipomxtf8qbwe4ppxxa[2] = uqitfc00xwe |rtuq1m6b67r7u;
  assign saq0lc9n82nipomxtf8qbwe4ppxxa[3] = i3t5mrrybl5 |dr32dt_a9g|uu7kphuq|cnluzxjjp1rcx|jctnij88_5a|mydhpyzp8hjwy;
  assign saq0lc9n82nipomxtf8qbwe4ppxxa[4] = ~(|saq0lc9n82nipomxtf8qbwe4ppxxa[3:0]);
                                         
                                         
                                         
                                         
                                         
                                         
                                         
                                         
                                         
                                         

wire hfssxn5khy43v3a;
wire ajb17ean3ect1us1;
wire [64-1:0] r8yaegh9ba96e1xa;
wire myn68i_ltybiz;
wire zlnee34lfscldxwt3;
wire t0l90nkbwz79s1q42wap9;
wire dnr9zcx_qdh6g53nn1w;
wire s9dhkac1gv9te6mkan;
wire w1csh43sefsn_8nvmg;
wire dfjomq32ksndlo1aqjznt; 
wire fv9hkqkehb6wk48yj1;
wire u40859qtkt50jkwp04lb;
wire eqg6rkyibf01gty;
wire v7kpw07shxecer5jmti; 
wire f2ky3p7ovwuqwa;
wire [63:0] cf4e81a2boubhxs6z22x;
wire [63:0] d22k4tfhcgdvbq5u1d;
wire [63:0] x0ztyrc8qvou4ss8s2f4p;
wire [63:0] mwznoddeyvujj40zt5lzje3;
wire vqf3_nc_dhkahnygcokxg4jo8mkuq3; 
wire [64+3:0] brn_oq7q18eeqdh;
wire xby1k5c7ixtjcr9ppd9;
wire ejocqibvbev5ibu9f8kdpm;
wire oribprqsoi187_50wv07vj;
wire wticntujbmn7m65pu;
wire ypsxwp1_n11vs652ej7u6anyne;
wire ix6y65ige9etghm_5izamhmitft;
wire ze12zuivp7nb1lrz5ddrrz8_m7r50; 
wire [4-1:0] qbpmsk2;               
wire upak0d1ulubm5kj31p0;
wire xgd98yfjs0wg1vjg;
wire q1xiho2m38dg2no_jw479l;
wire bn3hs_059enxzslhk7;
wire zb7_0qoubehnq5_pbeisyo0v;
wire ddu9petr88tlm28sdlv_a;
wire c05m65au78yv406zviubh21ja;
wire fsv9kaj739xkvpb5ihvn7f;
wire qdpmuly3a8cy2favjid0jvmbti8uznl;
wire rbxu9j6nyq8gd_m7v23k6qyil_7;
wire gpnwd_zd2tkt6d2c3v55_18;
wire wk8ixhma96scwieifpc_tu5suu7;
wire qnresap5l13vb0l9fpg3239b; 
wire z6vd_4woxg18gl39ld535x4p;
wire dzbgqblk3n4f9meoze_5kqt;
wire ssc2jog4ea621jss4q93x2lzvbr9u7z;
wire vgdkw2way6depe9y9xlft2qy_s;
wire bdintq29s9wqs4wl3maq;
wire dzf7_ria7p_gb3ncss2_6rm4j_2p2i;
wire r_ncsbcmokm3vu4u4e4mxha_6nnwu; 
wire bw07fgglb3daiy4zwcx3i; 
wire po6d8hzv709mhrjry7d40bw34;
wire e0sutlsxfldkk2qtrc5zcbaubgsc7;
wire r27dn114subbz1mkpqrh8u_nt;
wire tl1zdy8w4zowrfvngxabhgyryi;
wire y508vkh83pjbiyb4s9gee51;
wire my82zyk_j07wn20ac18;
wire lbvwt_z2shtjwj; 
wire jx5yr6oawedvf6yx9yhxwn; 
wire u9lxxlbiwci218dqtstuzuass;
wire [7:0] t23d5a2_5c3czou9eyx2;
wire [3:0] km_egpxwk5_g_t16kwy31x9;
wire [3:0] ljz5sb430nt2daz;
wire [64-1:0] lex655pvopbg;
wire [64-1:0] qpl4vprbks3eyas;
wire mxwmmibxvjzkawbzq7wln;
wire rwsukdwq5hi04;
wire p49z763fixgor;
wire o9baey2y_w0y;
wire [1:0] z69c2t8z03l1c3m9ksrqsyhps3l2ia9;
wire [1:0] fo0chd_icdt7p603t_pnmu3qmz5;
wire ql35edzw8pm;
wire qm1du4l3;
wire a63upddr;
wire [4:0] neomyeq8kehehvjcv0va7nnnx9q9;

localparam jwxxo5dwz741q1 = 604;
wire [jwxxo5dwz741q1-1:0] w7g88jocpgez2tluuo2;
wire [jwxxo5dwz741q1-1:0] y7p1icoagb3n59fpqnu8im;

    assign w7g88jocpgez2tluuo2 = {
                               t_998ilixet4pdvdkju
                              ,a2o96wlgs_5sqzm2a7ba_
                              ,l7mctsr6ttfp83pl8jo7
                              ,hxv8akm9tnbagx
                              ,oyxjs3av0z67vqd9z93
                              ,b43ixz6gjo_3lsem91csma
                              ,i23hpo2hianl9_xpewemf
                              ,jj1e19z04mdd1903k6
                              ,l_mrsjnfjwcw23l
                              ,xbbag3r7y2il4kz_fdcb 
                              ,laksv6w2w3g85egjh
                              ,obyenny15k41m98a7jhajt
                              ,t124x7d61613qbluy3
                              ,chgsl3e3omcgzcmhcdwnd9 
                              ,usrh37qm6nz8yamj6_h_pmbv5
                              ,mipc_c8bfwk8khoqgtsj65f1f
                              ,pm3m6aucefl9oas0vqgwfm
                              ,yc5f_bw94gu1iari4qpmo269z
                              ,qhmdzlcppcq8
                              ,scmnbmg4dt1z5dy2efq2oclr2rrw 
                              ,xcp0v_slt0baqx9h6px
                              ,znsowcs8aawt14bwmm7pw028ej
                              ,qm58hvuf0bd4w3wh45efr0cm3_hg
                              ,sm_kcjumavrifsevqbr07v0146ebrc 
                              ,gjexwhnf55ge45we9zlwto5i_ 
                              ,q41nhsca9cpo8c5nxkf06aiaq9l5rtqk4ewc0
                              ,fk79f3abowqk6mjcsntt5r2yo505028bazs
                              ,wj49kn8i8h4pmijeabgtzdr5_lhgmj4cuthy 
                              ,jsz4fvx2s3ijb5                
                              ,gdebc5b6o6bv57ax1bw
                              ,lygqe2977b3fd_0eit3wg_nnfirn
                              ,w363n7ci30h3kw2g1oktlj1puysbju
                              ,vz2rm7lc9ctulrdhe1kv8wdmobft
                              ,th583ebkp2cj56crsivefzygk81o65_h2
                              ,hlmhgsbtxsmi7y1a7oshnntydp27pj
                              ,dshcfm3k8zhyftxq_xw9j106j59z7notf
                              ,hf3_u19xhtm47jygm346ih5592f
                              ,fwyll5w8ae07xgdgo39mexv4ixjyh2v6h 
                              ,i326youmut2f1nc3n5g954hksk2i_xk8_ 
                              ,nvbe_d2m8frf6lhejs370g
                              ,nqrawbn8solmf6u8m2qj256f0kiqc
                              ,uph5v1440arp4wwekqz3w5epcssoq
                              ,upbbycb5makv3xss7d_ueoxns88bj
                              ,gnql1wtsvs8lc_ilos7_mf2 
                              ,br30p3wqrhus0g438nkl08fe033ge
                              ,ss3dr3dcf16zyxd7vzqkavqcfsg67a
                              ,ci22asx1f0mb9cas2qyhxdbjz7 
                              ,l1fkxm0gnih0xhcg05fcz2g9h3q6r0wm7f
                              ,dpr2g7tab1p_jkdlwh1uh6f0pk
                              ,m1srzg1de1n94hnbvq4vdq 
                              ,lq2yw3ecpj0d3nv481jxvgb8ocz
                              ,d3mzo0dhh20fvpjk45g58qkdakf
                              ,gqdeg_zyb4xaw4ewd8lcc0ppphj
                              ,mwbdq5y4q2vm_jjdra48kiwmnhgdmw2o
                              ,i66_7g0ft50oteolikly2sl
                              ,a0qgw4hnfjjkdr_nhqk3i 
                              ,t5r22u8u84ja1kz 
                              ,lhe9qqf_zddxeoabsci_jsy2o 
                              ,ubyk3d30hk8vuj7jjny689v146curyxy
                              ,l5ufd9cta9ufq6cd7a7r 
                              ,kdd7zbk_2mtjb7hi2ezxsetsb11i00 
                              ,pcko5kg7h0yh1z    
                              ,amgi_rqhtd007
                              ,kfgyebl8h3dbx234323 
                              ,lokgn5ampy2sq813dph9iluv99z
                              ,nsmvy4s6iv7_wyo2_otdx6ka79
                              ,hbgz8fj2
                              ,jctnij88_5a
                              ,mydhpyzp8hjwy
                              ,q73_mo9ywdxgnaqt5j3bkgy
                              ,yr49c02b6h4zwd
                              ,rkd9qofi1kl4toh4
                              ,f1fq641fouvrm9yr1i 
                              ,saq0lc9n82nipomxtf8qbwe4ppxxa
    };

    assign                  {
                               hfssxn5khy43v3a
                              ,ajb17ean3ect1us1
                              ,r8yaegh9ba96e1xa
                              ,myn68i_ltybiz
                              ,zlnee34lfscldxwt3
                              ,t0l90nkbwz79s1q42wap9
                              ,dnr9zcx_qdh6g53nn1w
                              ,s9dhkac1gv9te6mkan
                              ,w1csh43sefsn_8nvmg
                              ,dfjomq32ksndlo1aqjznt 
                              ,fv9hkqkehb6wk48yj1
                              ,u40859qtkt50jkwp04lb
                              ,eqg6rkyibf01gty
                              ,v7kpw07shxecer5jmti 
                              ,cf4e81a2boubhxs6z22x
                              ,d22k4tfhcgdvbq5u1d
                              ,x0ztyrc8qvou4ss8s2f4p
                              ,mwznoddeyvujj40zt5lzje3
                              ,f2ky3p7ovwuqwa
                              ,vqf3_nc_dhkahnygcokxg4jo8mkuq3 
                              ,brn_oq7q18eeqdh 
                              ,xby1k5c7ixtjcr9ppd9
                              ,ejocqibvbev5ibu9f8kdpm
                              ,oribprqsoi187_50wv07vj 
                              ,wticntujbmn7m65pu 
                              ,ypsxwp1_n11vs652ej7u6anyne
                              ,ix6y65ige9etghm_5izamhmitft
                              ,ze12zuivp7nb1lrz5ddrrz8_m7r50 
                              ,qbpmsk2                
                              ,upak0d1ulubm5kj31p0
                              ,xgd98yfjs0wg1vjg
                              ,q1xiho2m38dg2no_jw479l
                              ,bn3hs_059enxzslhk7
                              ,zb7_0qoubehnq5_pbeisyo0v
                              ,ddu9petr88tlm28sdlv_a
                              ,c05m65au78yv406zviubh21ja
                              ,fsv9kaj739xkvpb5ihvn7f
                              ,qdpmuly3a8cy2favjid0jvmbti8uznl 
                              ,rbxu9j6nyq8gd_m7v23k6qyil_7 
                              ,gpnwd_zd2tkt6d2c3v55_18
                              ,wk8ixhma96scwieifpc_tu5suu7
                              ,qnresap5l13vb0l9fpg3239b
                              ,z6vd_4woxg18gl39ld535x4p
                              ,dzbgqblk3n4f9meoze_5kqt 
                              ,ssc2jog4ea621jss4q93x2lzvbr9u7z
                              ,vgdkw2way6depe9y9xlft2qy_s
                              ,bdintq29s9wqs4wl3maq 
                              ,dzf7_ria7p_gb3ncss2_6rm4j_2p2i
                              ,r_ncsbcmokm3vu4u4e4mxha_6nnwu 
                              ,bw07fgglb3daiy4zwcx3i 
                              ,po6d8hzv709mhrjry7d40bw34
                              ,e0sutlsxfldkk2qtrc5zcbaubgsc7
                              ,r27dn114subbz1mkpqrh8u_nt
                              ,tl1zdy8w4zowrfvngxabhgyryi
                              ,y508vkh83pjbiyb4s9gee51
                              ,my82zyk_j07wn20ac18 
                              ,lbvwt_z2shtjwj 
                              ,jx5yr6oawedvf6yx9yhxwn 
                              ,u9lxxlbiwci218dqtstuzuass
                              ,t23d5a2_5c3czou9eyx2 
                              ,km_egpxwk5_g_t16kwy31x9 
                              ,lex655pvopbg    
                              ,qpl4vprbks3eyas    
                              ,ljz5sb430nt2daz 
                              ,z69c2t8z03l1c3m9ksrqsyhps3l2ia9
                              ,fo0chd_icdt7p603t_pnmu3qmz5
                              ,ql35edzw8pm
                              ,qm1du4l3
                              ,a63upddr
                              ,mxwmmibxvjzkawbzq7wln
                              ,rwsukdwq5hi04
                              ,p49z763fixgor
                              ,o9baey2y_w0y 
                              ,neomyeq8kehehvjcv0va7nnnx9q9
                             } = y7p1icoagb3n59fpqnu8im;


wire  wjblnj3zxv26betgtpwtxz85mlz;
assign izj2me9tmzxitrpzl1tr = pzhh8hyzbdb80ac8sdd_49 & wjblnj3zxv26betgtpwtxz85mlz;
wire   mxeyuvtl7iodvi9lm7qutkla = tvdvyldvwqhx7g8r9di & pzhh8hyzbdb80ac8sdd_49;
assign rgcs7q5ke7h8fte8jecm = tvdvyldvwqhx7g8r9di & wjblnj3zxv26betgtpwtxz85mlz;
 ux607_gnrl_pipe_stage # (
  .CUT_READY(0),
  .DP(1),
  .DW(jwxxo5dwz741q1)
 ) if1uo6nwhd78_9scnac (
   .i_vld(mxeyuvtl7iodvi9lm7qutkla), 
   .i_rdy(wjblnj3zxv26betgtpwtxz85mlz), 
   .i_dat(w7g88jocpgez2tluuo2  ),
   .o_vld(cwmxezrc3jv6hzxcfc), 
   .o_rdy(uig3ujuyq0_61kqb), 
   .o_dat(y7p1icoagb3n59fpqnu8im),
 
   .clk  (gf33atgy  ),
   .rst_n(ru_wi)  
  );



wire royh8kfx4l6z206rgv;
wire [64-1:0] cmdsrflujxwd007q;

lxot_pmljpjs9pco4am4pfh5r xrytmm0lw1o2u5xbyc8ppi72s7(
     .oyxjs3av0z67vqd9z93             (zlnee34lfscldxwt3) ,
     .laksv6w2w3g85egjh           (fv9hkqkehb6wk48yj1),
     .jj1e19z04mdd1903k6            (s9dhkac1gv9te6mkan),
     .obyenny15k41m98a7jhajt          (u40859qtkt50jkwp04lb),
     .b43ixz6gjo_3lsem91csma      (t0l90nkbwz79s1q42wap9),
     .i23hpo2hianl9_xpewemf      (dnr9zcx_qdh6g53nn1w),
     .l_mrsjnfjwcw23l            (w1csh43sefsn_8nvmg),
     .xbbag3r7y2il4kz_fdcb        (dfjomq32ksndlo1aqjznt),
     .t124x7d61613qbluy3          (eqg6rkyibf01gty),
     .chgsl3e3omcgzcmhcdwnd9      (v7kpw07shxecer5jmti),
     .usrh37qm6nz8yamj6_h_pmbv5       (cf4e81a2boubhxs6z22x),
     .mipc_c8bfwk8khoqgtsj65f1f       (d22k4tfhcgdvbq5u1d),
     .pm3m6aucefl9oas0vqgwfm       (x0ztyrc8qvou4ss8s2f4p),
     .yc5f_bw94gu1iari4qpmo269z       (mwznoddeyvujj40zt5lzje3),
     .k6c8aiwomjglm9ok9zt4wb        (cmdsrflujxwd007q), 
     .etcizv32c63_xdl3f60          (royh8kfx4l6z206rgv ) 
);



 
  wire deio5fy869cl5z0kt   = q1xiho2m38dg2no_jw479l | xgd98yfjs0wg1vjg; 
  wire ha5_nthmqq8a1b3 = zb7_0qoubehnq5_pbeisyo0v | bn3hs_059enxzslhk7; 
  wire [63:0] v4wb_ti29jdb4ieh7s5x321jdjg0hh5c = u9lxxlbiwci218dqtstuzuass ? {32'b0,32'h7fffffff} : {17'b0,32'h7fffffff,15'b0};
  wire c2w073rogzl = gpnwd_zd2tkt6d2c3v55_18 | bdintq29s9wqs4wl3maq |  y508vkh83pjbiyb4s9gee51 | bw07fgglb3daiy4zwcx3i;
  wire xb965l0fnqcjd = c2w073rogzl  & vqf3_nc_dhkahnygcokxg4jo8mkuq3 ;
  wire h16j5g6h4qze_20ud9ix = upak0d1ulubm5kj31p0 & lex655pvopbg [31];
  wire cqycxk2rfiyv2uf7m5a3o0u = upak0d1ulubm5kj31p0 & lex655pvopbg [63];
  wire zmxck2ys1tqf6aio41lqxzhzor = d22k4tfhcgdvbq5u1d[63];
  wire [63:0] v37ldix2i_j_gihlsim = {{32{h16j5g6h4qze_20ud9ix}}, lex655pvopbg[31:0]};
  wire [63:0] nwahql0hdil255akcnj02n = {{32{cqycxk2rfiyv2uf7m5a3o0u}}, lex655pvopbg[63:32]};
  wire [63:0] ppy6fe856k1_rda    =  ({64{gpnwd_zd2tkt6d2c3v55_18 | bdintq29s9wqs4wl3maq 
                                         | bw07fgglb3daiy4zwcx3i | po6d8hzv709mhrjry7d40bw34}} & v37ldix2i_j_gihlsim)
                                   |  ({64{e0sutlsxfldkk2qtrc5zcbaubgsc7}} & {v37ldix2i_j_gihlsim[48:0],15'b0})
                                   |  ({64{r27dn114subbz1mkpqrh8u_nt}} & {v37ldix2i_j_gihlsim[47:0],16'b0})
                                   |  ({64{tl1zdy8w4zowrfvngxabhgyryi}} & {v37ldix2i_j_gihlsim[31:0],32'b0})
                                   ;
  wire [63:0] js993ji4rw4f0iywaz7ozrkxnz =  ({64{gpnwd_zd2tkt6d2c3v55_18 | bdintq29s9wqs4wl3maq 
                                         | bw07fgglb3daiy4zwcx3i | po6d8hzv709mhrjry7d40bw34}} & nwahql0hdil255akcnj02n)
                                   |  ({64{e0sutlsxfldkk2qtrc5zcbaubgsc7}} & {nwahql0hdil255akcnj02n[48:0],15'b0})
                                   |  ({64{r27dn114subbz1mkpqrh8u_nt}} & {nwahql0hdil255akcnj02n[47:0],16'b0})
                                   |  ({64{tl1zdy8w4zowrfvngxabhgyryi}} & {nwahql0hdil255akcnj02n[31:0],32'b0})
                                   ;

  wire [32:0] e4gxec3zjbv25o5rf8wai1do = xgd98yfjs0wg1vjg ? {1'b0,v4wb_ti29jdb4ieh7s5x321jdjg0hh5c[31:0]}   : {1'b0,cf4e81a2boubhxs6z22x[31:0] };
  wire [32:0] br3rbue4woi7_rety29v2ku0yi = xgd98yfjs0wg1vjg ? 33'b0 : {(upak0d1ulubm5kj31p0 & cf4e81a2boubhxs6z22x[63]),cf4e81a2boubhxs6z22x[63:32]};
  wire [32:0] y5tou6wv8wpsep2d7nvz2 = xgd98yfjs0wg1vjg ? 33'b0 : {(upak0d1ulubm5kj31p0 & d22k4tfhcgdvbq5u1d[31]),d22k4tfhcgdvbq5u1d[31:0] };
  wire [32:0] b9s062tfzpxix6i364q8997ve = xgd98yfjs0wg1vjg ? {1'b0,v4wb_ti29jdb4ieh7s5x321jdjg0hh5c[63:32]}: {(upak0d1ulubm5kj31p0 & d22k4tfhcgdvbq5u1d[63]),d22k4tfhcgdvbq5u1d[63:32]};
  wire [32:0] ka97f3isuhin5zjf537_xzb4l = bn3hs_059enxzslhk7 ? {1'b0,v4wb_ti29jdb4ieh7s5x321jdjg0hh5c[31:0]}   : {1'b0,x0ztyrc8qvou4ss8s2f4p[31:0] };
  wire [32:0] qfqtz2j7nx_vphe1s9mq8lvb_ = bn3hs_059enxzslhk7 ? 33'b0 : {(upak0d1ulubm5kj31p0 & x0ztyrc8qvou4ss8s2f4p[63]),x0ztyrc8qvou4ss8s2f4p[63:32]};
  wire [32:0] xb2vqfv1me2hqy9bovai5uro = bn3hs_059enxzslhk7 ? 33'b0 : {(upak0d1ulubm5kj31p0 & mwznoddeyvujj40zt5lzje3[31]),mwznoddeyvujj40zt5lzje3[31:0] };
  wire [32:0] gb2x6jead6bokztqfctlgihone = bn3hs_059enxzslhk7 ? {1'b0,v4wb_ti29jdb4ieh7s5x321jdjg0hh5c[63:32]}: {(upak0d1ulubm5kj31p0 & mwznoddeyvujj40zt5lzje3[63]),mwznoddeyvujj40zt5lzje3[63:32]};
  wire [63:0] ppccyfh77m_wis5 =  cf4e81a2boubhxs6z22x;
  wire [63:0] gv8wbubo_bik7kj = d22k4tfhcgdvbq5u1d;

  wire [32:0] hplpy12njwr2n5atmn6x5qq9 = 33'b0;
  wire [32:0] sp8bh60rd8y0rg63n_iy1omu = ({33{z69c2t8z03l1c3m9ksrqsyhps3l2ia9[0]}} & {17'h1ffff,16'h0});
  wire [32:0] qkojw9k46swimy74csh3u8vk6te = ({33{z69c2t8z03l1c3m9ksrqsyhps3l2ia9[0]}} & {17'h1ffff,16'h0});
  wire [32:0] og2hab4t9g5bja_lhgqdyf_ = ({33{z69c2t8z03l1c3m9ksrqsyhps3l2ia9[1]}} & {17'h1ffff,16'h0})
                                     | ({33{z69c2t8z03l1c3m9ksrqsyhps3l2ia9[0]}} & 33'h1ffffffff)
                                     ;
  wire [32:0] bbs_zs12hm1yzwvyi6ouup8f = 33'b0;
  wire [32:0] y1y6hyewgqgll1127wp043 = ({33{fo0chd_icdt7p603t_pnmu3qmz5[0]}} & {17'h1ffff,16'h0});
  wire [32:0] pf6tyxmf2miiw2uhxk0mzwtn0eb = ({33{fo0chd_icdt7p603t_pnmu3qmz5[0]}} & {17'h1ffff,16'h0});
  wire [32:0] x6ob94k6ng8guck7udbs5n1 = ({33{fo0chd_icdt7p603t_pnmu3qmz5[1]}} & {17'h1ffff,16'h0})
                                     | ({33{fo0chd_icdt7p603t_pnmu3qmz5[0]}} & 33'h1ffffffff)
                                     ;

  wire [32:0] s9e3pj73edsa2hn8i_ = (~hplpy12njwr2n5atmn6x5qq9) & e4gxec3zjbv25o5rf8wai1do;
  wire [32:0] ownboagykdrscrtsqd9p = (~sp8bh60rd8y0rg63n_iy1omu) & br3rbue4woi7_rety29v2ku0yi;
  wire [32:0] fx3o1jdmucfaay24ofp = (~qkojw9k46swimy74csh3u8vk6te) & y5tou6wv8wpsep2d7nvz2;
  wire [32:0] q_zvoz2dbvlqcz57g = (~og2hab4t9g5bja_lhgqdyf_) & b9s062tfzpxix6i364q8997ve;
  wire [32:0] nmm1mrkr7bp3gn3bi = (~bbs_zs12hm1yzwvyi6ouup8f) & ka97f3isuhin5zjf537_xzb4l;
  wire [32:0] zd160q5aoqunimwla4j = (~y1y6hyewgqgll1127wp043) & qfqtz2j7nx_vphe1s9mq8lvb_;
  wire [32:0] d6f56s081ckjmdip0wg9bo = (~pf6tyxmf2miiw2uhxk0mzwtn0eb) & xb2vqfv1me2hqy9bovai5uro;
  wire [32:0] yjwjuu_4_eojh71_wp7v9h = (~x6ob94k6ng8guck7udbs5n1) & gb2x6jead6bokztqfctlgihone;


  
  
  wire [33:0] vu_6ed56hxoy_ = 
                                      ({34{ljz5sb430nt2daz[uneg70cdsrth1_hntmv]}} & {19'b0,1'b1,14'b0})
                                    | ({34{ljz5sb430nt2daz[vlce4jn2kvx35c3mp]}} & {18'b0,1'b1,15'b0})
                                    | ({34{ljz5sb430nt2daz[vrk4v02ziadwgyqaph8]}} & {3'b0,1'b1,30'b0})
                                    | ({34{ljz5sb430nt2daz[kcvaxstqpset40tc9xb]}} & {2'b0,1'b1,31'b0}) 
                                    | ({34{a63upddr}} & (34'h7fffffff))
                                    | ({34{qm1du4l3}} & {2'b0,32'hffffffff})
                                    ;

  wire [64:0] a2yt83mznut1_0e = ({65{fsv9kaj739xkvpb5ihvn7f}} & {{32{s9e3pj73edsa2hn8i_[32]}}, s9e3pj73edsa2hn8i_})
                                | ({65{bdintq29s9wqs4wl3maq | dzbgqblk3n4f9meoze_5kqt}} & {{33{upak0d1ulubm5kj31p0 & ppccyfh77m_wis5[31]}}, ppccyfh77m_wis5[31:0]})
                                | ({65{gpnwd_zd2tkt6d2c3v55_18}} & {{49{upak0d1ulubm5kj31p0 & ppccyfh77m_wis5[15]}}, ppccyfh77m_wis5[15:0]})
                                | ({65{z6vd_4woxg18gl39ld535x4p}} & {57'b0, brn_oq7q18eeqdh[7:0]})
                                ;
  wire [64:0] s07o1zmeybz9jboy5 = ({65{fsv9kaj739xkvpb5ihvn7f}} & {{16{ownboagykdrscrtsqd9p[32]}}, ownboagykdrscrtsqd9p, 16'b0}) 
                                | ({65{bdintq29s9wqs4wl3maq | dzbgqblk3n4f9meoze_5kqt}} & {{33{upak0d1ulubm5kj31p0 & ppccyfh77m_wis5[63]}}, ppccyfh77m_wis5[63:32]})
                                | ({65{gpnwd_zd2tkt6d2c3v55_18}} & {{49{upak0d1ulubm5kj31p0 & ppccyfh77m_wis5[31]}}, ppccyfh77m_wis5[31:16]})
                                | ({65{z6vd_4woxg18gl39ld535x4p}} & {57'b0, brn_oq7q18eeqdh[15:8]})
                                ;
  wire [64:0] r4d0t4rij_pmo8z = ({65{fsv9kaj739xkvpb5ihvn7f}} & {{16{fx3o1jdmucfaay24ofp[32]}}, fx3o1jdmucfaay24ofp, 16'b0}) 
                                | ({65{gpnwd_zd2tkt6d2c3v55_18}} & {{49{upak0d1ulubm5kj31p0 & ppccyfh77m_wis5[47]}}, ppccyfh77m_wis5[47:32]})
                                | ({65{z6vd_4woxg18gl39ld535x4p}} & {57'b0, brn_oq7q18eeqdh[23:16]})
                                ;
  wire [64:0] t2664jbiy_07vcj = ({65{(fsv9kaj739xkvpb5ihvn7f)}} & {q_zvoz2dbvlqcz57g, 32'b0})
                                | ({65{gpnwd_zd2tkt6d2c3v55_18}} & {{49{upak0d1ulubm5kj31p0 & ppccyfh77m_wis5[63]}}, ppccyfh77m_wis5[63:48]})
                                | ({65{z6vd_4woxg18gl39ld535x4p}} & {57'b0, brn_oq7q18eeqdh[31:24]})
                                ;
  wire [64:0] giwetg9prnn_pkn6n = ({65{qdpmuly3a8cy2favjid0jvmbti8uznl }} & {{32{nmm1mrkr7bp3gn3bi[32]}}, nmm1mrkr7bp3gn3bi})
                                | ({65{dzf7_ria7p_gb3ncss2_6rm4j_2p2i | ssc2jog4ea621jss4q93x2lzvbr9u7z}} & {{33{upak0d1ulubm5kj31p0 & gv8wbubo_bik7kj[31]}}, gv8wbubo_bik7kj[31:0]})
                                | ({65{wk8ixhma96scwieifpc_tu5suu7}} & {{49{upak0d1ulubm5kj31p0 & gv8wbubo_bik7kj[15]}}, gv8wbubo_bik7kj[15:0]})
                                | ({65{z6vd_4woxg18gl39ld535x4p}} & {57'b0, brn_oq7q18eeqdh[39:32]})
                                ;
  wire [64:0] f2ehiqbtbjxg4y9 = ({65{qdpmuly3a8cy2favjid0jvmbti8uznl }} & {{16{zd160q5aoqunimwla4j[32]}}, zd160q5aoqunimwla4j, 16'b0}) 
                                | ({65{dzf7_ria7p_gb3ncss2_6rm4j_2p2i | ssc2jog4ea621jss4q93x2lzvbr9u7z}} & {{33{upak0d1ulubm5kj31p0 & gv8wbubo_bik7kj[63]}}, gv8wbubo_bik7kj[63:32]})
                                | ({65{wk8ixhma96scwieifpc_tu5suu7}} & {{49{upak0d1ulubm5kj31p0 & gv8wbubo_bik7kj[31]}}, gv8wbubo_bik7kj[31:16]})
                                | ({65{z6vd_4woxg18gl39ld535x4p}} & {57'b0, brn_oq7q18eeqdh[47:40]})
                                ;
  wire [64:0] fn2pawdixwjekf8fx5m7 = ({65{qdpmuly3a8cy2favjid0jvmbti8uznl }} & {{16{d6f56s081ckjmdip0wg9bo[32]}}, d6f56s081ckjmdip0wg9bo, 16'b0}) 
                                | ({65{wk8ixhma96scwieifpc_tu5suu7}} & {{49{upak0d1ulubm5kj31p0 & gv8wbubo_bik7kj[47]}}, gv8wbubo_bik7kj[47:32]})
                                | ({65{z6vd_4woxg18gl39ld535x4p}} & {57'b0, brn_oq7q18eeqdh[55:48]})
                                ;
  wire [64:0] exrj57dd1ydis6e = ({65{(qdpmuly3a8cy2favjid0jvmbti8uznl )}} & {yjwjuu_4_eojh71_wp7v9h, 32'b0})
                                | ({65{wk8ixhma96scwieifpc_tu5suu7}} & {{49{upak0d1ulubm5kj31p0 & gv8wbubo_bik7kj[63]}}, gv8wbubo_bik7kj[63:48]})
                                | ({65{z6vd_4woxg18gl39ld535x4p}} & {57'b0, brn_oq7q18eeqdh[63:56]})
                                ;
  wire [64:0] cgj8zznqs9_rs4vig8ladd7r = 65'b0;
  wire [64:0] hjwsds5xurs0hi_i85wc8a0 = 65'b0;
  wire [64:0] khklv6b9bmk2wx5r690vq4eq = 65'b0;
  wire [64:0] r754ox21een4i0cwj3236klex3a = 65'b0;
  wire [64:0] p_tiyp08xvouxfizm5t9r8 = ({65{rbxu9j6nyq8gd_m7v23k6qyil_7}} & {{32{nmm1mrkr7bp3gn3bi[32]}}, nmm1mrkr7bp3gn3bi})
                                | ({65{r_ncsbcmokm3vu4u4e4mxha_6nnwu | vgdkw2way6depe9y9xlft2qy_s}} & {{33{upak0d1ulubm5kj31p0 & gv8wbubo_bik7kj[31]}}, gv8wbubo_bik7kj[31:0]})
                                | ({65{qnresap5l13vb0l9fpg3239b}} & {{49{upak0d1ulubm5kj31p0 & gv8wbubo_bik7kj[15]}}, gv8wbubo_bik7kj[15:0]})
                                ;
  wire [64:0] f2gsnr9qfeecwca292lnku227 = ({65{rbxu9j6nyq8gd_m7v23k6qyil_7}} & {{16{zd160q5aoqunimwla4j[32]}}, zd160q5aoqunimwla4j, 16'b0}) 
                                | ({65{r_ncsbcmokm3vu4u4e4mxha_6nnwu | vgdkw2way6depe9y9xlft2qy_s}} & {{33{upak0d1ulubm5kj31p0 & gv8wbubo_bik7kj[63]}}, gv8wbubo_bik7kj[63:32]})
                                | ({65{qnresap5l13vb0l9fpg3239b}} & {{49{upak0d1ulubm5kj31p0 & gv8wbubo_bik7kj[31]}}, gv8wbubo_bik7kj[31:16]})
                                ;
  wire [64:0] ymmuidv3lbgpkx1ioh2kvp6l0y9 = ({65{rbxu9j6nyq8gd_m7v23k6qyil_7}} & {{16{d6f56s081ckjmdip0wg9bo[32]}}, d6f56s081ckjmdip0wg9bo, 16'b0}) 
                                | ({65{qnresap5l13vb0l9fpg3239b}} & {{49{upak0d1ulubm5kj31p0 & gv8wbubo_bik7kj[47]}}, gv8wbubo_bik7kj[47:32]})
                                ;
  wire [64:0] kvvjjve90m_n0ob9ara8pl = ({65{(rbxu9j6nyq8gd_m7v23k6qyil_7)}} & {yjwjuu_4_eojh71_wp7v9h, 32'b0})
                                | ({65{qnresap5l13vb0l9fpg3239b}} & {{49{upak0d1ulubm5kj31p0 & gv8wbubo_bik7kj[63]}}, gv8wbubo_bik7kj[63:48]})
                                ;
  wire indrji2q4p5ysbyc4ynor6ckc = t23d5a2_5c3czou9eyx2[0];
  wire smvhlyuq50g5ld5o6fj_qg = t23d5a2_5c3czou9eyx2[1];
  wire aqooyt2h952qunj08gbwa6 = t23d5a2_5c3czou9eyx2[2];
  wire miz7vhxylfl1_5pztf7tvdt = t23d5a2_5c3czou9eyx2[3];
  wire c66i3cfpsq7jkgu046yc_y = t23d5a2_5c3czou9eyx2[4];
  wire pxdgia8y6_s1m9_el8mgxg7 = t23d5a2_5c3czou9eyx2[5];
  wire mzypp3mzj0ujf_0ae3jxd = t23d5a2_5c3czou9eyx2[6];
  wire fuqfaq7wca9i0qix4qjsd = t23d5a2_5c3czou9eyx2[7];
  wire k2uwwh6g_7ege_it5w25l5hpjnlt = km_egpxwk5_g_t16kwy31x9[0];
  wire iw4x95o42r6pym0mvgcz5s4g5r597_y2 = km_egpxwk5_g_t16kwy31x9[1];
  wire nam6ou62takz82lrg7_1dvl53ekw = km_egpxwk5_g_t16kwy31x9[2];
  wire ot9r5h3f2snedshy4f4gcubnbewl = km_egpxwk5_g_t16kwy31x9[3];

  wire [63:0] zdflw28wxlss1vaq    = 
                                     ({64{ql35edzw8pm}}    & {qpl4vprbks3eyas})
                                    |({64{my82zyk_j07wn20ac18}} & lex655pvopbg)
                                    |({64{c2w073rogzl}} & {ppy6fe856k1_rda})
                                    ;
  wire [64:0] yk90y6l5d_cln9qkt =  {(upak0d1ulubm5kj31p0 & zdflw28wxlss1vaq[63]), zdflw28wxlss1vaq}; 
  wire [64:0] wb0um2oh903cf4gl = indrji2q4p5ysbyc4ynor6ckc ?  (~a2yt83mznut1_0e) : a2yt83mznut1_0e; 
  wire [64:0] bmhyj5vzy18r_ = smvhlyuq50g5ld5o6fj_qg ?  (~s07o1zmeybz9jboy5) : s07o1zmeybz9jboy5; 
  wire [64:0] li1txsi8gtc6 = aqooyt2h952qunj08gbwa6 ?  (~r4d0t4rij_pmo8z) : r4d0t4rij_pmo8z; 
  wire [64:0] jz7v41221fbhg = miz7vhxylfl1_5pztf7tvdt ?  (~t2664jbiy_07vcj) : t2664jbiy_07vcj; 
  wire [64:0] a9dk06q6nvg9bwjh = c66i3cfpsq7jkgu046yc_y ?  (~giwetg9prnn_pkn6n) : giwetg9prnn_pkn6n; 
  wire [64:0] c2f1e9sa022qp = pxdgia8y6_s1m9_el8mgxg7 ?  (~f2ehiqbtbjxg4y9) : f2ehiqbtbjxg4y9; 
  wire [64:0] j826amcloaye9z2zu = mzypp3mzj0ujf_0ae3jxd ?  (~fn2pawdixwjekf8fx5m7) : fn2pawdixwjekf8fx5m7; 
  wire [64:0] kw5ya9ro03kb4 = fuqfaq7wca9i0qix4qjsd ?  (~exrj57dd1ydis6e) : exrj57dd1ydis6e; 

  wire [63:0] rltcqngg8fkiy0nyt3u1kp0ig0t = ({64{xb965l0fnqcjd}} & {js993ji4rw4f0iywaz7ozrkxnz});
  wire [64:0] szz25lqlbfjr_1do40m_nu =  {(upak0d1ulubm5kj31p0 & rltcqngg8fkiy0nyt3u1kp0ig0t[63]), rltcqngg8fkiy0nyt3u1kp0ig0t}; 
  wire [64:0] ofaynbeg20l468n550bzr = 65'b0;
  wire [64:0] t_a7piunj72_ruymfveo = 65'b0;
  wire [64:0] a7bsg64noz2hzrcvy5_fyxx = 65'b0;
  wire [64:0] tlftjsdq0om1ij7yvi74q8 = 65'b0;
  wire [64:0] zp4oxmmrtd0jm6xmpu9exo07 = k2uwwh6g_7ege_it5w25l5hpjnlt ?  (~p_tiyp08xvouxfizm5t9r8) : p_tiyp08xvouxfizm5t9r8; 
  wire [64:0] w9pgray5cmbdb83rsvyu = iw4x95o42r6pym0mvgcz5s4g5r597_y2 ?  (~f2gsnr9qfeecwca292lnku227) : f2gsnr9qfeecwca292lnku227; 
  wire [64:0] aq55569spbv4o2f0j2iv_orw = nam6ou62takz82lrg7_1dvl53ekw ?  (~ymmuidv3lbgpkx1ioh2kvp6l0y9) : ymmuidv3lbgpkx1ioh2kvp6l0y9; 
  wire [64:0] dyl1osrbprq47ppt60zx1zw = ot9r5h3f2snedshy4f4gcubnbewl ?  (~kvvjjve90m_n0ob9ara8pl) : kvvjjve90m_n0ob9ara8pl; 
  wire [33:0] psh56cjgmkcgxminibqe    = deio5fy869cl5z0kt ? 34'b0 : vu_6ed56hxoy_;
  wire [33:0] w4zf9xctmenumbjjuqcxbpe3jw    = ha5_nthmqq8a1b3 ? 34'b0 : vu_6ed56hxoy_;
  wire [34:0]  fvq8btmrm7czfzb9ag_8d89tn = 
                           ({35{xby1k5c7ixtjcr9ppd9}} & 35'd1)
                         | ({35{ejocqibvbev5ibu9f8kdpm}} & 35'd2)
                         | ({35{oribprqsoi187_50wv07vj}} & {35'd4})
                         | ({35{wticntujbmn7m65pu}} & {35'd8})
                         | ({35{z6vd_4woxg18gl39ld535x4p}} & {31'd0,brn_oq7q18eeqdh[64+3:64]})
                         ;
  wire [34:0]  gzddmt2dswaw7jvitpe5hgt61zb255 = 
                           ({35{ypsxwp1_n11vs652ej7u6anyne}} & 35'd1)
                         | ({35{ix6y65ige9etghm_5izamhmitft}} & 35'd2)
                         | ({35{ze12zuivp7nb1lrz5ddrrz8_m7r50}} & {35'd4})
                         ;
  wire [66:0] of41hddih6s4bcn_3nwrp9;
  wire [66:0] mqn5zl56qb4wkr4l5wjwjajufy9;

cwe8y4czjwvbx6znvqv5wg09qsfw i4ftq_qev5t1f_ic3jp0xba83b(
  .ho7hbln__5mzkxd(yk90y6l5d_cln9qkt ),
  .e7e6yf3rwo5s(wb0um2oh903cf4gl ),
  .zpa9wht92mu(bmhyj5vzy18r_ ),
  .mx84o3rvy8(li1txsi8gtc6 ),
  .l6dri5njf3xti3j(jz7v41221fbhg ),
  .d986vh8a8wdpib0(a9dk06q6nvg9bwjh ),
  .xfnf1gelth(c2f1e9sa022qp ),
  .n2t6qssk9yjxv(j826amcloaye9z2zu ),
  .nvjphm8kit9(kw5ya9ro03kb4 ),
  .yj4jcdxd_qu6m3mon       (psh56cjgmkcgxminibqe    ),
  .af86r5akqaznjghqqft (fvq8btmrm7czfzb9ag_8d89tn),
  .wrcjvt7pl1j_           (of41hddih6s4bcn_3nwrp9)
);

cwe8y4czjwvbx6znvqv5wg09qsfw jb4h4rd2igitfd_nsl80g_6l5wf_8cqtf16(
  .ho7hbln__5mzkxd(szz25lqlbfjr_1do40m_nu ),
  .e7e6yf3rwo5s(ofaynbeg20l468n550bzr ),
  .zpa9wht92mu(t_a7piunj72_ruymfveo ),
  .mx84o3rvy8(a7bsg64noz2hzrcvy5_fyxx ),
  .l6dri5njf3xti3j(tlftjsdq0om1ij7yvi74q8 ),
  .d986vh8a8wdpib0(zp4oxmmrtd0jm6xmpu9exo07 ),
  .xfnf1gelth(w9pgray5cmbdb83rsvyu ),
  .n2t6qssk9yjxv(aq55569spbv4o2f0j2iv_orw ),
  .nvjphm8kit9(dyl1osrbprq47ppt60zx1zw ),
  .yj4jcdxd_qu6m3mon       (w4zf9xctmenumbjjuqcxbpe3jw    ),
  .af86r5akqaznjghqqft (gzddmt2dswaw7jvitpe5hgt61zb255),
  .wrcjvt7pl1j_           (mqn5zl56qb4wkr4l5wjwjajufy9)
);



  assign xc2becmsn4fcniw6ks = 1'b0;
                                               
  wire [32:0] dl7jvynj91yjq_ubriyt8rb5y1ksoen = 
                                           ({33{neomyeq8kehehvjcv0va7nnnx9q9[0]}} & of41hddih6s4bcn_3nwrp9[47:15])
                                         | ({33{neomyeq8kehehvjcv0va7nnnx9q9[1]}} & of41hddih6s4bcn_3nwrp9[48:16])
                                         | ({33{neomyeq8kehehvjcv0va7nnnx9q9[2]}} & of41hddih6s4bcn_3nwrp9[63:31])
                                         | ({33{neomyeq8kehehvjcv0va7nnnx9q9[3]}} & of41hddih6s4bcn_3nwrp9[64:32])
                                         | ({33{neomyeq8kehehvjcv0va7nnnx9q9[4]}} & of41hddih6s4bcn_3nwrp9[32:0])
                                         ;
  wire [32:0] g4o3eqh6nb2enoez45n88_wji8vd4 = 
                                           vqf3_nc_dhkahnygcokxg4jo8mkuq3 ? 
                                           ( ({33{neomyeq8kehehvjcv0va7nnnx9q9[0]}} & mqn5zl56qb4wkr4l5wjwjajufy9[47:15])
                                           | ({33{neomyeq8kehehvjcv0va7nnnx9q9[1]}} & mqn5zl56qb4wkr4l5wjwjajufy9[48:16])
                                           | ({33{neomyeq8kehehvjcv0va7nnnx9q9[2]}} & mqn5zl56qb4wkr4l5wjwjajufy9[63:31])
                                           | ({33{neomyeq8kehehvjcv0va7nnnx9q9[3]}} & mqn5zl56qb4wkr4l5wjwjajufy9[64:32])
                                           | ({33{neomyeq8kehehvjcv0va7nnnx9q9[4]}} & mqn5zl56qb4wkr4l5wjwjajufy9[32:0])
                                           ) : 
                                          of41hddih6s4bcn_3nwrp9[64:32];

  wire oyfgg_lfe45lc6el4jliokey58s   = rwsukdwq5hi04 & (dl7jvynj91yjq_ubriyt8rb5y1ksoen[32] & (~dl7jvynj91yjq_ubriyt8rb5y1ksoen[31]));
  wire e19bnjn_4s7whygso_r2koe_zzywlec = rwsukdwq5hi04 & (g4o3eqh6nb2enoez45n88_wji8vd4[32] & (~g4o3eqh6nb2enoez45n88_wji8vd4[31]));
  wire um41wkknnjh9udu8fdp06cdq = p49z763fixgor & (of41hddih6s4bcn_3nwrp9[64] & (~of41hddih6s4bcn_3nwrp9[63]));
  wire dih5lzug3zjlibji1cv3es26ul3 = o9baey2y_w0y & of41hddih6s4bcn_3nwrp9[66];

  wire kqz_c9hcgqb073u1cfs7na6a9jxz = (rwsukdwq5hi04 | mxwmmibxvjzkawbzq7wln ) & ((~dl7jvynj91yjq_ubriyt8rb5y1ksoen[32]) & dl7jvynj91yjq_ubriyt8rb5y1ksoen[31]); 
  wire g0jhd96dai4zuw94p6wnaoy90o9sh = (rwsukdwq5hi04 | mxwmmibxvjzkawbzq7wln ) & ((~g4o3eqh6nb2enoez45n88_wji8vd4[32]) & g4o3eqh6nb2enoez45n88_wji8vd4[31]); 
  wire mt2coznzoc3g0qkmqqvlk38ya = p49z763fixgor & ((~of41hddih6s4bcn_3nwrp9[64]) & of41hddih6s4bcn_3nwrp9[63]);
  wire j4e0_g8rg6u94qgpijpsj2pq = o9baey2y_w0y & ((~of41hddih6s4bcn_3nwrp9[66]) & (of41hddih6s4bcn_3nwrp9[65] | of41hddih6s4bcn_3nwrp9[64]));
  wire eiz1b4o4cqyrkrcm3fc =
                          oyfgg_lfe45lc6el4jliokey58s | kqz_c9hcgqb073u1cfs7na6a9jxz
                        | um41wkknnjh9udu8fdp06cdq | dih5lzug3zjlibji1cv3es26ul3
                        | mt2coznzoc3g0qkmqqvlk38ya | j4e0_g8rg6u94qgpijpsj2pq 
                        | q1xiho2m38dg2no_jw479l 
                        | ddu9petr88tlm28sdlv_a 
                        ;
  wire zi95lhlhuj1go8fk3qlnsc =
                          e19bnjn_4s7whygso_r2koe_zzywlec | g0jhd96dai4zuw94p6wnaoy90o9sh
                        | um41wkknnjh9udu8fdp06cdq   | dih5lzug3zjlibji1cv3es26ul3
                        | mt2coznzoc3g0qkmqqvlk38ya   | j4e0_g8rg6u94qgpijpsj2pq 
                        | zb7_0qoubehnq5_pbeisyo0v | c05m65au78yv406zviubh21ja
                        ;

  wire dt8rxjgth2bpc7ca = xgd98yfjs0wg1vjg;
  wire f49rkd3tra9rncu1ztlg = bn3hs_059enxzslhk7;

wire p8ccsbqbhzb9m1xhre = 
                        eiz1b4o4cqyrkrcm3fc 
                      | dt8rxjgth2bpc7ca
                      | zi95lhlhuj1go8fk3qlnsc 
                      | f49rkd3tra9rncu1ztlg
                      ;

  assign vjkz8n6i44pc7o = cwmxezrc3jv6hzxcfc & uig3ujuyq0_61kqb &
                             ( (hfssxn5khy43v3a  & ajb17ean3ect1us1)
                              |(myn68i_ltybiz        & royh8kfx4l6z206rgv) 
                              |(f2ky3p7ovwuqwa      & p8ccsbqbhzb9m1xhre))
                              ;

 wire [63:0] l4gwj3afpn4uqn7y0mj8e;
 assign  l4gwj3afpn4uqn7y0mj8e[31:0] = ( eiz1b4o4cqyrkrcm3fc ? 
                                        (
                                            ({32{oyfgg_lfe45lc6el4jliokey58s}} & 32'h80000000)
                                          | ({32{kqz_c9hcgqb073u1cfs7na6a9jxz | q1xiho2m38dg2no_jw479l }} & 32'h7fffffff)
                                          | ({32{ddu9petr88tlm28sdlv_a}} & 32'h7fff)
                                          | ({32{um41wkknnjh9udu8fdp06cdq | dih5lzug3zjlibji1cv3es26ul3}}& 32'h0)
                                          | ({32{mt2coznzoc3g0qkmqqvlk38ya | j4e0_g8rg6u94qgpijpsj2pq}} & 32'hffffffff)
                                        )
                                        : dl7jvynj91yjq_ubriyt8rb5y1ksoen[31:0]
                                      );

  assign  l4gwj3afpn4uqn7y0mj8e[63:32] = (zi95lhlhuj1go8fk3qlnsc ?
                                       (
                                           ({32{e19bnjn_4s7whygso_r2koe_zzywlec}} & 32'h80000000)
                                         | ({32{g0jhd96dai4zuw94p6wnaoy90o9sh | zb7_0qoubehnq5_pbeisyo0v }} & 32'h7fffffff)
                                         | ({32{c05m65au78yv406zviubh21ja}} & 32'h7fff)
                                         | ({32{um41wkknnjh9udu8fdp06cdq}} & 32'h80000000)
                                         | ({32{mt2coznzoc3g0qkmqqvlk38ya}} & 32'h7fffffff)
                                         | ({32{j4e0_g8rg6u94qgpijpsj2pq}} & 32'hffffffff)
                                         | ({32{dih5lzug3zjlibji1cv3es26ul3}} & 32'h0)
                                       )
                                       : lbvwt_z2shtjwj ? {32{nb3w1rq_ny95rvrt[31]}} : g4o3eqh6nb2enoez45n88_wji8vd4[31:0]
                                      );
  assign  nb3w1rq_ny95rvrt[31:0] =
                                        ({32{hfssxn5khy43v3a}} & r8yaegh9ba96e1xa[31:0]) 
                                      | ({32{myn68i_ltybiz      }} & cmdsrflujxwd007q[31:0]) 
                                      | ({32{f2ky3p7ovwuqwa    }} & l4gwj3afpn4uqn7y0mj8e[31:0]) 
                                      ;

  assign  nb3w1rq_ny95rvrt[63:32] =
                                        ({32{hfssxn5khy43v3a}} & r8yaegh9ba96e1xa[63:32]) 
                                      | ({32{myn68i_ltybiz      }} & cmdsrflujxwd007q[63:32]) 
                                      | ({32{f2ky3p7ovwuqwa    }} & l4gwj3afpn4uqn7y0mj8e[63:32]) 
                                      ;

  assign p_yx415so7q1vohijb = qbpmsk2;


endmodule
        










































































module i6tr_dyutx06rp9skham4 # (
  parameter ctu6y0yy1_ = 5   
) (
  
  
  
  input  [64-1:0] amgi_rqhtd007,       
  input  [64-1:0] h33_crpt0l75o,    
  input  [64-1:0] g7tawq8tp6,
  input  [64-1:0] jmf1rwo8,
  input  [64-1:0] xo5bwsw4j8a,        
  input  [105-1:0] xlkm1ikvsatc2,

  
  
  
  
  output lzal8kswefl9gv4kqdclkfx23, 
  output [64-1:0] udhgtu0ck3hr1aj,
  output [5:0] so4zxlxtb1t9lx,
  input  [64-1:0] q7c4bjf1j8kujxtvei,

  
  
  
  
  output bdd_smghkpbtvkxlxpdyq2perm, 
  output [64-1:0] sznwd73uhzrymh69lt9dcfpa,
  output [ctu6y0yy1_-1:0] l4ik_e9aa1bhu66b138,
  input  [64-1:0] zvnjpa2uy_h98fk1u8zei9w,

  
  
  
  
  output sazh4of6fhumdu0qyo1yjk2u00eee, 
  output [64-1:0] m9e0b_s90djin0iqc0ts9v,
  output [64-1:0] yqf19lhru49yxe2r5x0diu,
  input  [64-1:0] yhru2nhdb63arfxbb25pgcp,

  
  
  
  output [64-1:0] nb3w1rq_ny95rvrt,
    
  output vjkz8n6i44pc7o,
    
  input  m6ouh9hkcy63fxj02, 

  
  
  input  gf33atgy,
  input  ru_wi 

  );

localparam yk7 = 2;
localparam m0qq = 4;
localparam dk34z = 8;









wire vuz9jubu4     = xlkm1ikvsatc2[11:11];
wire i2ouxsq7e     = xlkm1ikvsatc2[12:12];
wire gxr7nn3    = xlkm1ikvsatc2[13:13];
wire mx3rzhyu8f34    = xlkm1ikvsatc2[14:14];
wire xb6zb0of    = xlkm1ikvsatc2[15:15];
wire ou2t9osgil39    = xlkm1ikvsatc2[16:16];

wire [5:0] v4an2pt_ara = xlkm1ikvsatc2[10:5];





wire [4:0] smo9yw4mrr0p_;
wire [31:0] b1k_vgv9hjhr7h2;

assign smo9yw4mrr0p_[2:0] = v4an2pt_ara[2:0];
assign smo9yw4mrr0p_[4:3] = {
                         ({2{(vuz9jubu4 | i2ouxsq7e)}} & {2'b0}) |
                         ({2{(gxr7nn3 | mx3rzhyu8f34)}} & {1'b0,v4an2pt_ara[3]}) |
                         ({2{(xb6zb0of | ou2t9osgil39)}} & {v4an2pt_ara[4:3]})
						};


genvar i;
generate 
	for(i=0; i<32; i=i+1) begin: r0pwqlpmco
		assign b1k_vgv9hjhr7h2[i] = (smo9yw4mrr0p_==i[4:0]);    
	end
endgenerate


wire [31:0] abm09env4nq25q4yk;


wire [31:0] nrznb44cczc12ko9;

generate 
	for(i=0; i<32; i=i+1) begin: aon0u5bpt_tjqf
		assign nrznb44cczc12ko9[i] = |b1k_vgv9hjhr7h2[i:0];
	end
endgenerate

assign abm09env4nq25q4yk = ~nrznb44cczc12ko9;

wire [64-1:0] dowh377m4y1o = amgi_rqhtd007;












wire [dk34z-1:0] dcwpqmycx30;
wire [dk34z-1:0] q0sbhwkxjdq56;






wire [m0qq-1:0]  k6bpq_fej6maw;
wire [m0qq-1:0]  f8libiup_8xtk;



wire [31:0]    db_w4igipz8oag = abm09env4nq25q4yk;
wire [31:0]    f7ywgzs25mvcjk1do = nrznb44cczc12ko9;
wire [15:0]    sp_mih3885s0so0_3 = abm09env4nq25q4yk[15:0];
wire [15:0]    af5vksf5srbn1 = nrznb44cczc12ko9[15:0];
wire [ 7:0]    cujm807_npq0dq2k  = abm09env4nq25q4yk[7:0];
wire [ 7:0]    mnjb617natbpvf  = nrznb44cczc12ko9[7:0];
wire [yk7-1:0]  a1w3tnd5vr3n;
wire [yk7-1:0]  axkj4dvy_e_cde_z;

gr40tady98ryto733e #(
    .yk7(yk7),
    .m0qq(m0qq),
    .dk34z(dk34z)
)  q0jzdszo0hdxo9q0sobo (
	.c5qrwj5sm0vc      ( dowh377m4y1o      ),     
	.of4kpekzgop8    ( 64'b0 ),     
	.l59fhx3o23g9ig ( 64'b0 ),     
	.p2v9igi9t66348 ( 64'b0 ),     
	.utwav9is_83yd6ng0 ( db_w4igipz8oag  ),     
	.sdmfqus_d4n5v3k ( f7ywgzs25mvcjk1do  ),     
	.ghpvhjxwavld6r6r0w2 ( sp_mih3885s0so0_3  ),     
	.berx62p9_hc2bfcnyn0 ( af5vksf5srbn1  ),     
	.ky3ucnc3e8n4c_iz  ( cujm807_npq0dq2k   ),     
	.v98eqhdqs8d1wk_qf2  ( mnjb617natbpvf   ),     
	.p2tb25qpyet2a_c    (               ),     
	.wms1mxki5gyfyc    (               ),     
	.tkuhwm5tyjr    ( a1w3tnd5vr3n   ),     
	.rg1trb_7w92    ( axkj4dvy_e_cde_z   ),     
	.a1bp0x22t5vu4q    ( k6bpq_fej6maw   ),     
	.rgxbhxlvt61yfzn    ( f8libiup_8xtk   ),     
	.jpltrmmj8jw4lh_  (               ),     
	.gs2s9lvzd_phhnv  (               ),     
	.j694o6frj_680_g     ( dcwpqmycx30    ),     
	.n2nedhasxux7buh     ( q0sbhwkxjdq56    ),     
	.fnv_7okzmo6y4ne85   (               ),     
	.u_frczxmkmo88ujnp   (               )      
);


wire [yk7-1:0] vkezs43ppvgfxm;
wire [m0qq-1:0] l7sxt6i5wgf0;
wire [dk34z-1:0] ptzoc7dl32t9u7;

generate 
	for(i=0; i<yk7; i=i+1) begin: v25k3tdkvl6rnd56c
        assign vkezs43ppvgfxm[i] = dowh377m4y1o[i*32+31];
	end
endgenerate

generate 
	for(i=0; i<m0qq; i=i+1) begin: yapihobpzjdh3
        assign l7sxt6i5wgf0[i] = dowh377m4y1o[i*16+15];
	end
endgenerate

generate 
	for(i=0; i<dk34z; i=i+1) begin: qfiu1hh7vlgjrd
        assign ptzoc7dl32t9u7[i] = dowh377m4y1o[i*8+7];
	end
endgenerate

wire [yk7-1:0] sxoos4_vgs3kfcq;
wire [yk7-1:0] ciqq1yyzkp_9a5ssv;
wire [yk7-1:0] sonxjnnyfadhdpt6qqzilre;
wire [yk7-1:0] r8ftllfi_osy0q4wv213;
wire [31:0]   epp_b2cftx920o50zt[yk7-1:0];
wire [m0qq-1:0] u5va18k93w84464;
wire [m0qq-1:0] fetsdr04nryh85t;
wire [m0qq-1:0] bzvao_bivg2r9edn5d;
wire [m0qq-1:0] mjqmdpme83lhf1369;
wire [15:0]   o4wf4fb79_qnhywmbapm[m0qq-1:0];
wire [dk34z-1:0] zl3qk4gsg2ttv1m;
wire [dk34z-1:0] szkb51g7fmynxa;
wire [dk34z-1:0] vsc2c4dt3pu3_h2lmlgl;
wire [dk34z-1:0] jixyajtkls74wq_ivfl;
wire [7:0] fioltoxti5m3lhgyr04vq[dk34z-1:0];

generate 
	for(i=0; i<yk7; i=i+1) begin: qe8iuuxvwmc74rvhluin
        assign sxoos4_vgs3kfcq[i]           = (ou2t9osgil39 & ~vkezs43ppvgfxm[i] & ~a1w3tnd5vr3n[i]) | 
                                              (xb6zb0of & ~vkezs43ppvgfxm[i] & ~a1w3tnd5vr3n[i]) |
                                              (xb6zb0of &  vkezs43ppvgfxm[i] & ~axkj4dvy_e_cde_z[i]);
        
        assign ciqq1yyzkp_9a5ssv[i]           = (ou2t9osgil39 & ~vkezs43ppvgfxm[i] &  a1w3tnd5vr3n[i]) |
                                              (xb6zb0of & ~vkezs43ppvgfxm[i] &  a1w3tnd5vr3n[i]); 
        
        assign sonxjnnyfadhdpt6qqzilre[i]        = (xb6zb0of &  vkezs43ppvgfxm[i] &  axkj4dvy_e_cde_z[i]);
        
        assign r8ftllfi_osy0q4wv213[i]          = (ou2t9osgil39 &  vkezs43ppvgfxm[i]);
        
        assign epp_b2cftx920o50zt[i]        = sxoos4_vgs3kfcq[i]    ? dowh377m4y1o[i*32+31:i*32] :
                                              ciqq1yyzkp_9a5ssv[i]    ? abm09env4nq25q4yk :
                                              sonxjnnyfadhdpt6qqzilre[i] ? nrznb44cczc12ko9 : 32'b0;
	end
endgenerate

wire [15:0] nbrsrkf6kgv1s5i[m0qq-1:0];

generate 
	for(i=0; i<m0qq; i=i+1) begin: kips6mgae59lg_p40o
		assign nbrsrkf6kgv1s5i[i]     = dowh377m4y1o[i*16+15:i*16];

		assign u5va18k93w84464[i]  = (mx3rzhyu8f34 & ~l7sxt6i5wgf0[i] & ~k6bpq_fej6maw[i]) | 
		                             (gxr7nn3 & ~l7sxt6i5wgf0[i] & ~k6bpq_fej6maw[i]) |
		                             (gxr7nn3 & l7sxt6i5wgf0[i]  & ~f8libiup_8xtk[i]);
 
		assign fetsdr04nryh85t[i]  = (mx3rzhyu8f34 & ~l7sxt6i5wgf0[i] & k6bpq_fej6maw[i]) |
		                             (gxr7nn3 & ~l7sxt6i5wgf0[i] & k6bpq_fej6maw[i]); 

		assign bzvao_bivg2r9edn5d[i]= (gxr7nn3 & l7sxt6i5wgf0[i] & f8libiup_8xtk[i]);

		assign mjqmdpme83lhf1369[i]  = (mx3rzhyu8f34 & l7sxt6i5wgf0[i]);

		assign o4wf4fb79_qnhywmbapm[i]= u5va18k93w84464[i] ? nbrsrkf6kgv1s5i[i] :
		                              fetsdr04nryh85t[i] ? abm09env4nq25q4yk[15:0] :
		                              bzvao_bivg2r9edn5d[i] ? nrznb44cczc12ko9[15:0] : 16'h0;
	end

endgenerate

wire [7:0] vi50mb99o93uu[dk34z-1:0];
assign vi50mb99o93uu[0] = dowh377m4y1o[7:0];
assign vi50mb99o93uu[1] = dowh377m4y1o[15:8];
assign vi50mb99o93uu[2] = dowh377m4y1o[23:16];
assign vi50mb99o93uu[3] = dowh377m4y1o[31:24];

generate 
	for(i=0; i<dk34z; i=i+1) begin: v6mu_d6dvwqjjmx43z
		assign vi50mb99o93uu[i]      = dowh377m4y1o[i*8+7:i*8];
		assign zl3qk4gsg2ttv1m[i]   = (i2ouxsq7e & ~ptzoc7dl32t9u7[i] & ~dcwpqmycx30[i]) | 
		                             (vuz9jubu4 & ~ptzoc7dl32t9u7[i] & ~dcwpqmycx30[i]) |
		                             (vuz9jubu4 & ptzoc7dl32t9u7[i]  & ~q0sbhwkxjdq56[i]);
 
		assign szkb51g7fmynxa[i]   = (i2ouxsq7e & ~ptzoc7dl32t9u7[i] & dcwpqmycx30[i]) |
		                             (vuz9jubu4 & ~ptzoc7dl32t9u7[i] & dcwpqmycx30[i]); 

		assign vsc2c4dt3pu3_h2lmlgl[i]= (vuz9jubu4 & ptzoc7dl32t9u7[i] & q0sbhwkxjdq56[i]);

		assign jixyajtkls74wq_ivfl[i]  = (i2ouxsq7e & ptzoc7dl32t9u7[i]);

		assign fioltoxti5m3lhgyr04vq[i]= zl3qk4gsg2ttv1m[i] ? vi50mb99o93uu[i] :
		                             szkb51g7fmynxa[i] ? abm09env4nq25q4yk[7:0] :
		                             vsc2c4dt3pu3_h2lmlgl[i] ? nrznb44cczc12ko9[7:0] : 8'h0;
	end

endgenerate

wire b8pejgc4p = (ou2t9osgil39 | xb6zb0of);
wire q0pof4ypop = (mx3rzhyu8f34 | gxr7nn3);
wire lyzbi5  = (i2ouxsq7e  | vuz9jubu4 );

wire [64-1:0] huf4d5e5ey8_pj9r6_;
assign huf4d5e5ey8_pj9r6_ = b8pejgc4p ? {epp_b2cftx920o50zt[1],epp_b2cftx920o50zt[0]}:
                          q0pof4ypop ? {o4wf4fb79_qnhywmbapm[3],o4wf4fb79_qnhywmbapm[2],o4wf4fb79_qnhywmbapm[1],o4wf4fb79_qnhywmbapm[0]} :
                          {fioltoxti5m3lhgyr04vq[7],fioltoxti5m3lhgyr04vq[6],fioltoxti5m3lhgyr04vq[5],fioltoxti5m3lhgyr04vq[4],fioltoxti5m3lhgyr04vq[3],fioltoxti5m3lhgyr04vq[2],fioltoxti5m3lhgyr04vq[1],fioltoxti5m3lhgyr04vq[0]};

wire lkoe_jcrsl9h3;
assign lkoe_jcrsl9h3    = b8pejgc4p ? ~(&sxoos4_vgs3kfcq) :
                          q0pof4ypop ? ~(&u5va18k93w84464) :
						  lyzbi5  ? ~(&zl3qk4gsg2ttv1m)  :
						  1'b0;

wire zby8wjkievope63 = vuz9jubu4 | i2ouxsq7e | gxr7nn3 | mx3rzhyu8f34 | xb6zb0of | ou2t9osgil39;














wire vgwjh46b2 = xlkm1ikvsatc2[17:17];
wire niqd13o6pl6 = xlkm1ikvsatc2[18:18];
wire bmunld04drsu = xlkm1ikvsatc2[19:19];
wire eprzju601h4a = xlkm1ikvsatc2[20:20];
wire hs24zc9dxe8i = xlkm1ikvsatc2[21:21];
wire okgyx6mwq_36 = xlkm1ikvsatc2[22:22];
wire r89bv6_v_ = xlkm1ikvsatc2[23:23];
wire vh4cec1h_x4g = xlkm1ikvsatc2[24:24];
wire ghj6n9znmzg = xlkm1ikvsatc2[25:25];
wire e3_b_jyl7dz5 = xlkm1ikvsatc2[26:26];


wire [15:0] w3i7fmc5_fpu = {{8{amgi_rqhtd007[7]}}, amgi_rqhtd007[7:0]};
wire [15:0] bwr0xd58 = {{8{amgi_rqhtd007[15]}}, amgi_rqhtd007[15:8]};
wire [15:0] tq1r41ocd = {{8{amgi_rqhtd007[23]}}, amgi_rqhtd007[23:16]};
wire [15:0] aod8pj9v9 = {{8{amgi_rqhtd007[31]}}, amgi_rqhtd007[31:24]};
wire [15:0] gwt775m0yeh = {{8{amgi_rqhtd007[39]}}, amgi_rqhtd007[39:32]};
wire [15:0] yjuatb12wo_v0 = {{8{amgi_rqhtd007[47]}}, amgi_rqhtd007[47:40]};
wire [15:0] caqo7gtetxj9pg = {{8{amgi_rqhtd007[55]}}, amgi_rqhtd007[55:48]};
wire [15:0] vjnxnk3kju = {{8{amgi_rqhtd007[63]}}, amgi_rqhtd007[63:56]};


wire [15:0] r0qh3j03 = {8'h0, amgi_rqhtd007[7:0]};
wire [15:0] ghebcpe_ikm = {8'h0, amgi_rqhtd007[15:8]};
wire [15:0] e0avt8ih2o = {8'h0, amgi_rqhtd007[23:16]};
wire [15:0] dtcb6qvfx0mqm = {8'h0, amgi_rqhtd007[31:24]};
wire [15:0] j5bs8a69iapw = {{8{1'b0}}, amgi_rqhtd007[39:32]};
wire [15:0] f5rca544us9 = {{8{1'b0}}, amgi_rqhtd007[47:40]};
wire [15:0] aw397dqrask_vf = {{8{1'b0}}, amgi_rqhtd007[55:48]};
wire [15:0] cn9kzckwrh224h = {{8{1'b0}}, amgi_rqhtd007[63:56]};

wire [64-1:0] p7e55yl2xz_s76csdl;
assign p7e55yl2xz_s76csdl = ({64{vgwjh46b2}} & {yjuatb12wo_v0,gwt775m0yeh,bwr0xd58,w3i7fmc5_fpu}) |
                            ({64{niqd13o6pl6}} & {caqo7gtetxj9pg,gwt775m0yeh,tq1r41ocd,w3i7fmc5_fpu}) |
                            ({64{bmunld04drsu}} & {vjnxnk3kju,gwt775m0yeh,aod8pj9v9,w3i7fmc5_fpu}) |
                            ({64{eprzju601h4a}} & {vjnxnk3kju,yjuatb12wo_v0,aod8pj9v9,bwr0xd58}) |
                            ({64{hs24zc9dxe8i}} & {vjnxnk3kju,caqo7gtetxj9pg,aod8pj9v9,tq1r41ocd}) |
                            ({64{okgyx6mwq_36}} & {f5rca544us9,j5bs8a69iapw,ghebcpe_ikm,r0qh3j03}) |
                            ({64{r89bv6_v_}} & {aw397dqrask_vf,j5bs8a69iapw,e0avt8ih2o,r0qh3j03}) |
                            ({64{vh4cec1h_x4g}} & {cn9kzckwrh224h,j5bs8a69iapw,dtcb6qvfx0mqm,r0qh3j03}) |
                            ({64{ghj6n9znmzg}} & {cn9kzckwrh224h,f5rca544us9,dtcb6qvfx0mqm,ghebcpe_ikm}) |
                            ({64{e3_b_jyl7dz5}} & {cn9kzckwrh224h,aw397dqrask_vf,dtcb6qvfx0mqm,e0avt8ih2o}) ;

wire cg_xvkpcb5oe4ov3r = 
                          vgwjh46b2 |
                          niqd13o6pl6 |
                          bmunld04drsu |
                          eprzju601h4a |
                          hs24zc9dxe8i |
                          okgyx6mwq_36 |
                          r89bv6_v_ |
                          vh4cec1h_x4g |
                          ghj6n9znmzg |
                          e3_b_jyl7dz5;












wire i_9e3rjoddz0u = xlkm1ikvsatc2[27:27];
wire zf6n5ojitnzc = xlkm1ikvsatc2[28:28];
wire l80mr2fy = xlkm1ikvsatc2[29:29];
wire d5cfr3w4s7he9 = xlkm1ikvsatc2[30:30];
wire ei02jqe0nb = xlkm1ikvsatc2[56:56];
wire fjl7lngye = xlkm1ikvsatc2[57:57];
wire vfqtv67tls8p = xlkm1ikvsatc2[58:58];
wire rfu_9o52ml0w = xlkm1ikvsatc2[59:59];

wire [64-1:0] qyh4fb808wpe28g8;
assign qyh4fb808wpe28g8 = ({64{i_9e3rjoddz0u}} & {amgi_rqhtd007[47:32],g7tawq8tp6[47:32],amgi_rqhtd007[15: 0],g7tawq8tp6[15: 0]}) |
                          ({64{zf6n5ojitnzc}} & {amgi_rqhtd007[47:32],g7tawq8tp6[63:48],amgi_rqhtd007[15: 0],g7tawq8tp6[31:16]}) |
                          ({64{l80mr2fy}} & {amgi_rqhtd007[63:48],g7tawq8tp6[47:32],amgi_rqhtd007[31:16],g7tawq8tp6[15: 0]}) |
                          ({64{d5cfr3w4s7he9}} & {amgi_rqhtd007[63:48],g7tawq8tp6[63:48],amgi_rqhtd007[31:16],g7tawq8tp6[31:16]}) |
                          ({64{ei02jqe0nb}} & {amgi_rqhtd007[31: 0],g7tawq8tp6[31: 0]}) |
                          ({64{fjl7lngye}} & {amgi_rqhtd007[31: 0],g7tawq8tp6[63:32]}) |
                          ({64{vfqtv67tls8p}} & {amgi_rqhtd007[63:32],g7tawq8tp6[31: 0]}) |
                          ({64{rfu_9o52ml0w}} & {amgi_rqhtd007[63:32],g7tawq8tp6[63:32]});

wire ccm19fkdl1_0ex2 = 
                        i_9e3rjoddz0u |
                        zf6n5ojitnzc |
                        l80mr2fy |
                        d5cfr3w4s7he9 |
                        ei02jqe0nb |
                        fjl7lngye |
                        vfqtv67tls8p |
                        rfu_9o52ml0w;













wire vmirs3c3sk  = xlkm1ikvsatc2[39:39];
wire qosva   = xlkm1ikvsatc2[40:40];
wire r61tzvs   = xlkm1ikvsatc2[41:41];
wire wseodi = xlkm1ikvsatc2[42:42];
wire q7sm7ubc  = xlkm1ikvsatc2[43:43];
wire n5vmjq_  = xlkm1ikvsatc2[44:44];
wire m9d8wlbj = xlkm1ikvsatc2[45:45];
wire s5_j28hb4  = xlkm1ikvsatc2[46:46];
wire uqnc92  = xlkm1ikvsatc2[47:47];

wire cnuj = vmirs3c3sk | qosva | r61tzvs;
wire am6ee = wseodi | q7sm7ubc | n5vmjq_;
wire wcxui5h = m9d8wlbj | s5_j28hb4 | uqnc92;
wire zra9dfflxqu = vmirs3c3sk | wseodi;
wire y11_ = zra9dfflxqu | m9d8wlbj;

wire [31:0] iocihvyxfkea[yk7-1:0];
wire [31:0] f83otta4ue5fult[yk7-1:0];
wire [31:0] fi9c7sy7[yk7-1:0];
wire [31:0] bn0xke0e2[yk7-1:0];
wire [32:0] fbox7ssd7[yk7-1:0];
wire [31:0] bv9nyvtl6ox[yk7-1:0];
wire [yk7-1:0]         ebs5_h3sb5sl;
wire [5:0]            aeh7ngbsvis5xa[yk7-1:0];



generate 
	for(i=0; i<yk7; i=i+1) begin: dlf0j049jp3yhgv_9rq2iqs
        assign iocihvyxfkea[i]  =({32{wcxui5h}} & amgi_rqhtd007[i*32+31:i*32]);
        
        assign f83otta4ue5fult[i] = y11_ ? {iocihvyxfkea[i][30:0], ~iocihvyxfkea[i][31]} : iocihvyxfkea[i];
        assign ebs5_h3sb5sl[i]  = s5_j28hb4 ? 1'b0 : m9d8wlbj ? amgi_rqhtd007[i*32+31] : 1'b1;
        assign fbox7ssd7[i]       = {bn0xke0e2[i],1'b1};
	end

endgenerate

genvar j;

generate 
	for(j=0; j<yk7; j=j+1) begin: f07r9wn6_fqqnndhcfpo
	    for(i=0; i<32; i=i+1) begin: vmxcdfimeka1eljtc0
	    	assign fi9c7sy7[j][i] = ebs5_h3sb5sl[j] ^ f83otta4ue5fult[j][i];
	    	assign bn0xke0e2[j][i] = |fi9c7sy7[j][31:i];
	    	assign bv9nyvtl6ox[j][i] = ~fbox7ssd7[j][i+1] & fbox7ssd7[j][i];
	    end
	end
endgenerate


generate 
	for(i=0; i<yk7; i=i+1) begin: x3_eqgu489sw7m0lrl8d15y

qlm10lcv_tyz847h7k qah8ibwsvidu_t6jawju
(
	.wz0wek1lz0  ( bv9nyvtl6ox[i]  ),
	.i8vml4gn     ( aeh7ngbsvis5xa[i] ) 
);

	end

endgenerate


wire [16:0] z30vfsxam[m0qq-1:0];
wire [15:0] kk2p2ihzu4l5zpc2iv2[m0qq-1:0];
wire [15:0] g_csjzq02dcf7ty65stph[m0qq-1:0];
wire [15:0] emereeit[m0qq-1:0];
wire [15:0] ocq7bbomyap[m0qq-1:0];
wire [15:0] h3bjjr6eh0hvyii[m0qq-1:0];
wire [m0qq-1:0] hgmb3wx5bucb;
wire [4:0] vc3jrp5f4guyd3[m0qq-1:0];

generate 
	for(i=0; i<m0qq; i=i+1) begin: xf9e9l8qah0i9amook1sns
        assign kk2p2ihzu4l5zpc2iv2[i] = ({16{am6ee}} & amgi_rqhtd007[i*16+15:i*16]);
        
        assign g_csjzq02dcf7ty65stph[i] = wseodi ? {kk2p2ihzu4l5zpc2iv2[i][14:0], ~kk2p2ihzu4l5zpc2iv2[i][15]} : kk2p2ihzu4l5zpc2iv2[i];
        
        assign hgmb3wx5bucb[i] = q7sm7ubc ? 1'b0 : wseodi ? amgi_rqhtd007[i*16+15] : 1'b1;
        assign z30vfsxam[i] = {emereeit[i],1'b1};
	end

endgenerate

generate 
	for(j=0; j<m0qq; j=j+1) begin: fcy26p_kz2gscqx8j1no7
	    for(i=0; i<16; i=i+1) begin: g5myv2ya67ic5ujsqzhpq
	    	assign ocq7bbomyap[j][i] = hgmb3wx5bucb[j] ^ g_csjzq02dcf7ty65stph[j][i];
	    	assign emereeit[j][i] = |ocq7bbomyap[j][15:i];
	    	assign h3bjjr6eh0hvyii[j][i] = ~z30vfsxam[j][i+1] & z30vfsxam[j][i];
	    end
	end
endgenerate

generate 
	for(i=0; i<m0qq; i=i+1) begin: nb8rnqriutgxdrpfud9g

h09sftk403rm5tnmsmed j87vwe6v9ixiztmi087
(
	.wz0wek1lz0  ( h3bjjr6eh0hvyii[i]  ),
	.i8vml4gn     ( vc3jrp5f4guyd3[i] ) 
);

	end

endgenerate


wire [8:0] ypxxakedfe2wh[dk34z-1:0];
wire [7:0] dhg7cetpwwek6iy[dk34z-1:0];
wire [7:0] xjlaag0hyk7_adr9nw[dk34z-1:0];
wire [7:0] wr4f86a4wwry[dk34z-1:0];
wire [7:0] pfo4ugw6u9evh[dk34z-1:0];
wire [7:0] wqcuzfrqkdn6b2r34[dk34z-1:0];
wire [dk34z-1:0] irjvmserpbwmy6xgwuad;
wire [3:0] lpsqexg2b4gjrah_cib[dk34z-1:0];

generate 
	for(i=0; i<dk34z; i=i+1) begin: ymv48nz0nz1twi1phpgw
        assign dhg7cetpwwek6iy[i] = amgi_rqhtd007[i*8+7:i*8];
        assign xjlaag0hyk7_adr9nw[i] = vmirs3c3sk ? {dhg7cetpwwek6iy[i][6:0], ~dhg7cetpwwek6iy[i][7]} : dhg7cetpwwek6iy[i];
        
        assign irjvmserpbwmy6xgwuad[i] = qosva ? 1'b0 : vmirs3c3sk ? amgi_rqhtd007[i*8+7] : 1'b1;
        assign ypxxakedfe2wh[i] = {wr4f86a4wwry[i],1'b1};
	end
endgenerate

generate 
	for(j=0; j<dk34z; j=j+1) begin: w_072rw5emfatxpa883
	    for(i=0; i<8; i=i+1) begin: w_072rw5emfatxpa883
	    	assign pfo4ugw6u9evh[j][i] = irjvmserpbwmy6xgwuad[j] ^ xjlaag0hyk7_adr9nw[j][i];
	    	assign wr4f86a4wwry[j][i] = |pfo4ugw6u9evh[j][7:i];
	    	assign wqcuzfrqkdn6b2r34[j][i] = ~ypxxakedfe2wh[j][i+1] & ypxxakedfe2wh[j][i];
	    end
	end
endgenerate


generate 
	for(i=0; i<dk34z; i=i+1) begin: vms19i7p4uzsvybfij
sqkb0d8aic395m2pbugz ch1umbyoxoc9w4z1d2vtv
(
	.wz0wek1lz0  ( wqcuzfrqkdn6b2r34[i]  ),
	.i8vml4gn     ( lpsqexg2b4gjrah_cib[i] ) 
);
	end
endgenerate

wire [64-1:0] xx_4lcsv8bjm23ylo;
assign xx_4lcsv8bjm23ylo = cnuj ?  {4'b0, lpsqexg2b4gjrah_cib[7],4'b0, lpsqexg2b4gjrah_cib[6],4'b0, lpsqexg2b4gjrah_cib[5],4'b0, lpsqexg2b4gjrah_cib[4],4'b0, lpsqexg2b4gjrah_cib[3],4'b0, lpsqexg2b4gjrah_cib[2],4'b0, lpsqexg2b4gjrah_cib[1],4'b0, lpsqexg2b4gjrah_cib[0]} :
                        am6ee ? {11'b0, vc3jrp5f4guyd3[3], 11'b0, vc3jrp5f4guyd3[2],11'b0, vc3jrp5f4guyd3[1], 11'b0, vc3jrp5f4guyd3[0]} :
                        {26'b0,aeh7ngbsvis5xa[1],26'b0,aeh7ngbsvis5xa[0]};

wire uq3eiceihlgu = 
                      vmirs3c3sk  | 
                      qosva   | 
                      r61tzvs   | 
                      wseodi | 
                      q7sm7ubc  | 
                      n5vmjq_  | 
                      m9d8wlbj | 
                      s5_j28hb4  | 
                      uqnc92  ;















wire vfjyij  = xlkm1ikvsatc2[48:48];
wire us171m8a = xlkm1ikvsatc2[49:49];
wire [5:0] s119d6od = xlkm1ikvsatc2[10:5]; 
wire [ctu6y0yy1_-1:0] tv5o2dgsibw = g7tawq8tp6[ctu6y0yy1_-1:0];

wire [ctu6y0yy1_-1:0] eni83nk = ({ctu6y0yy1_{vfjyij}}  & tv5o2dgsibw[ctu6y0yy1_-1:0]) |
                          ({ctu6y0yy1_{us171m8a}} & s119d6od[ctu6y0yy1_-1:0]);





wire [64-1:0] item2h0zpygqk9zeo;
i6_4g5fspqlv1svn #(64) wlvhd378om0a9(amgi_rqhtd007, item2h0zpygqk9zeo);



wire pfj780v6il2rtp;
assign lzal8kswefl9gv4kqdclkfx23 = pfj780v6il2rtp;
assign udhgtu0ck3hr1aj = item2h0zpygqk9zeo;
assign so4zxlxtb1t9lx = ~eni83nk;

wire [64-1:0] k69l77w397qhwjeh;

assign k69l77w397qhwjeh = q7c4bjf1j8kujxtvei;
assign pfj780v6il2rtp = us171m8a | vfjyij;











wire onyfmj  = xlkm1ikvsatc2[50:50];
wire t7ia9se062 = xlkm1ikvsatc2[51:51];
wire [5:0] sy6s77blv256 = xlkm1ikvsatc2[10:5];
wire [4:0] o8jezj1t9w85e = sy6s77blv256[4:0];
wire gkjybnhfjsie3o;

wire [4:0] k_n_y9t30mvy4j5 = ({5{onyfmj}} & g7tawq8tp6[4:0]) |
                            ({5{t7ia9se062}} & o8jezj1t9w85e[4:0]);


assign bdd_smghkpbtvkxlxpdyq2perm = gkjybnhfjsie3o;
assign sznwd73uhzrymh69lt9dcfpa       = amgi_rqhtd007;
assign l4ik_e9aa1bhu66b138       = {1'b0,k_n_y9t30mvy4j5};
assign sazh4of6fhumdu0qyo1yjk2u00eee = 1'b0;
assign m9e0b_s90djin0iqc0ts9v = 64'b0;   
assign yqf19lhru49yxe2r5x0diu = 64'b0;

wire [64-1:0] slmojwuw5628djvr;

assign slmojwuw5628djvr = {{32{zvnjpa2uy_h98fk1u8zei9w[31]}},zvnjpa2uy_h98fk1u8zei9w[31:0]};
assign gkjybnhfjsie3o = onyfmj | t7ia9se062;





wire mezhady2w = xlkm1ikvsatc2 [52:52];

wire [64-1:0] n8v1vqp24ko3fof;
assign n8v1vqp24ko3fof = (jmf1rwo8 & amgi_rqhtd007) | (~jmf1rwo8 & g7tawq8tp6);

wire dzs4lvfhrbn6q = mezhady2w;





wire e_vv = xlkm1ikvsatc2[53:53];
wire [5:0] iy6znwx03 = xlkm1ikvsatc2 [10:5];
wire a1fqfh04bor = (iy6znwx03[2:0] == 3'b000) & e_vv; 
wire mpovguulfu = (iy6znwx03[2:0] == 3'b001) & e_vv;
wire xzujh5p5lh2qk3 = (iy6znwx03[2:0] == 3'b010) & e_vv;
wire l6jbfhfho5 = (iy6znwx03[2:0] == 3'b011) & e_vv;
wire aio46bn_krne = (iy6znwx03[2:0] == 3'b100) & e_vv; 
wire dn819og59mg7 = (iy6znwx03[2:0] == 3'b101) & e_vv;
wire cuz3l4ac7ygj = (iy6znwx03[2:0] == 3'b110) & e_vv;
wire jytc3ic8pgzqg4_ = (iy6znwx03[2:0] == 3'b111) & e_vv;
wire [64-1:0] tkuokqnj0qhz = {{8{jytc3ic8pgzqg4_}}, {8{cuz3l4ac7ygj}}, {8{dn819og59mg7}}, {8{aio46bn_krne}},{8{l6jbfhfho5}}, {8{xzujh5p5lh2qk3}}, {8{mpovguulfu}}, {8{a1fqfh04bor}}};
wire [64-1:0] fja3sq8t73lm0x = {8{amgi_rqhtd007[7:0]}};

wire [64-1:0] lfkclmsw9nw8cco_8c;
assign lfkclmsw9nw8cco_8c = (tkuokqnj0qhz & fja3sq8t73lm0x) | (~tkuokqnj0qhz & xo5bwsw4j8a);
wire ut1dkcj1azkbznfp = e_vv;






wire soa15g4rw8  = xlkm1ikvsatc2[54:54];
wire r3zfud = xlkm1ikvsatc2[55:55];

wire [64-1:0] q96ft3lmyjaeecp_2x45p;
assign q96ft3lmyjaeecp_2x45p = ({64{soa15g4rw8}} & {amgi_rqhtd007[55:48],amgi_rqhtd007[63:56],amgi_rqhtd007[39:32],amgi_rqhtd007[47:40],amgi_rqhtd007[23:16],amgi_rqhtd007[31:24],amgi_rqhtd007[7:0],amgi_rqhtd007[15:8]}) |
                          ({64{r3zfud}} & {amgi_rqhtd007[47:32],amgi_rqhtd007[63:48],amgi_rqhtd007[15:0],amgi_rqhtd007[31:16]});

wire z0v1bqkq5qn284wu = soa15g4rw8 | r3zfud;








wire pldtey61 = xlkm1ikvsatc2[31];
wire vribxr_dbn = xlkm1ikvsatc2[32];
wire l5bnwm = xlkm1ikvsatc2[33];
wire lgnvbn = xlkm1ikvsatc2[34];
wire ksxzc99stv9 = xlkm1ikvsatc2[35];
wire z_hjy_5 = xlkm1ikvsatc2[36];
wire f9ojncwk = xlkm1ikvsatc2[37];
wire chwsbsq = xlkm1ikvsatc2[38];

wire [64-1:0] qi8_x06autspcyhhv;
assign qi8_x06autspcyhhv = ({64{pldtey61}} & {8{amgi_rqhtd007[7:0]}})
                        | ({64{vribxr_dbn}} & {8{amgi_rqhtd007[15:8]}})
                        | ({64{l5bnwm}} & {8{amgi_rqhtd007[23:16]}})
                        | ({64{lgnvbn}} & {8{amgi_rqhtd007[31:24]}})
                        | ({64{ksxzc99stv9}} & {8{amgi_rqhtd007[39:32]}})
                        | ({64{z_hjy_5}} & {8{amgi_rqhtd007[47:40]}})
                        | ({64{f9ojncwk}} & {8{amgi_rqhtd007[55:48]}})
                        | ({64{chwsbsq}} & {8{amgi_rqhtd007[63:56]}})
                        ;
wire zid3nz9u293bss6f4 = pldtey61 | vribxr_dbn | l5bnwm | lgnvbn | ksxzc99stv9 | z_hjy_5 | f9ojncwk | chwsbsq;                        





assign nb3w1rq_ny95rvrt = ({64{zby8wjkievope63}}   & huf4d5e5ey8_pj9r6_   ) |
                         ({64{cg_xvkpcb5oe4ov3r}} & p7e55yl2xz_s76csdl ) | 
                         ({64{ccm19fkdl1_0ex2}}   & qyh4fb808wpe28g8   ) | 
                         ({64{uq3eiceihlgu}}     & xx_4lcsv8bjm23ylo     ) | 
                         ({64{pfj780v6il2rtp}}     & k69l77w397qhwjeh     ) | 
                         ({64{gkjybnhfjsie3o}}   & slmojwuw5628djvr     ) | 
                         ({64{dzs4lvfhrbn6q}}     & n8v1vqp24ko3fof     ) | 
                         ({64{ut1dkcj1azkbznfp}}   & lfkclmsw9nw8cco_8c   ) |
                         ({64{z0v1bqkq5qn284wu}}   & q96ft3lmyjaeecp_2x45p   ) |
                         ({64{zid3nz9u293bss6f4}}   & qi8_x06autspcyhhv   )  
                         ;

assign vjkz8n6i44pc7o = zby8wjkievope63 & lkoe_jcrsl9h3;    



























endmodule




















module lxot_pmljpjs9pco4am4pfh5r(
    input oyxjs3av0z67vqd9z93,
    input laksv6w2w3g85egjh,
    input jj1e19z04mdd1903k6,
    input obyenny15k41m98a7jhajt,
    input b43ixz6gjo_3lsem91csma,
    input i23hpo2hianl9_xpewemf,
    input l_mrsjnfjwcw23l,
    input t124x7d61613qbluy3,
    input xbbag3r7y2il4kz_fdcb,
    input chgsl3e3omcgzcmhcdwnd9,
    input [63:0] usrh37qm6nz8yamj6_h_pmbv5,
    input [63:0] mipc_c8bfwk8khoqgtsj65f1f,
    input [63:0] pm3m6aucefl9oas0vqgwfm,
    input [63:0] yc5f_bw94gu1iari4qpmo269z,
    output [64-1:0] k6c8aiwomjglm9ok9zt4wb, 
    output etcizv32c63_xdl3f60 
);



  wire [31:0] kjjn1ogtam6o58b;                
  wire [31:0] ou8kz8uo9vsrehd;                
  wire [31:0] px82_aza1j05o;                
  wire [31:0] fqnmhf1gsvfiaq_ir;                

  wire [7:0] ppuytgyus4cq5ss;
  assign  ppuytgyus4cq5ss[0] = oyxjs3av0z67vqd9z93   & ((~usrh37qm6nz8yamj6_h_pmbv5[15]) & usrh37qm6nz8yamj6_h_pmbv5[14]);
  assign  ppuytgyus4cq5ss[1] = oyxjs3av0z67vqd9z93   & ((~usrh37qm6nz8yamj6_h_pmbv5[31]) & usrh37qm6nz8yamj6_h_pmbv5[30]);
  assign  ppuytgyus4cq5ss[2] = oyxjs3av0z67vqd9z93   & ((~usrh37qm6nz8yamj6_h_pmbv5[47]) & usrh37qm6nz8yamj6_h_pmbv5[46]);
  assign  ppuytgyus4cq5ss[3] = oyxjs3av0z67vqd9z93   & ((~usrh37qm6nz8yamj6_h_pmbv5[63]) & usrh37qm6nz8yamj6_h_pmbv5[62]);
  assign  ppuytgyus4cq5ss[4] = laksv6w2w3g85egjh & ((~mipc_c8bfwk8khoqgtsj65f1f[15]) & mipc_c8bfwk8khoqgtsj65f1f[14]);
  assign  ppuytgyus4cq5ss[5] = laksv6w2w3g85egjh & ((~mipc_c8bfwk8khoqgtsj65f1f[31]) & mipc_c8bfwk8khoqgtsj65f1f[30]);
  assign  ppuytgyus4cq5ss[6] = laksv6w2w3g85egjh & ((~mipc_c8bfwk8khoqgtsj65f1f[47]) & mipc_c8bfwk8khoqgtsj65f1f[46]);
  assign  ppuytgyus4cq5ss[7] = laksv6w2w3g85egjh & ((~mipc_c8bfwk8khoqgtsj65f1f[63]) & mipc_c8bfwk8khoqgtsj65f1f[62]);
  assign kjjn1ogtam6o58b[7:0]    = {8{oyxjs3av0z67vqd9z93}} & (ppuytgyus4cq5ss[0] ? 8'h7f : usrh37qm6nz8yamj6_h_pmbv5[14:7] );
  assign kjjn1ogtam6o58b[15:8]   = {8{oyxjs3av0z67vqd9z93}} & (ppuytgyus4cq5ss[1] ? 8'h7f : usrh37qm6nz8yamj6_h_pmbv5[30:23]); 
  assign kjjn1ogtam6o58b[23:16]  = {8{oyxjs3av0z67vqd9z93}} & (ppuytgyus4cq5ss[2] ? 8'h7f : usrh37qm6nz8yamj6_h_pmbv5[46:39]);
  assign kjjn1ogtam6o58b[31:24]  = {8{oyxjs3av0z67vqd9z93}} & (ppuytgyus4cq5ss[3] ? 8'h7f : usrh37qm6nz8yamj6_h_pmbv5[62:55]);
  assign ou8kz8uo9vsrehd[7:0]    = {8{laksv6w2w3g85egjh}} & (ppuytgyus4cq5ss[4] ? 8'h7f : mipc_c8bfwk8khoqgtsj65f1f[14:7] );
  assign ou8kz8uo9vsrehd[15:8]   = {8{laksv6w2w3g85egjh}} & (ppuytgyus4cq5ss[5] ? 8'h7f : mipc_c8bfwk8khoqgtsj65f1f[30:23]); 
  assign ou8kz8uo9vsrehd[23:16]  = {8{laksv6w2w3g85egjh}} & (ppuytgyus4cq5ss[6] ? 8'h7f : mipc_c8bfwk8khoqgtsj65f1f[46:39]);
  assign ou8kz8uo9vsrehd[31:24]  = {8{laksv6w2w3g85egjh}} & (ppuytgyus4cq5ss[7] ? 8'h7f : mipc_c8bfwk8khoqgtsj65f1f[62:55]);

  wire [3:0] vlf9vi0glv438el76vu;
  assign  vlf9vi0glv438el76vu[0] =   jj1e19z04mdd1903k6 & ((~usrh37qm6nz8yamj6_h_pmbv5[31]) &  usrh37qm6nz8yamj6_h_pmbv5[30]);
  assign  vlf9vi0glv438el76vu[1] =   b43ixz6gjo_3lsem91csma & ((~usrh37qm6nz8yamj6_h_pmbv5[63]) &  usrh37qm6nz8yamj6_h_pmbv5[62]);
  assign  vlf9vi0glv438el76vu[2] =   b43ixz6gjo_3lsem91csma & ((~mipc_c8bfwk8khoqgtsj65f1f[31]) &  mipc_c8bfwk8khoqgtsj65f1f[30]);
  assign  vlf9vi0glv438el76vu[3] =   b43ixz6gjo_3lsem91csma & ((~mipc_c8bfwk8khoqgtsj65f1f[63]) &  mipc_c8bfwk8khoqgtsj65f1f[62]); 

  assign px82_aza1j05o[15:0]  =  {16{jj1e19z04mdd1903k6}} & (vlf9vi0glv438el76vu[0] ? 16'h7fff : usrh37qm6nz8yamj6_h_pmbv5[30:15]);

  assign px82_aza1j05o[31:16] = ({16{b43ixz6gjo_3lsem91csma}} & (vlf9vi0glv438el76vu[1] ? 16'h7fff : usrh37qm6nz8yamj6_h_pmbv5[62:47]))
                              | ({16{i23hpo2hianl9_xpewemf &  px82_aza1j05o[15]}})
                              ;

  assign fqnmhf1gsvfiaq_ir[15:0]  = ({16{b43ixz6gjo_3lsem91csma}} & (vlf9vi0glv438el76vu[2] ? 16'h7fff : mipc_c8bfwk8khoqgtsj65f1f[30:15]))
                                | ({16{i23hpo2hianl9_xpewemf &  px82_aza1j05o[15]}})
                                ;
  assign fqnmhf1gsvfiaq_ir[31:16] =  ({16{b43ixz6gjo_3lsem91csma}} & (vlf9vi0glv438el76vu[3] ? 16'h7fff : mipc_c8bfwk8khoqgtsj65f1f[62:47]))
                                |  ({16{i23hpo2hianl9_xpewemf &  px82_aza1j05o[15]}})
                                ;


  wire [1:0] wl89ragxbngypbuube; 
  assign wl89ragxbngypbuube[0] = l_mrsjnfjwcw23l & ((~usrh37qm6nz8yamj6_h_pmbv5[31]) & usrh37qm6nz8yamj6_h_pmbv5[30]);
  assign wl89ragxbngypbuube[1] = t124x7d61613qbluy3 & ((~mipc_c8bfwk8khoqgtsj65f1f[31]) & mipc_c8bfwk8khoqgtsj65f1f[30]);



  wire [31:0] t9amokzo0kvsc0 =   {32{l_mrsjnfjwcw23l}} & (wl89ragxbngypbuube[0] ? 32'h7fffffff : {usrh37qm6nz8yamj6_h_pmbv5[30:0],1'b0});
  wire [31:0] o3j1m8xuh_ttqj1x0 =   {32{t124x7d61613qbluy3}} & (wl89ragxbngypbuube[1] ? 32'h7fffffff : {mipc_c8bfwk8khoqgtsj65f1f[30:0],1'b0});


  wire [32-1:0] q32s364d3mb118st6wa   = kjjn1ogtam6o58b | px82_aza1j05o | t9amokzo0kvsc0;
  wire [32-1:0] lxxferqtffzn5m_3ksu = ou8kz8uo9vsrehd | fqnmhf1gsvfiaq_ir |  o3j1m8xuh_ttqj1x0;
 
  assign etcizv32c63_xdl3f60 = (|ppuytgyus4cq5ss) | (|vlf9vi0glv438el76vu) | (|wl89ragxbngypbuube);

  wire [32-1:0] jso0sqe03do   = usrh37qm6nz8yamj6_h_pmbv5[31:0];
  wire [32-1:0] fioukloavng4sc = usrh37qm6nz8yamj6_h_pmbv5[63:32];

  wire [32-1:0] k2exu2r61fdq62e6tmt   = xbbag3r7y2il4kz_fdcb   ? q32s364d3mb118st6wa   : jso0sqe03do;
  wire [32-1:0] b3ejb414ewpnoqb1s4tdm4 = chgsl3e3omcgzcmhcdwnd9 ? lxxferqtffzn5m_3ksu : fioukloavng4sc;
  assign k6c8aiwomjglm9ok9zt4wb = {b3ejb414ewpnoqb1s4tdm4,k2exu2r61fdq62e6tmt};

endmodule
                       





















module qhqypfyt2lgewc2ne9xw(

  
  
  
  input [105-1:0] a4p3huz_qaf92as,
  input [105-1:0] e4_5otstd9ttd5eebgmf,
  input [50-1:0] n6izg3jvgts,
  input [64-1:0] amgi_rqhtd007,
  input [64-1:0] g7tawq8tp6,
  output w363n7ci30h3kw2g1oktlj1puysbju, 
  output lygqe2977b3fd_0eit3wg_nnfirn, 
  output th583ebkp2cj56crsivefzygk81o65_h2, 
  output vz2rm7lc9ctulrdhe1kv8wdmobft, 
  output hlmhgsbtxsmi7y1a7oshnntydp27pj,
  output dshcfm3k8zhyftxq_xw9j106j59z7notf,
  output [63 : 0] usrh37qm6nz8yamj6_h_pmbv5,           
  output [63 : 0] mipc_c8bfwk8khoqgtsj65f1f,           
  output [63 : 0] pm3m6aucefl9oas0vqgwfm,           
  output [63 : 0] yc5f_bw94gu1iari4qpmo269z,           
  output gdebc5b6o6bv57ax1bw
  );


  wire s7g459       = a4p3huz_qaf92as[15]; 
  wire xlr2qc65_      = 1'b0;
  wire pftfitai1lu     = 1'b0;
  wire scq1d7kkv5gs      = a4p3huz_qaf92as[16]; 
  wire wb1h98355      = a4p3huz_qaf92as[9];
  wire ko179gi1u      = a4p3huz_qaf92as[17];
  wire m5ne7y3kl2      = a4p3huz_qaf92as[18];
  wire gi8jcn9      = a4p3huz_qaf92as[19];
  wire crgxw_h6k      = a4p3huz_qaf92as[20];
  wire lsg8wa99uix9      = a4p3huz_qaf92as[21];
  wire qdf_fu8f      = a4p3huz_qaf92as[22];
  wire uttgo7lrg     = a4p3huz_qaf92as[10];
  wire nv4o0dey0     = a4p3huz_qaf92as[5];
  wire va5gdfkqpm56v7    = a4p3huz_qaf92as[6];
  wire cf8eoeq2c     = a4p3huz_qaf92as[7];
  wire p50g8hfzog    = a4p3huz_qaf92as[8];
  wire j33bi1i7w      = a4p3huz_qaf92as[11];
  wire c2d0jswv     = a4p3huz_qaf92as[12];
  wire qq9ppwd9      = a4p3huz_qaf92as[13];
  wire tdqo_isxb8_y     = a4p3huz_qaf92as[14];
  wire ytse6qk3     = e4_5otstd9ttd5eebgmf[48];
  wire lldmuweh65     = e4_5otstd9ttd5eebgmf[49];
  wire zqew83r8d     = e4_5otstd9ttd5eebgmf[50];
  wire uualc9afpol     = e4_5otstd9ttd5eebgmf[7];
  wire qm1du4l3      = e4_5otstd9ttd5eebgmf[8];
  wire a63upddr     = e4_5otstd9ttd5eebgmf[9];
  wire jyts2vkzi24kms    = e4_5otstd9ttd5eebgmf[10];
  wire l7n1yzahgthjb     = e4_5otstd9ttd5eebgmf[11];
  wire dfh3b4t_     = e4_5otstd9ttd5eebgmf[12];
  wire q1l2has7i4yu     = e4_5otstd9ttd5eebgmf[13];
  wire pszkdprqk6epwd    = e4_5otstd9ttd5eebgmf[14];
  wire pbwpday5027k     = e4_5otstd9ttd5eebgmf[15];
  wire lgy1y5tai    = e4_5otstd9ttd5eebgmf[16];
  wire n5cih6basb    = e4_5otstd9ttd5eebgmf[17];
  wire p4ew2ern4ea8      = e4_5otstd9ttd5eebgmf[6];
  wire jh6b6i12xnr0     = e4_5otstd9ttd5eebgmf[5];
  wire dota0x0h6ai5na    = e4_5otstd9ttd5eebgmf[18];
  wire sl6afay324me    = e4_5otstd9ttd5eebgmf[19];
  wire zi97mwha9ela   = e4_5otstd9ttd5eebgmf[20];
  wire cva1rq8nyf3    = e4_5otstd9ttd5eebgmf[21];
  wire b4shesc7j0liph   = e4_5otstd9ttd5eebgmf[22];
  wire egxho2viil87     = e4_5otstd9ttd5eebgmf[23];
  wire kqj6ekeqi0    = e4_5otstd9ttd5eebgmf[24];
  wire yd8mqaqh5       = e4_5otstd9ttd5eebgmf[25];
  wire khqacvet      = e4_5otstd9ttd5eebgmf[26];
  wire eumjbmutd       = e4_5otstd9ttd5eebgmf[27];
  wire hpbnc6go      = e4_5otstd9ttd5eebgmf[28];
  wire c586vep6      = e4_5otstd9ttd5eebgmf[29];
  wire trik6is2rd6m      = e4_5otstd9ttd5eebgmf[30];
  wire z7vkp91kvo      = e4_5otstd9ttd5eebgmf[31];
  wire dd0zqlm      = e4_5otstd9ttd5eebgmf[32];
  wire drfueow8g      = e4_5otstd9ttd5eebgmf[33];
  wire emvuyj8q5978k     = e4_5otstd9ttd5eebgmf[34];
  wire tzu0chnkec8      = e4_5otstd9ttd5eebgmf[35];
  wire w52f9xwl     = e4_5otstd9ttd5eebgmf[36];
  wire pb0jnx9gx     = e4_5otstd9ttd5eebgmf[37];
  wire dikgckhr      = e4_5otstd9ttd5eebgmf[38];
  wire nnhhc_ndfd     = e4_5otstd9ttd5eebgmf[39];
  wire l37c86_r      = e4_5otstd9ttd5eebgmf[40];
  wire a619145es      = e4_5otstd9ttd5eebgmf[41];
  wire agmkl2blti1    = e4_5otstd9ttd5eebgmf[42];
  wire wlxmne8wur     = e4_5otstd9ttd5eebgmf[43];
  wire pbgu2zjwf_     = e4_5otstd9ttd5eebgmf[44];
  wire aub52c3h     = e4_5otstd9ttd5eebgmf[45];
  wire u5qia7e705cb    = e4_5otstd9ttd5eebgmf[46];
  wire ykb5bh5g8d    = e4_5otstd9ttd5eebgmf[47];
  wire ql35edzw8pm       = e4_5otstd9ttd5eebgmf[51];
  wire kbxabqgwv9x8     = e4_5otstd9ttd5eebgmf[52];
  wire zqha84xel8     = e4_5otstd9ttd5eebgmf[53];
  wire uif2kv76     = e4_5otstd9ttd5eebgmf[54];
  wire ag7xsrfle7axh     = e4_5otstd9ttd5eebgmf[55];
  wire kmbjany88n1_0a    = e4_5otstd9ttd5eebgmf[56];
  wire lz6wwdpjxrj7e_    = e4_5otstd9ttd5eebgmf[57];
  wire kudyj9anu     = e4_5otstd9ttd5eebgmf[58];
  wire k2k_g5ru4q3vk    = e4_5otstd9ttd5eebgmf[59];
  wire faxp_tntmr8w     = e4_5otstd9ttd5eebgmf[60];
  wire cjtfl1k8q7376     = e4_5otstd9ttd5eebgmf[61];
  wire kbf5wps3bwl     = e4_5otstd9ttd5eebgmf[62];
  wire pqkp66hss2hu     = e4_5otstd9ttd5eebgmf[63];
  wire vyvkpez4tk5    = e4_5otstd9ttd5eebgmf[64];
  wire p1nfq2d77    = e4_5otstd9ttd5eebgmf[65];
  wire k6v0y53i3v03q     = e4_5otstd9ttd5eebgmf[66];
  wire mf7yezsyfa     = e4_5otstd9ttd5eebgmf[67];
  wire mw107xxcio4xz     = e4_5otstd9ttd5eebgmf[96];
  wire mp8ovnj      = e4_5otstd9ttd5eebgmf[97];
  wire i6ul4edu28m6     = e4_5otstd9ttd5eebgmf[98];
  wire ct0bff_7      = e4_5otstd9ttd5eebgmf[99];
  wire axpllj15ze9      = e4_5otstd9ttd5eebgmf[100];
  wire ojp0rsxys5     = e4_5otstd9ttd5eebgmf[101];
  wire rpc06tnfa_u     = e4_5otstd9ttd5eebgmf[102];
  wire ix_p044rqd     = e4_5otstd9ttd5eebgmf[103];
  wire lmc5kuujz1ue    = e4_5otstd9ttd5eebgmf[104];
  wire fme237kyf6i    = e4_5otstd9ttd5eebgmf[68];
  wire jtt_4jgy4r9a    = e4_5otstd9ttd5eebgmf[69];
  wire h_2kos5aq5l    = e4_5otstd9ttd5eebgmf[70];
  wire u0_9klg0dwfbyu    = e4_5otstd9ttd5eebgmf[71];
  wire ltxfa9scjc    = e4_5otstd9ttd5eebgmf[72];
  wire w9y5m7h97ob9v    = e4_5otstd9ttd5eebgmf[73];
  wire ebjrf08wpu     = e4_5otstd9ttd5eebgmf[74 ];
  wire lgd_52ezs     = e4_5otstd9ttd5eebgmf[75 ];
  wire sdg_mdde53r     = e4_5otstd9ttd5eebgmf[76 ];
  wire es5f1193zfutlpl   = e4_5otstd9ttd5eebgmf[77];   
  wire r789g6d1e6_   = e4_5otstd9ttd5eebgmf[78];   
  wire fgcvletq0c   = e4_5otstd9ttd5eebgmf[79];   
  wire npnmecyw6yf8x    = e4_5otstd9ttd5eebgmf[80 ];   
  wire zt38wq5knk    = e4_5otstd9ttd5eebgmf[81 ];   
  wire nksarbtyv7d3    = e4_5otstd9ttd5eebgmf[82 ];   
  wire i88x9z6wh1g    = e4_5otstd9ttd5eebgmf[83 ];   
  wire k7p4lhmq6ip   = e4_5otstd9ttd5eebgmf[84];   
  wire bg30eiom3ga7     = e4_5otstd9ttd5eebgmf[85  ];   
  wire fb9u6xhxy    = e4_5otstd9ttd5eebgmf[86 ];   
  wire qpgrwyn1vt    = e4_5otstd9ttd5eebgmf[87 ];   
  wire h34ave6xbfid4v   = e4_5otstd9ttd5eebgmf[88];   
  wire bltyctxgbkrkac4   = e4_5otstd9ttd5eebgmf[89];   
  wire t4t3u8572n8    = e4_5otstd9ttd5eebgmf[90 ];   
  wire aqe95jz9p48m21   = e4_5otstd9ttd5eebgmf[91];   
  wire jdck4rxqtx7zn     = e4_5otstd9ttd5eebgmf[92  ];   
  wire vb4fv39_hqam3    = e4_5otstd9ttd5eebgmf[93 ];   
  wire hkx0hr49lgrsxh    = e4_5otstd9ttd5eebgmf[94 ];   
        

  wire jl5uafxavxn4ffun =  n6izg3jvgts[10];


  wire b4wi1969mw9n534p = n6izg3jvgts[9];
  wire k5795hlk3_q   =  n6izg3jvgts[11];

  wire x1kaexv26aa2fd_7nz8w2t = n6izg3jvgts[13];
                                
                                


  wire hf3_u19xhtm47jygm346ih5592f = n6izg3jvgts[28]; 
  wire niiot38ff0zsxxncd0u_5fljm__dl = n6izg3jvgts[27];
  wire pm3poaltg6mtmffm_87yhorfj9eort_ = n6izg3jvgts[29]; 
  wire hxv8akm9tnbagx      = n6izg3jvgts[14];



  wire [31:0] tt2c87mcx6t7l4nazopbi8tufyyx2a;
  wire [31:0] hexy9i9cx278g_gq1xa85w735098s;
  wire [31:0] scnc2o0onmfzkunfbqlwf96_dqibfx5;
  wire [31:0] ofydji25el_rhpy7qm466hp1a414dn;

  wire [64-1:0] u3sluj7j2sehfsy = ({64{k5795hlk3_q}} & amgi_rqhtd007)
                                      ;
  wire [64-1:0] xtl841cb0zo01b1f = ({64{k5795hlk3_q}} & g7tawq8tp6)
                                      ;

  wire y1fgyae1uzj7ujuxqi3znyfnbb19hjsl = n6izg3jvgts[30];
  wire sfwi4o77fiwv1s1kb4mmixcewjetb_1 = n6izg3jvgts[31];
  wire oboq9ew68wxfv1zbbzbw6ovxumvp4ms = n6izg3jvgts[32];
  wire ozipqe_4brzi2opcs5pi232jtqiu7_m6kuv = n6izg3jvgts[33];
  wire imwjfayr9ztr86owxp26dtq0onjtd6dp = n6izg3jvgts[34];
  wire n38usa0n35mgmntamkuxh2l5pd2gcwghz = n6izg3jvgts[35];
  wire gm3156cuu5w0z0iabqd970k351i652n1u = n6izg3jvgts[36];
  wire n93vkxau7xxglljhnhsxg_4jddx13kcy = n6izg3jvgts[37];
  wire t88i3logg39o9_7fi_4qgfve8slrofj4j = n6izg3jvgts[38];
  wire e7ilxivhp9g8urh1klgvakcpqfmwjd5tw = n6izg3jvgts[39];
  wire hhf5vk7i4v5m5s0diu0q2m6pmxzvm7zeyiv7r = n6izg3jvgts[40];
  wire e9gctcgx_15frdmbcrevvtf_2lldmasrmr9gp = n6izg3jvgts[41];
  wire wj4suc8dinc_9d5409y_to9toxtea5b3afqoc = n6izg3jvgts[42];
  wire o44zcer7fjl2e666o3w3zxacak78idnwavnn = n6izg3jvgts[43];
  wire iue4b0u82l97gr25u35a4wkzrr64s8kyxgwm = n6izg3jvgts[44];
  wire mr9h2nuumis0_vx1kbbu849xvlx89du725kw = n6izg3jvgts[45];
  wire k0ly3yt_k96klqrmoe2jg2fjd6qz2edc5j87l = n6izg3jvgts[46];
  wire tivrapwmioo0momgw9hmmlzhrcqyoa8a6wdu2yh = n6izg3jvgts[47];
  wire s89z9cptleb2csl1iyj0lg_altgx5k1f6316m1h = n6izg3jvgts[48];
  wire oy_6emad9374dtcw5eu89i4o6o5kuiqu26hsgcb = n6izg3jvgts[49];



  assign tt2c87mcx6t7l4nazopbi8tufyyx2a   =
                                     ({32{y1fgyae1uzj7ujuxqi3znyfnbb19hjsl}} & {amgi_rqhtd007[31:0]})
                                   | ({32{sfwi4o77fiwv1s1kb4mmixcewjetb_1}} & {{16{amgi_rqhtd007[15]}},amgi_rqhtd007[15:0]})
                                   | ({32{oboq9ew68wxfv1zbbzbw6ovxumvp4ms}} & {{16{amgi_rqhtd007[31]}},amgi_rqhtd007[31:16]})
                                   | ({32{ozipqe_4brzi2opcs5pi232jtqiu7_m6kuv}} & {{16{g7tawq8tp6[15]}},g7tawq8tp6[15:0]})
                                   | ({32{imwjfayr9ztr86owxp26dtq0onjtd6dp}} & {amgi_rqhtd007[63:32]})
                                   ;

  



  assign hexy9i9cx278g_gq1xa85w735098s   = 
                                     ({32{n38usa0n35mgmntamkuxh2l5pd2gcwghz}} & {g7tawq8tp6[31:0]})
                                   | ({32{gm3156cuu5w0z0iabqd970k351i652n1u}} & {{16{g7tawq8tp6[15]}},g7tawq8tp6[15:0]})
                                   | ({32{n93vkxau7xxglljhnhsxg_4jddx13kcy}} & {{16{g7tawq8tp6[31]}},g7tawq8tp6[31:16]})
                                   | ({32{t88i3logg39o9_7fi_4qgfve8slrofj4j}} & {{15{g7tawq8tp6[15]}},g7tawq8tp6[15:0],1'b0})
                                   | ({32{e7ilxivhp9g8urh1klgvakcpqfmwjd5tw}} & {{15{g7tawq8tp6[31]}},g7tawq8tp6[31:16],1'b0})
                                   ;


  assign scnc2o0onmfzkunfbqlwf96_dqibfx5 =
                                     ({32{hhf5vk7i4v5m5s0diu0q2m6pmxzvm7zeyiv7r}} & {amgi_rqhtd007[63:32]})
                                   | ({32{e9gctcgx_15frdmbcrevvtf_2lldmasrmr9gp}} & {{16{amgi_rqhtd007[47]}},amgi_rqhtd007[47:32]})
                                   | ({32{wj4suc8dinc_9d5409y_to9toxtea5b3afqoc}} & {{16{amgi_rqhtd007[63]}},amgi_rqhtd007[63:48]})
                                   | ({32{o44zcer7fjl2e666o3w3zxacak78idnwavnn}} & {{16{g7tawq8tp6[47]}},g7tawq8tp6[47:32]})
                                   | ({32{iue4b0u82l97gr25u35a4wkzrr64s8kyxgwm}} & {amgi_rqhtd007[31:0]})
                                     ;

  assign ofydji25el_rhpy7qm466hp1a414dn =
                                     ({32{mr9h2nuumis0_vx1kbbu849xvlx89du725kw}} & {g7tawq8tp6[63:32]})
                                   | ({32{k0ly3yt_k96klqrmoe2jg2fjd6qz2edc5j87l}} & {{16{g7tawq8tp6[47]}},g7tawq8tp6[47:32]})
                                   | ({32{tivrapwmioo0momgw9hmmlzhrcqyoa8a6wdu2yh}} & {{16{g7tawq8tp6[63]}},g7tawq8tp6[63:48]})
                                   | ({32{s89z9cptleb2csl1iyj0lg_altgx5k1f6316m1h}} & {{15{g7tawq8tp6[47]}},g7tawq8tp6[47:32],1'b0})
                                   | ({32{oy_6emad9374dtcw5eu89i4o6o5kuiqu26hsgcb}} & {{15{g7tawq8tp6[63]}},g7tawq8tp6[63:48],1'b0})
                                     ;

  

  assign gdebc5b6o6bv57ax1bw = n6izg3jvgts[0];

  wire fxk_v35ltu7y0_q6aadrtlvrl = agmkl2blti1;                           


  e2pg9lpkkc1p07id6ljjmll1r hsorf_so0wrjcn5p7gyhidxo(
    .u3sluj7j2sehfsy              (u3sluj7j2sehfsy),
    .xtl841cb0zo01b1f              (xtl841cb0zo01b1f),
    .tt2c87mcx6t7l4nazopbi8tufyyx2a  (tt2c87mcx6t7l4nazopbi8tufyyx2a),
    .hexy9i9cx278g_gq1xa85w735098s  (hexy9i9cx278g_gq1xa85w735098s),
    .scnc2o0onmfzkunfbqlwf96_dqibfx5(scnc2o0onmfzkunfbqlwf96_dqibfx5),
    .ofydji25el_rhpy7qm466hp1a414dn(ofydji25el_rhpy7qm466hp1a414dn),
    .gdebc5b6o6bv57ax1bw           (gdebc5b6o6bv57ax1bw),
    .jl5uafxavxn4ffun               (jl5uafxavxn4ffun),
    .b4wi1969mw9n534p               (b4wi1969mw9n534p),
    .hf3_u19xhtm47jygm346ih5592f   (hf3_u19xhtm47jygm346ih5592f),
    .niiot38ff0zsxxncd0u_5fljm__dl (niiot38ff0zsxxncd0u_5fljm__dl),
    .pm3poaltg6mtmffm_87yhorfj9eort_(pm3poaltg6mtmffm_87yhorfj9eort_),
    .x1kaexv26aa2fd_7nz8w2t     (x1kaexv26aa2fd_7nz8w2t),
    .usrh37qm6nz8yamj6_h_pmbv5       (usrh37qm6nz8yamj6_h_pmbv5),
    .mipc_c8bfwk8khoqgtsj65f1f       (mipc_c8bfwk8khoqgtsj65f1f),
    .pm3m6aucefl9oas0vqgwfm       (pm3m6aucefl9oas0vqgwfm),
    .yc5f_bw94gu1iari4qpmo269z       (yc5f_bw94gu1iari4qpmo269z),
    .fxk_v35ltu7y0_q6aadrtlvrl     (fxk_v35ltu7y0_q6aadrtlvrl) 
  );


  wire [15:0] eerenuij1zyae3gifzsq3e6h6ahnp1 = ({16{(wlxmne8wur | pbgu2zjwf_
                                                  | u0_9klg0dwfbyu | ltxfa9scjc
                                                  | fme237kyf6i | jtt_4jgy4r9a 
                                                  | es5f1193zfutlpl | r789g6d1e6_
                                                  )}} & amgi_rqhtd007[15:0])
                                            | ({16{
                                                   aub52c3h
                                                 | w9y5m7h97ob9v | h_2kos5aq5l | fgcvletq0c
                                                  }} & amgi_rqhtd007[31:16])
                                            ; 
  wire [15:0] o6xi4lbf659woe65xbsqramzut382y72448ibsogc2 = ({16{( u0_9klg0dwfbyu | ltxfa9scjc | fme237kyf6i 
                                                           | jtt_4jgy4r9a | es5f1193zfutlpl | r789g6d1e6_)}} & amgi_rqhtd007[47:32])
                                                    | ({16{ w9y5m7h97ob9v | h_2kos5aq5l | fgcvletq0c }} & amgi_rqhtd007[63:48])
                                                    ; 

  wire [15:0] ad84kle0972tfpz4bzmhq3d_8pxu8_5         = ({16{(wlxmne8wur | sl6afay324me | zi97mwha9ela 
                                                          | ojp0rsxys5 | n5cih6basb
                                                          | u0_9klg0dwfbyu | fme237kyf6i | es5f1193zfutlpl
                                                          )}} & g7tawq8tp6[15:0])
                                                    | ({16{aub52c3h | pbgu2zjwf_ | cva1rq8nyf3 
                                                         | b4shesc7j0liph | rpc06tnfa_u | dota0x0h6ai5na
                                                          | ltxfa9scjc | jtt_4jgy4r9a | r789g6d1e6_
                                                          | w9y5m7h97ob9v | h_2kos5aq5l | fgcvletq0c
                                                         }} & g7tawq8tp6[31:16])
                                                    ; 
  wire [15:0] v_1f43tv2phai790a5k7t0o73vdl2g2a8vkqdw5eth = ({16{( sl6afay324me | zi97mwha9ela 
                                                           | ojp0rsxys5 | n5cih6basb
                                                           | u0_9klg0dwfbyu | fme237kyf6i | es5f1193zfutlpl
                                                            )}} & g7tawq8tp6[47:32])
                                                    | ({16{ cva1rq8nyf3 | b4shesc7j0liph 
                                                          | rpc06tnfa_u | dota0x0h6ai5na 
                                                          | ltxfa9scjc | jtt_4jgy4r9a | r789g6d1e6_
                                                          | w9y5m7h97ob9v | h_2kos5aq5l | fgcvletq0c
                                                          }} & g7tawq8tp6[63:48])
                                                    ; 

  wire c68ttj4idrbl1pav4aj68wy3zype7cbg = (eerenuij1zyae3gifzsq3e6h6ahnp1 == 16'h8000);
  wire jb6hpl55u7jfxk7y6uky3_n0p2o8pxv5nwe = (ad84kle0972tfpz4bzmhq3d_8pxu8_5 == 16'h8000);
  wire hunxkdngkabivw0cufin9uxcecbp_60k08v = (amgi_rqhtd007[31:0] == 32'h80000000);
  wire a17_ebmjt2tcwty1g6cz8hj1o0a6u0y2rb = (g7tawq8tp6[31:0] == 32'h80000000);
  wire hhf1ceimjq8kjjpsou6s3mvvf0n72jdf_c9 = (o6xi4lbf659woe65xbsqramzut382y72448ibsogc2 == 16'h8000);
  wire cew8da95sd_55r5lzo4eboas9f1cynswrh = (v_1f43tv2phai790a5k7t0o73vdl2g2a8vkqdw5eth == 16'h8000);
  wire fh5aamygxzkui2he_rq32pa_b8abmhvrh_bs9q = (amgi_rqhtd007[63:32] == 32'h80000000);
  wire isr_e4xbysrx4yfled1d4k56rugd2r9g49 = (g7tawq8tp6[63:32] == 32'h80000000);
  assign w363n7ci30h3kw2g1oktlj1puysbju = (  hunxkdngkabivw0cufin9uxcecbp_60k08v &
                                   ( ((ojp0rsxys5 |rpc06tnfa_u   | n5cih6basb |dota0x0h6ai5na )   & jb6hpl55u7jfxk7y6uky3_n0p2o8pxv5nwe)  
                                   | ((i6ul4edu28m6 |jyts2vkzi24kms)                            & a17_ebmjt2tcwty1g6cz8hj1o0a6u0y2rb)
                                   ))
                                   ;
  assign th583ebkp2cj56crsivefzygk81o65_h2 = (fh5aamygxzkui2he_rq32pa_b8abmhvrh_bs9q &
                                   ( ((ojp0rsxys5 |rpc06tnfa_u   | n5cih6basb |dota0x0h6ai5na )   & cew8da95sd_55r5lzo4eboas9f1cynswrh)  
                                   | ((i6ul4edu28m6 |jyts2vkzi24kms)                            & isr_e4xbysrx4yfled1d4k56rugd2r9g49)
                                   ))
                                   ;
  assign hlmhgsbtxsmi7y1a7oshnntydp27pj = jb6hpl55u7jfxk7y6uky3_n0p2o8pxv5nwe & c68ttj4idrbl1pav4aj68wy3zype7cbg
                                    & (u0_9klg0dwfbyu | ltxfa9scjc | w9y5m7h97ob9v)
                                    ;
  assign dshcfm3k8zhyftxq_xw9j106j59z7notf = cew8da95sd_55r5lzo4eboas9f1cynswrh & hhf1ceimjq8kjjpsou6s3mvvf0n72jdf_c9
                                    & (u0_9klg0dwfbyu | ltxfa9scjc | w9y5m7h97ob9v)
                                    ;
  assign lygqe2977b3fd_0eit3wg_nnfirn  = jb6hpl55u7jfxk7y6uky3_n0p2o8pxv5nwe &
                                   ( (hunxkdngkabivw0cufin9uxcecbp_60k08v & (sl6afay324me | zi97mwha9ela |cva1rq8nyf3 |b4shesc7j0liph))
                                    |(c68ttj4idrbl1pav4aj68wy3zype7cbg & (wlxmne8wur | pbgu2zjwf_ | aub52c3h
                                                                        | fme237kyf6i | jtt_4jgy4r9a | h_2kos5aq5l
                                                                        | es5f1193zfutlpl | r789g6d1e6_ | fgcvletq0c
                                                                         ))
                                   );
  assign vz2rm7lc9ctulrdhe1kv8wdmobft  = cew8da95sd_55r5lzo4eboas9f1cynswrh &
                                   ( (fh5aamygxzkui2he_rq32pa_b8abmhvrh_bs9q & (sl6afay324me | zi97mwha9ela |cva1rq8nyf3 |b4shesc7j0liph))
                                   | (hhf1ceimjq8kjjpsou6s3mvvf0n72jdf_c9 & ( fme237kyf6i | jtt_4jgy4r9a | h_2kos5aq5l
                                                                           | es5f1193zfutlpl | r789g6d1e6_ | fgcvletq0c
                                                                           ))
                                   );

 
  

endmodule                                           

module opvhnxssc7yjqmd3 #(
  parameter onr7l = 106 
)(
  input [onr7l-1:0] frgfco,
  input [onr7l-1:0] ii,
  input [onr7l-1:0] fij51v,
  output [onr7l-1:0] c,
  output [onr7l-1:0] s 
);

assign s = (frgfco ^ ii) ^ fij51v;

wire [onr7l-1:0] oz7_y5 = (frgfco & ii) | (frgfco & fij51v) | (ii & fij51v);

assign c = {oz7_y5[onr7l-2:0], 1'b0};

endmodule

module gg0ubjxsd5riswv #(
    parameter onr7l = 106 
)(
  input [onr7l-1:0] frgfco,
  input [onr7l-1:0] ii,
  input [onr7l-1:0] fij51v,
  input [onr7l-1:0] cuzhl9,
  output [onr7l-1:0] c,
  output [onr7l-1:0] s 
);

   wire [onr7l-1:0] i885 = (frgfco & ii) | (ii & fij51v) | (frgfco & fij51v);
   wire [onr7l-1:0] smqrocit = {i885[onr7l-2:0], 1'b0};

   wire [onr7l-1:0] tqxp_8 = smqrocit ^ cuzhl9;
   wire [onr7l-1:0] ddaxu87 = (frgfco ^ ii) ^ fij51v;

   assign s = tqxp_8 ^ ddaxu87;

   wire [onr7l-1:0] hgtxv = (ddaxu87 & cuzhl9) |  (cuzhl9 & smqrocit) | (smqrocit & ddaxu87);

   assign c = {hgtxv[onr7l-2:0], 1'b0};

endmodule
                       





















module s20vasmduccat9_3(

  

  input[80-1:0]  pugy9o4i2pr3ns8yo3 ,
  input[80-1:0]  qg0gj_1bem7nt1wek5w2bc ,
  input[2:0]   wip5afkxmbs5dou  , 
  input[3:0]   dgvew5k86brk_8uip   , 
  input        phlh_dccd75w7xikxtg03 , 
  input        jqnqhlv1gjf2k3xg4 ,
  output[64-1:0] vvoozaywykiwmels   ,
  output[64-1:0] m50l82p03g15y_ehxthx1  ,
  output       hsvg_y2njolj1bl      


  );

  wire [80-1:0] duhacqzewc4p;
  wire [80-1:0] xt0_dl4l5jwlesp;
  wire [2:0]  pxscquhi78;
  wire [3:0]  ck6o6flrt;
  wire        lvhs9fkt_6d9;
  
  
  
  

  localparam wxbg7z6hn_1rfi1anz2 = 80+80+3+4+1;

  assign  {
    duhacqzewc4p
   ,xt0_dl4l5jwlesp
   ,pxscquhi78      
   ,ck6o6flrt      
   ,lvhs9fkt_6d9     
    }
    = 
        ({wxbg7z6hn_1rfi1anz2{jqnqhlv1gjf2k3xg4}} & {
             pugy9o4i2pr3ns8yo3 
            ,qg0gj_1bem7nt1wek5w2bc 
            ,wip5afkxmbs5dou 
            ,dgvew5k86brk_8uip 
            ,phlh_dccd75w7xikxtg03      
           })
        ;


  
  
  
  
  wire khqzwdn7t8_cfub9p = (ck6o6flrt == 4'b0000) & (pxscquhi78 == 3'b000) & lvhs9fkt_6d9;
  wire b6hhq101tety5ku7 = (ck6o6flrt == 4'b0000) & (pxscquhi78 == 3'b100) & lvhs9fkt_6d9;

  wire o9a1t19_k87qejl6jpfi   = ~duhacqzewc4p[78]   & duhacqzewc4p[77];
  wire pp2p4uy2pjiute0aisyq   = ~duhacqzewc4p[68]   & duhacqzewc4p[67];
  wire uldmmclkihym2tt40frjit2q   = ~duhacqzewc4p[58]   & duhacqzewc4p[57];
  wire ej44tix3xlo9b3ek8rnk935m   = ~duhacqzewc4p[48]   & duhacqzewc4p[47];
  wire f89mew8l_3vd3yfsgi2wzadp9   = ~duhacqzewc4p[38]   & duhacqzewc4p[37];
  wire fjpavfi27v774sm0uye3k   = ~duhacqzewc4p[28]   & duhacqzewc4p[27];
  wire cxpr5eviejhjiumtij5p9vb_   = ~duhacqzewc4p[18]   & duhacqzewc4p[17];
  wire z_xfo1ho0xh2ws9pfxze_   = ~duhacqzewc4p[8 ]   & duhacqzewc4p[7 ];

  
  wire vhivszyvssfd9yt_dbqzbbx   = duhacqzewc4p[78]   & ~duhacqzewc4p[77];
  wire c4lry4ezrmeprxk927cg   = duhacqzewc4p[68]   & ~duhacqzewc4p[67];
  wire u968xct45kalhavp7qadwy   = duhacqzewc4p[58]   & ~duhacqzewc4p[57];
  wire igcyyvmr2dcfu7h5mgrf35cg   = duhacqzewc4p[48]   & ~duhacqzewc4p[47];
  wire rtm_ujfus2gjnzom57x4   = duhacqzewc4p[38]   & ~duhacqzewc4p[37];
  wire s9uxc4pu0neakyknw1ryjr9wy   = duhacqzewc4p[28]   & ~duhacqzewc4p[27];
  wire iqibu_1drkoqe34m3rxsu1xj   = duhacqzewc4p[18]   & ~duhacqzewc4p[17];
  wire jzq5ma17wgzv_p7sihacj   = duhacqzewc4p[8 ]   & ~duhacqzewc4p[7 ];

  wire[64-1:0] utgqzem07taxie245 = {64{khqzwdn7t8_cfub9p | b6hhq101tety5ku7}} & {
        ({1'b0,{7{o9a1t19_k87qejl6jpfi}}}) | ({8{vhivszyvssfd9yt_dbqzbbx}} & 8'h80) | ({8{~o9a1t19_k87qejl6jpfi & ~vhivszyvssfd9yt_dbqzbbx}} & duhacqzewc4p[77:70]),
        ({1'b0,{7{pp2p4uy2pjiute0aisyq}}}) | ({8{c4lry4ezrmeprxk927cg}} & 8'h80) | ({8{~pp2p4uy2pjiute0aisyq & ~c4lry4ezrmeprxk927cg}} & duhacqzewc4p[67:60]),
        ({1'b0,{7{uldmmclkihym2tt40frjit2q}}}) | ({8{u968xct45kalhavp7qadwy}} & 8'h80) | ({8{~uldmmclkihym2tt40frjit2q & ~u968xct45kalhavp7qadwy}} & duhacqzewc4p[57:50]),
        ({1'b0,{7{ej44tix3xlo9b3ek8rnk935m}}}) | ({8{igcyyvmr2dcfu7h5mgrf35cg}} & 8'h80) | ({8{~ej44tix3xlo9b3ek8rnk935m & ~igcyyvmr2dcfu7h5mgrf35cg}} & duhacqzewc4p[47:40]),
        ({1'b0,{7{f89mew8l_3vd3yfsgi2wzadp9}}}) | ({8{rtm_ujfus2gjnzom57x4}} & 8'h80) | ({8{~f89mew8l_3vd3yfsgi2wzadp9 & ~rtm_ujfus2gjnzom57x4}} & duhacqzewc4p[37:30]),
        ({1'b0,{7{fjpavfi27v774sm0uye3k}}}) | ({8{s9uxc4pu0neakyknw1ryjr9wy}} & 8'h80) | ({8{~fjpavfi27v774sm0uye3k & ~s9uxc4pu0neakyknw1ryjr9wy}} & duhacqzewc4p[27:20]),
        ({1'b0,{7{cxpr5eviejhjiumtij5p9vb_}}}) | ({8{iqibu_1drkoqe34m3rxsu1xj}} & 8'h80) | ({8{~cxpr5eviejhjiumtij5p9vb_ & ~iqibu_1drkoqe34m3rxsu1xj}} & duhacqzewc4p[17:10]),
        ({1'b0,{7{z_xfo1ho0xh2ws9pfxze_}}}) | ({8{jzq5ma17wgzv_p7sihacj}} & 8'h80) | ({8{~z_xfo1ho0xh2ws9pfxze_ & ~jzq5ma17wgzv_p7sihacj}} & duhacqzewc4p[7 : 0])
       };


  wire bsc70kh_r2id7wwj7   =  (khqzwdn7t8_cfub9p | b6hhq101tety5ku7) & (
                              (o9a1t19_k87qejl6jpfi | pp2p4uy2pjiute0aisyq | uldmmclkihym2tt40frjit2q | ej44tix3xlo9b3ek8rnk935m | 
                               vhivszyvssfd9yt_dbqzbbx | c4lry4ezrmeprxk927cg | u968xct45kalhavp7qadwy | igcyyvmr2dcfu7h5mgrf35cg
                              ) | 
                              (f89mew8l_3vd3yfsgi2wzadp9 | fjpavfi27v774sm0uye3k | cxpr5eviejhjiumtij5p9vb_ | z_xfo1ho0xh2ws9pfxze_ | 
                               rtm_ujfus2gjnzom57x4 | s9uxc4pu0neakyknw1ryjr9wy | iqibu_1drkoqe34m3rxsu1xj | jzq5ma17wgzv_p7sihacj 
                              ));


  wire w3wxllzvry4npxh = bsc70kh_r2id7wwj7 
                   ;

  
  wire otvnx5pkt5aw = (ck6o6flrt == 4'b0001) & (pxscquhi78 == 3'b000) & lvhs9fkt_6d9;
  wire[64-1:0] mta9g3ta_8x7b3tqa = {64{otvnx5pkt5aw}} & {
                             ({8{~(duhacqzewc4p[78])}} & duhacqzewc4p[77:70]),
                             ({8{~(duhacqzewc4p[68])}} & duhacqzewc4p[67:60]),
                             ({8{~(duhacqzewc4p[58])}} & duhacqzewc4p[57:50]),
                             ({8{~(duhacqzewc4p[48])}} & duhacqzewc4p[47:40]),
                             ({8{~(duhacqzewc4p[38])}} & duhacqzewc4p[37:30]),
                             ({8{~(duhacqzewc4p[28])}} & duhacqzewc4p[27:20]),
                             ({8{~(duhacqzewc4p[18])}} & duhacqzewc4p[17:10]),
                             ({8{~(duhacqzewc4p[08])}} & duhacqzewc4p[07:00])};

  wire g1j_85l4zzhsb = otvnx5pkt5aw & (
                            duhacqzewc4p[78] | duhacqzewc4p[68] |duhacqzewc4p[58] |duhacqzewc4p[48] |
                            duhacqzewc4p[38] | duhacqzewc4p[28] |duhacqzewc4p[18] |duhacqzewc4p[8] 
                          );

  
  wire t9r50zrh89s7ztk = (ck6o6flrt == 4'b0001) & (pxscquhi78 == 3'b000) & ~lvhs9fkt_6d9;
  wire[64-1:0] uxo500z5tj5fa1j = {64{t9r50zrh89s7ztk}} & {
                              ({8{duhacqzewc4p[78]}} | duhacqzewc4p[77:70]),
                              ({8{duhacqzewc4p[68]}} | duhacqzewc4p[67:60]),
                              ({8{duhacqzewc4p[58]}} | duhacqzewc4p[57:50]),
                              ({8{duhacqzewc4p[48]}} | duhacqzewc4p[47:40]), 
                              ({8{duhacqzewc4p[38]}} | duhacqzewc4p[37:30]),
                              ({8{duhacqzewc4p[28]}} | duhacqzewc4p[27:20]),
                              ({8{duhacqzewc4p[18]}} | duhacqzewc4p[17:10]),
                              ({8{duhacqzewc4p[8 ]}} | duhacqzewc4p[7 :0] )};
  wire sy1xledv0xcnby3 = t9r50zrh89s7ztk &( 
                              (duhacqzewc4p[78] | duhacqzewc4p[68] |duhacqzewc4p[58] |duhacqzewc4p[48])|
                              (duhacqzewc4p[38] | duhacqzewc4p[28] |duhacqzewc4p[18] |duhacqzewc4p[8])
                            );

  
  wire ush3kg4qf4rchvxt    = (ck6o6flrt == 4'b0010) & (pxscquhi78 == 3'b001) & lvhs9fkt_6d9;
  wire q8cq6922962cszd1w1ibpy = (ck6o6flrt == 4'b0010) & (pxscquhi78 == 3'b101) & lvhs9fkt_6d9;
  
  wire j__th1ko8ws350t77itc = ~duhacqzewc4p[76] & duhacqzewc4p[75];
  wire qj6g_bez2aghkpev9c98nb = ~duhacqzewc4p[56] & duhacqzewc4p[55]; 
  wire hgdvb2s9bcix18l_idom = ~duhacqzewc4p[36] & duhacqzewc4p[35]; 
  wire b4f49ooi7xsqx0ie7ij6om = ~duhacqzewc4p[16] & duhacqzewc4p[15];

  
  wire w7fmivhceqetnlwmrdb = duhacqzewc4p[76] & ~duhacqzewc4p[75]; 
  wire lpxs5u9ssrumjxjriyl = duhacqzewc4p[56] & ~duhacqzewc4p[55];
  wire a9byi_8qwydluylgukur = duhacqzewc4p[36] & ~duhacqzewc4p[35]; 
  wire yjaozd_7pa5a173abfs_sd = duhacqzewc4p[16] & ~duhacqzewc4p[15];
  wire[64-1:0] i8hs0nk1rk1897rxqa = {64{ush3kg4qf4rchvxt | q8cq6922962cszd1w1ibpy}} & {
           (({1'b0,{15{j__th1ko8ws350t77itc}}}) | ({16{w7fmivhceqetnlwmrdb}} & 16'h8000) | ({16{~j__th1ko8ws350t77itc & ~w7fmivhceqetnlwmrdb}} & duhacqzewc4p[75:60])),
           (({1'b0,{15{qj6g_bez2aghkpev9c98nb}}}) | ({16{lpxs5u9ssrumjxjriyl}} & 16'h8000) | ({16{~qj6g_bez2aghkpev9c98nb & ~lpxs5u9ssrumjxjriyl}} & duhacqzewc4p[55:40])),
           (({1'b0,{15{hgdvb2s9bcix18l_idom}}}) | ({16{a9byi_8qwydluylgukur}} & 16'h8000) | ({16{~hgdvb2s9bcix18l_idom & ~a9byi_8qwydluylgukur}} & duhacqzewc4p[35:20])),
           (({1'b0,{15{b4f49ooi7xsqx0ie7ij6om}}}) | ({16{yjaozd_7pa5a173abfs_sd}} & 16'h8000) | ({16{~b4f49ooi7xsqx0ie7ij6om & ~yjaozd_7pa5a173abfs_sd}} & duhacqzewc4p[15:0 ]))
       };


  wire ogko3fr7jpuvbgb1mga   = (ush3kg4qf4rchvxt | q8cq6922962cszd1w1ibpy) & (
                               (j__th1ko8ws350t77itc | qj6g_bez2aghkpev9c98nb | w7fmivhceqetnlwmrdb | lpxs5u9ssrumjxjriyl) | 
                               (hgdvb2s9bcix18l_idom | b4f49ooi7xsqx0ie7ij6om | a9byi_8qwydluylgukur | yjaozd_7pa5a173abfs_sd)
                   ); 

  wire eio0m4xyepriqqk8wl5cvd =  1'b0; 
  wire mqo5q_91fbwq6p3r = ogko3fr7jpuvbgb1mga | eio0m4xyepriqqk8wl5cvd
                   ;  


  
  wire rtvs3qjdc4jbzne = (ck6o6flrt == 4'b0011) & (pxscquhi78 == 3'b001) & ~lvhs9fkt_6d9;
  wire[64-1:0] h59gmpawefdlc7erk9nq = {64{rtvs3qjdc4jbzne}} & {
                                ({16{duhacqzewc4p[76]}} | duhacqzewc4p[75:60]),({16{duhacqzewc4p[56]}} | duhacqzewc4p[55:40]), 
                                ({16{duhacqzewc4p[36]}} | duhacqzewc4p[35:20]),({16{duhacqzewc4p[16]}} | duhacqzewc4p[15:0 ])};
  wire e6tk2oatobnknne = rtvs3qjdc4jbzne & (
                         duhacqzewc4p[76] | duhacqzewc4p[56] |  
                         duhacqzewc4p[36] | duhacqzewc4p[16]
                        );
  
  
  wire u1xa8v9g_87fspma = (ck6o6flrt == 4'b0011) & (pxscquhi78 == 3'b001) & lvhs9fkt_6d9;
  wire[64-1:0] ek7dk29izkdtor =  {64{u1xa8v9g_87fspma}} & {
                                ({16{~(duhacqzewc4p[76])}} & duhacqzewc4p[75:60]),({16{~(duhacqzewc4p[56])}} & duhacqzewc4p[55:40]),
                                ({16{~(duhacqzewc4p[36])}} & duhacqzewc4p[35:20]),({16{~(duhacqzewc4p[16])}} & duhacqzewc4p[15:0 ])};

  wire suunz_obigrbmg8 = u1xa8v9g_87fspma & (
                               duhacqzewc4p[76] | duhacqzewc4p[56] |
                               duhacqzewc4p[36] | duhacqzewc4p[16]);


  
  wire megmtexkcejn7j4t    = (ck6o6flrt == 4'b0110) & (pxscquhi78 == 3'b000);
  wire v8g190egj7fkzr036wsol8d = (ck6o6flrt == 4'b0110) & (pxscquhi78 == 3'b100);
  wire qh5aqip9mi63us3tciq  = duhacqzewc4p[78] & (~duhacqzewc4p[77]);
  wire tjxuqq4zf_xju7a16bwou7  = duhacqzewc4p[68] & (~duhacqzewc4p[67]);
  wire vxbjkrru83c3walaqoyluwx  = duhacqzewc4p[58] & (~duhacqzewc4p[57]);
  wire mijs0a1t33e152qwd8di  = duhacqzewc4p[48] & (~duhacqzewc4p[47]);
  wire eshzy3_sakedorrju7wa  = duhacqzewc4p[38] & (~duhacqzewc4p[37]);
  wire rgz66rgl3mi4xotrz3  = duhacqzewc4p[28] & (~duhacqzewc4p[27]);
  wire mok9m6fs4y3hmgv5f6m  = duhacqzewc4p[18] & (~duhacqzewc4p[17]);
  wire fruw41264fd6a7t8sqk  = duhacqzewc4p[ 8] & (~duhacqzewc4p[ 7]);

  wire[64-1:0] qfnxty3b3r0wv5b_ = {64{megmtexkcejn7j4t | v8g190egj7fkzr036wsol8d}} & { 
     {1'b0,{7{qh5aqip9mi63us3tciq}}} | ({8{duhacqzewc4p[78] & duhacqzewc4p[77]}} & (~duhacqzewc4p[77:70])) | ({8{(~duhacqzewc4p[78]) & (~duhacqzewc4p[77])}} & duhacqzewc4p[77:70]) ,
     {1'b0,{7{tjxuqq4zf_xju7a16bwou7}}} | ({8{duhacqzewc4p[68] & duhacqzewc4p[67]}} & (~duhacqzewc4p[67:60])) | ({8{(~duhacqzewc4p[68]) & (~duhacqzewc4p[67])}} & duhacqzewc4p[67:60]) ,
     {1'b0,{7{vxbjkrru83c3walaqoyluwx}}} | ({8{duhacqzewc4p[58] & duhacqzewc4p[57]}} & (~duhacqzewc4p[57:50])) | ({8{(~duhacqzewc4p[58]) & (~duhacqzewc4p[57])}} & duhacqzewc4p[57:50]) ,
     {1'b0,{7{mijs0a1t33e152qwd8di}}} | ({8{duhacqzewc4p[48] & duhacqzewc4p[47]}} & (~duhacqzewc4p[47:40])) | ({8{(~duhacqzewc4p[48]) & (~duhacqzewc4p[47])}} & duhacqzewc4p[47:40]) , 
     {1'b0,{7{eshzy3_sakedorrju7wa}}} | ({8{duhacqzewc4p[38] & duhacqzewc4p[37]}} & (~duhacqzewc4p[37:30])) | ({8{(~duhacqzewc4p[38]) & (~duhacqzewc4p[37])}} & duhacqzewc4p[37:30]) ,
     {1'b0,{7{rgz66rgl3mi4xotrz3}}} | ({8{duhacqzewc4p[28] & duhacqzewc4p[27]}} & (~duhacqzewc4p[27:20])) | ({8{(~duhacqzewc4p[28]) & (~duhacqzewc4p[27])}} & duhacqzewc4p[27:20]) ,
     {1'b0,{7{mok9m6fs4y3hmgv5f6m}}} | ({8{duhacqzewc4p[18] & duhacqzewc4p[17]}} & (~duhacqzewc4p[17:10])) | ({8{(~duhacqzewc4p[18]) & (~duhacqzewc4p[17])}} & duhacqzewc4p[17:10]) ,
     {1'b0,{7{fruw41264fd6a7t8sqk}}} | ({8{duhacqzewc4p[ 8] & duhacqzewc4p[ 7]}} & (~duhacqzewc4p[7 :0 ])) | ({8{(~duhacqzewc4p[ 8]) & (~duhacqzewc4p[ 7])}} & duhacqzewc4p[7 :0 ]) };

  wire o0hw_mm_grdkap9ptct7 = (megmtexkcejn7j4t | v8g190egj7fkzr036wsol8d) &  
                       ( eshzy3_sakedorrju7wa  
                       | rgz66rgl3mi4xotrz3  
                       | mok9m6fs4y3hmgv5f6m  
                       | fruw41264fd6a7t8sqk
                       | qh5aqip9mi63us3tciq  
                       | tjxuqq4zf_xju7a16bwou7  
                       | vxbjkrru83c3walaqoyluwx  
                       | mijs0a1t33e152qwd8di
                       )
                       ;

  wire z8_ag3wbvbhcdp = o0hw_mm_grdkap9ptct7 
                 ;

  
  wire z03_wl6z1na1ebppos    = (ck6o6flrt == 4'b0110) & (pxscquhi78 == 3'b001);
  wire dl1k34qvje99ofpsjzadtq61  = (ck6o6flrt == 4'b0110) & (pxscquhi78 == 3'b101);
  wire ktbf6dfpqw7ullwvs0 = duhacqzewc4p[76] & (~duhacqzewc4p[75]);
  wire ryfbr1ol3w448dqtaictsz = duhacqzewc4p[56] & (~duhacqzewc4p[55]);
  wire o_j64jm_72wyhefzn9g7 = duhacqzewc4p[36] & (~duhacqzewc4p[35]);
  wire iktahd9pfcstthpcp_dnu = duhacqzewc4p[16] & (~duhacqzewc4p[15]);
  wire[64-1:0] dhroqc1noi7tp8jgubh =  {64{z03_wl6z1na1ebppos | dl1k34qvje99ofpsjzadtq61}} & {
     ({1'b0,{15{ktbf6dfpqw7ullwvs0}}} | ({16{duhacqzewc4p[76] & duhacqzewc4p[75]}} & (~duhacqzewc4p[75:60])) | ({16{(~duhacqzewc4p[76]) & (~duhacqzewc4p[75])}} & duhacqzewc4p[75:60])),
     ({1'b0,{15{ryfbr1ol3w448dqtaictsz}}} | ({16{duhacqzewc4p[56] & duhacqzewc4p[55]}} & (~duhacqzewc4p[55:40])) | ({16{(~duhacqzewc4p[56]) & (~duhacqzewc4p[55])}} & duhacqzewc4p[55:40])), 
     ({1'b0,{15{o_j64jm_72wyhefzn9g7}}} | ({16{duhacqzewc4p[36] & duhacqzewc4p[35]}} & (~duhacqzewc4p[35:20])) | ({16{(~duhacqzewc4p[36]) & (~duhacqzewc4p[35])}} & duhacqzewc4p[35:20])),
     ({1'b0,{15{iktahd9pfcstthpcp_dnu}}} | ({16{duhacqzewc4p[16] & duhacqzewc4p[15]}} & (~duhacqzewc4p[15:0 ])) | ({16{(~duhacqzewc4p[16]) & (~duhacqzewc4p[15])}} & duhacqzewc4p[15:0 ]))};
  
  wire ov3_mcecffyeq92798y4 = (z03_wl6z1na1ebppos | dl1k34qvje99ofpsjzadtq61) & (
                ktbf6dfpqw7ullwvs0 | ryfbr1ol3w448dqtaictsz |
                o_j64jm_72wyhefzn9g7 | iktahd9pfcstthpcp_dnu
              );
  wire jz527i0yzwr4knc0kjuzz = 1'b0;
  wire dpbsk_b28bd84i234    =  ov3_mcecffyeq92798y4 | jz527i0yzwr4knc0kjuzz;

  
  
  wire gadt0zg6g1b97hecbm_ = (ck6o6flrt == 4'b0111) & (pxscquhi78 == 3'b001);
  wire[64-1:0] jx3v45j8o22kd = {64{gadt0zg6g1b97hecbm_}} & {
                             ({16{duhacqzewc4p[76]}} | duhacqzewc4p[75:60]), ({16{~(duhacqzewc4p[56])}} & duhacqzewc4p[55:40]), 
                             ({16{duhacqzewc4p[36]}} | duhacqzewc4p[35:20]), ({16{~(duhacqzewc4p[16])}} & duhacqzewc4p[15:0 ])
                          };
  wire vztdr9wa4oxcxe = gadt0zg6g1b97hecbm_ & (
                            duhacqzewc4p[76] | duhacqzewc4p[56] |
                            duhacqzewc4p[36] | duhacqzewc4p[16]
                          );

  
  
  wire lrg2t_uhh4me2ix3ii = (ck6o6flrt == 4'b1000) & (pxscquhi78 == 3'b001);
  wire[64-1:0] s562ayhfwthes5 = {64{lrg2t_uhh4me2ix3ii}} & { 
                             ({16{~(duhacqzewc4p[76])}} & duhacqzewc4p[75:60]), ({16{duhacqzewc4p[56]}} | duhacqzewc4p[55:40]),    
                             ({16{~(duhacqzewc4p[36])}} & duhacqzewc4p[35:20]), ({16{duhacqzewc4p[16]}} | duhacqzewc4p[15:0 ])
                          };  
  wire i8trjvyz72w = lrg2t_uhh4me2ix3ii & (                             
                            duhacqzewc4p[76] | duhacqzewc4p[56] |
                            duhacqzewc4p[36] | duhacqzewc4p[16]
                          );

  
  
  wire mcr2vfu0w3r3d8spnrl = (ck6o6flrt == 4'b0111) & (pxscquhi78 == 3'b110);
  wire[64-1:0] dfwr3dn_zawt30y = {64{mcr2vfu0w3r3d8spnrl}} & {
                             ({32{duhacqzewc4p[72]}} | duhacqzewc4p[71:40]),  
                             ({32{~(duhacqzewc4p[32])}} & duhacqzewc4p[31:0 ])
                          };
  wire f9mkw5ch2tbrj = mcr2vfu0w3r3d8spnrl & (
                            duhacqzewc4p[72] | 
                            duhacqzewc4p[32]  
                          );

  
  wire puuohaeslh1xpmy = (ck6o6flrt == 4'b1000) & (pxscquhi78 == 3'b110);
  wire[64-1:0] qhu3idrzkhfjzcw0e1h = {64{puuohaeslh1xpmy}} & { 
                             ({32{~(duhacqzewc4p[72])}} & duhacqzewc4p[71:40]),
                             ({32{duhacqzewc4p[32]}} | duhacqzewc4p[31: 0])  
                          };  
  wire h8tkfq512i86f5 = puuohaeslh1xpmy & (                             
                            duhacqzewc4p[72] | 
                            duhacqzewc4p[32]  
                          );

  
  
  
  
  
  wire o8u0ps1oxtnnwr8u8h = (ck6o6flrt == 4'b0010) & (pxscquhi78 == 3'b010) & lvhs9fkt_6d9;
  wire bad1at5cv0jn3xqzjx = ~duhacqzewc4p[32] &  (|duhacqzewc4p[31:15]); 
  wire o4pl0c_i553kg5_as0tlgk =  duhacqzewc4p[32] & ~(&duhacqzewc4p[31:15]); 
  wire[64-1:0] i4l0fq5q10bfzz9h = {64{o8u0ps1oxtnnwr8u8h}} & (
          ({ {64-15{1'b0}}, {15{bad1at5cv0jn3xqzjx}} }) 
         |({64{o4pl0c_i553kg5_as0tlgk}} & {{64-32{1'b1}},32'hffff8000}) 
         |({64{~bad1at5cv0jn3xqzjx & ~o4pl0c_i553kg5_as0tlgk}} & {{64-16{duhacqzewc4p[32]}},duhacqzewc4p[15:0]} )
         );




  wire h4idev9r835k7 = o8u0ps1oxtnnwr8u8h & (bad1at5cv0jn3xqzjx | o4pl0c_i553kg5_as0tlgk);

  
  wire q0ycwm826m2lrqr = (ck6o6flrt == 4'b0011) & (pxscquhi78 == 3'b010) & lvhs9fkt_6d9;
  wire jtrfd3ax9bqg1my9hs = ~duhacqzewc4p[32] & (|duhacqzewc4p[31:16]); 
  wire gsag77aet1oqjbgz =  duhacqzewc4p[32]; 
  wire[64-1:0] kx4l6ahx1wqd388 = {64{q0ycwm826m2lrqr}} & (
           ({ {64-16{1'b0}}, {16{jtrfd3ax9bqg1my9hs}} }) 
         | ({64{~jtrfd3ax9bqg1my9hs & ~gsag77aet1oqjbgz}} & {{64-16{duhacqzewc4p[32]}}, duhacqzewc4p[15:0]}));
  wire kiasjfektpu75789v = q0ycwm826m2lrqr & (jtrfd3ax9bqg1my9hs | gsag77aet1oqjbgz);

  
  wire q2nmfs8kb443fb9 = (ck6o6flrt == 4'b0011) & (pxscquhi78 == 3'b010) & ~lvhs9fkt_6d9;
  wire rjo1wu6ovecxpkynwhq = (|duhacqzewc4p[32:16]); 
  wire[64-1:0] fyucfk2732ngvllwz39 = {64{q2nmfs8kb443fb9}} &
          (({ {64-16{1'b0}},{16{rjo1wu6ovecxpkynwhq}}}) | ({64{~rjo1wu6ovecxpkynwhq}} & {{64-16{1'b0}}, duhacqzewc4p[15:0]}));
  wire efuzf0v9fiwcx8 = q2nmfs8kb443fb9 & (rjo1wu6ovecxpkynwhq);

  

  wire vzv9psgyd30qoe = (ck6o6flrt == 4'b0100) & (pxscquhi78 == 3'b010) & lvhs9fkt_6d9;
  wire lx4ithjn8sb8_ez9al7ive8 = ~duhacqzewc4p[32] &  duhacqzewc4p[31]; 
  wire bblw_vqnu7n6p_h9wc2mx1ph =  duhacqzewc4p[32] & ~duhacqzewc4p[31]; 
  wire[64-1:0] o3uxjktahobimz2cuq = {64{vzv9psgyd30qoe}} & (
            ({ {64-31{1'b0}},{31{lx4ithjn8sb8_ez9al7ive8}} }) 
          | ({64{bblw_vqnu7n6p_h9wc2mx1ph}} & {{64-32{1'b1}}, 32'h80000000}) 
          | ({64{~lx4ithjn8sb8_ez9al7ive8 & ~bblw_vqnu7n6p_h9wc2mx1ph}} & {{64-32{duhacqzewc4p[32]}}, duhacqzewc4p[31:0]}));
  wire vxgf74c9k4wav = vzv9psgyd30qoe & (lx4ithjn8sb8_ez9al7ive8 | bblw_vqnu7n6p_h9wc2mx1ph);

  
  wire x30664wf1w8_fy9mpu = (ck6o6flrt == 4'b0101) & (pxscquhi78 == 3'b010) & lvhs9fkt_6d9;
  wire[64-1:0] fs7dqhxyc73iyp1 = {64{x30664wf1w8_fy9mpu}} & ({64{~duhacqzewc4p[32]}} & {{64-32{duhacqzewc4p[32]}}, duhacqzewc4p[31:0]});
  wire uldvolfjsstpft = x30664wf1w8_fy9mpu & (duhacqzewc4p[32]);

  
  wire hk5jt97w1cnrj8h1 = (ck6o6flrt == 4'b0101) & (pxscquhi78 == 3'b010) & ~lvhs9fkt_6d9;
  wire[64-1:0] ha0257hzj9t3v6jb = {64{hk5jt97w1cnrj8h1}} & {
           {64-32{1'b0}},
          (({32{duhacqzewc4p[32]}}) | ({32{~duhacqzewc4p[32]}} & duhacqzewc4p[31:0]))
          };
  wire wa6q6g2aaaon138i = hk5jt97w1cnrj8h1 & duhacqzewc4p[32];

  
  wire ya6g1fxkdo56ik = (ck6o6flrt == 4'b0100) & (pxscquhi78 == 3'b110) & lvhs9fkt_6d9;
  wire gxgjxbqnlk01_t0dzqx7id2v = ~duhacqzewc4p[72] &  duhacqzewc4p[71]; 
  wire t25wd_n4i31atn8pxcyn31jge3bj =  duhacqzewc4p[72] & ~duhacqzewc4p[71]; 
  wire cm5lyy2a6zojbs1y_cswigf90li = ~duhacqzewc4p[32] &  duhacqzewc4p[31]; 
  wire pbe2_4q8yoh_1q9zcw1kt8vh =  duhacqzewc4p[32] & ~duhacqzewc4p[31]; 
  wire[64-1:0] i0thro2gq50h4y = {64{ya6g1fxkdo56ik}} & {
              (({ 1'b0, {31{gxgjxbqnlk01_t0dzqx7id2v}} }) | ({32{t25wd_n4i31atn8pxcyn31jge3bj}} & 32'h80000000) 
            | ({32{~gxgjxbqnlk01_t0dzqx7id2v & ~t25wd_n4i31atn8pxcyn31jge3bj}} & duhacqzewc4p[71:40])), 
              (({ 1'b0, {31{cm5lyy2a6zojbs1y_cswigf90li}} }) | ({32{pbe2_4q8yoh_1q9zcw1kt8vh}} & 32'h80000000) 
            | ({32{~cm5lyy2a6zojbs1y_cswigf90li & ~pbe2_4q8yoh_1q9zcw1kt8vh}} & duhacqzewc4p[31: 0]))} ;
  wire sezz2frrpika9l8 = ya6g1fxkdo56ik & (gxgjxbqnlk01_t0dzqx7id2v | t25wd_n4i31atn8pxcyn31jge3bj | cm5lyy2a6zojbs1y_cswigf90li | pbe2_4q8yoh_1q9zcw1kt8vh);

  
  wire ux37hndoelyb7qgr_ = (ck6o6flrt == 4'b0101) & (pxscquhi78 == 3'b110) & lvhs9fkt_6d9;
  wire w6t3hserxetpk =  ~duhacqzewc4p[72]; 
  wire jxqr7cnincrvczzn4 =  ~duhacqzewc4p[32]; 
  wire[64-1:0] iksbn3wj9ty037ghle = {64{ux37hndoelyb7qgr_}} & {
              ({32{w6t3hserxetpk}} & duhacqzewc4p[71:40]), 
              ({32{jxqr7cnincrvczzn4}} & duhacqzewc4p[31: 0])} ;
  wire gg_e00der0k6v3zhpi = ux37hndoelyb7qgr_ & (~w6t3hserxetpk | ~jxqr7cnincrvczzn4);

  
  wire a24cdlzq0tq0u3g6 = (ck6o6flrt == 4'b0101) & (pxscquhi78 == 3'b110) & ~lvhs9fkt_6d9;
  wire onm_08po1ggfm2ljby_qyky = duhacqzewc4p[72]; 
  wire yfr6_6n84509z2l5h4dm2cx = duhacqzewc4p[32]; 
  wire[64-1:0] unmgl0ftbvgshye0 = {64{a24cdlzq0tq0u3g6}} & {
              ({32{onm_08po1ggfm2ljby_qyky}} | ({32{~onm_08po1ggfm2ljby_qyky}} & duhacqzewc4p[71:40])), 
              ({32{yfr6_6n84509z2l5h4dm2cx}} | ({32{~yfr6_6n84509z2l5h4dm2cx}} & duhacqzewc4p[31: 0]))} ;
  wire f_tovd0gdluco1rissz = a24cdlzq0tq0u3g6 & (onm_08po1ggfm2ljby_qyky | yfr6_6n84509z2l5h4dm2cx);






  
  wire rj2hmfjonjn6cac7r5q = (ck6o6flrt == 4'b0110) & (pxscquhi78 == 3'b010);
  wire gkj167gqqh8grv1hc = duhacqzewc4p[32] & (~duhacqzewc4p[31]);
  wire[31:0] mc9pvantv2ppcyam = {32{rj2hmfjonjn6cac7r5q}} &
       {{1'b0,{31{gkj167gqqh8grv1hc}}} | ({32{duhacqzewc4p[32] & duhacqzewc4p[31]}} & (~duhacqzewc4p[31:0 ])) | ({32{(~duhacqzewc4p[32]) & (~duhacqzewc4p[31])}} & duhacqzewc4p[31:0 ])};
  wire fr3icsm_kbjc = rj2hmfjonjn6cac7r5q & (gkj167gqqh8grv1hc);

  
  wire flrr6m298i_cx37q5_j2 = (ck6o6flrt == 4'b0110) & (pxscquhi78 == 3'b110);
  wire r9vm9lym204uz6sda48 = duhacqzewc4p[72] & (~duhacqzewc4p[71]);
  wire ics21s5hej6th338r0 = duhacqzewc4p[32] & (~duhacqzewc4p[31]);
  wire[63:0] ztd3zuipbi5y_eb8 = {64{flrr6m298i_cx37q5_j2}} & {
    ({1'b0,{31{r9vm9lym204uz6sda48}}}) | ({32{duhacqzewc4p[72] & duhacqzewc4p[71]}} & (~duhacqzewc4p[71:40])) | ({32{(~duhacqzewc4p[72]) & (~duhacqzewc4p[71])}} & duhacqzewc4p[71:40]),
    ({1'b0,{31{ics21s5hej6th338r0}}}) | ({32{duhacqzewc4p[32] & duhacqzewc4p[31]}} & (~duhacqzewc4p[31:0 ])) | ({32{(~duhacqzewc4p[32]) & (~duhacqzewc4p[31])}} & duhacqzewc4p[31:0 ])
    };
  wire gqe3pghk01419 = flrr6m298i_cx37q5_j2 & (ics21s5hej6th338r0 | r9vm9lym204uz6sda48);





  
  wire zxl27nzmujz1bwez = (ck6o6flrt == 4'b1001) & (pxscquhi78 == 3'b011) & lvhs9fkt_6d9;
  wire s63qmwsevfy071iudvvi0 = ~duhacqzewc4p[64] &  duhacqzewc4p[63]; 
  wire tzf8pfo3f5nctbpgrbp =  duhacqzewc4p[64] & ~duhacqzewc4p[63]; 
  wire[64-1:0] m_5k9yxib3e9ma019j = {64{zxl27nzmujz1bwez}} &
           (({64{s63qmwsevfy071iudvvi0}} & {32'h7fffffff,32'hffffffff}) 
          | ({64{tzf8pfo3f5nctbpgrbp}} & {1'b1,{64-1{1'b0}}}) 
          | ({64{(~s63qmwsevfy071iudvvi0 & ~tzf8pfo3f5nctbpgrbp)}} & duhacqzewc4p[64-1:0]));



  wire srcojqjcmmadp2u = zxl27nzmujz1bwez & (s63qmwsevfy071iudvvi0 | tzf8pfo3f5nctbpgrbp);

  
  wire hepglnwgst84t7c0g = (ck6o6flrt == 4'b1010) & (pxscquhi78 == 3'b011) & lvhs9fkt_6d9;
  wire[64-1:0] tlozsyh0dxincxc71ch = {64{hepglnwgst84t7c0g}} &
           (({64{duhacqzewc4p[64]}} & {64{1'b0}}) 
          | ({64{~duhacqzewc4p[64]}} & duhacqzewc4p[64-1:0]));
  wire xbnlp_yi87losqbct = hepglnwgst84t7c0g & (duhacqzewc4p[64]);

  
  wire euysszeuwmncykamhy = (ck6o6flrt == 4'b1010) & (pxscquhi78 == 3'b011) & ~lvhs9fkt_6d9;
  wire[64-1:0] ku2wkk7jsne7e8tja_9 = {64{euysszeuwmncykamhy}} &
           (({64{duhacqzewc4p[64]}} & {64{1'b1}}) 
          | ({64{~duhacqzewc4p[64]}} & duhacqzewc4p[64-1:0]));
  wire q0mfxbs3petvezf = euysszeuwmncykamhy & (duhacqzewc4p[64]);


  wire[64-1:0] ugh99u1va5po = 
          ({64{t9r50zrh89s7ztk   }}    &  {uxo500z5tj5fa1j})  
         |({64{khqzwdn7t8_cfub9p | b6hhq101tety5ku7 }}    
                                             &  {utgqzem07taxie245})  
         |({64{otvnx5pkt5aw    }}    &  {mta9g3ta_8x7b3tqa}) 
         |({64{megmtexkcejn7j4t |  v8g190egj7fkzr036wsol8d}}  
                                             &  {qfnxty3b3r0wv5b_}) 
         |({64{ush3kg4qf4rchvxt | q8cq6922962cszd1w1ibpy}}   
                                             &  {i8hs0nk1rk1897rxqa}) 
         |({64{rtvs3qjdc4jbzne }}    &  {h59gmpawefdlc7erk9nq}) 
         |({64{u1xa8v9g_87fspma  }}    &  {ek7dk29izkdtor}) 
         |({64{z03_wl6z1na1ebppos |  dl1k34qvje99ofpsjzadtq61}}
                                             &  {dhroqc1noi7tp8jgubh}) 
         |({64{gadt0zg6g1b97hecbm_ }}    &  {jx3v45j8o22kd})
         |({64{lrg2t_uhh4me2ix3ii }}    &  {s562ayhfwthes5}) 
         |({64{mcr2vfu0w3r3d8spnrl }}    &  {dfwr3dn_zawt30y}) 
         |({64{puuohaeslh1xpmy }}    &  {qhu3idrzkhfjzcw0e1h})
         |({64{o8u0ps1oxtnnwr8u8h }}      &  {i4l0fq5q10bfzz9h})                         
         |({64{q0ycwm826m2lrqr }}      &  {kx4l6ahx1wqd388})                         
         |({64{q2nmfs8kb443fb9 }}     &  {fyucfk2732ngvllwz39})                         
         |({64{vzv9psgyd30qoe }}      &  {o3uxjktahobimz2cuq})                         
         |({64{x30664wf1w8_fy9mpu }}      &  {fs7dqhxyc73iyp1})                         
         |({64{hk5jt97w1cnrj8h1 }}     &  {ha0257hzj9t3v6jb})                         
         |({64{rj2hmfjonjn6cac7r5q }}    &  {mc9pvantv2ppcyam})                         
         |({64{ya6g1fxkdo56ik }}     &  {i0thro2gq50h4y})                         
         |({64{ux37hndoelyb7qgr_ }}     &  {iksbn3wj9ty037ghle})                         
         |({64{a24cdlzq0tq0u3g6 }}    &  {unmgl0ftbvgshye0}) 
         |({64{zxl27nzmujz1bwez }}     &  m_5k9yxib3e9ma019j)                         
         |({64{hepglnwgst84t7c0g }}     &  tlozsyh0dxincxc71ch)                         
         |({64{euysszeuwmncykamhy}}     &  ku2wkk7jsne7e8tja_9)                         
         |({64{flrr6m298i_cx37q5_j2 }}  &  {ztd3zuipbi5y_eb8})                         
         ;

  wire a2u9_cwjyyq = sy1xledv0xcnby3   
              | w3wxllzvry4npxh  
              | g1j_85l4zzhsb  
              | z8_ag3wbvbhcdp 
              | mqo5q_91fbwq6p3r
              | e6tk2oatobnknne 
              | suunz_obigrbmg8
              | dpbsk_b28bd84i234
              | vztdr9wa4oxcxe  
              | i8trjvyz72w  
              | f9mkw5ch2tbrj  
              | h8tkfq512i86f5  
              | h4idev9r835k7
              | kiasjfektpu75789v
              | efuzf0v9fiwcx8 
              | vxgf74c9k4wav
              | uldvolfjsstpft
              | wa6q6g2aaaon138i 
              | sezz2frrpika9l8
              | gg_e00der0k6v3zhpi
              | f_tovd0gdluco1rissz 
              | fr3icsm_kbjc 
              | srcojqjcmmadp2u 
              | xbnlp_yi87losqbct 
              | q0mfxbs3petvezf
              | gqe3pghk01419 
                ;

            
            
            
assign vvoozaywykiwmels = ugh99u1va5po;
assign m50l82p03g15y_ehxthx1 = {64{1'b0}};
assign hsvg_y2njolj1bl    = a2u9_cwjyyq ;

endmodule                                      
                                               






















module uq9oowb3c0mb0eda15rcw5 # (
  parameter ctu6y0yy1_ = 5   
) (
  input                   f218verzay1lfg_t73r7h    ,      
  input                   wvyn3jdt7m5qk570c1zta     ,      
  input  [64-1:0] v2k5ixyb1cco74jghjt          ,      
  input  [ctu6y0yy1_-1:0]      mhres_bf8ykyi80s          ,      
  output [64-1:0] jhqv9u46f4ilao8a7rqc    ,      
  output [64-1:0] en2fwj8b2lksbcaz8_f            

  );

wire j4qv5sod = f218verzay1lfg_t73r7h | f218verzay1lfg_t73r7h;

wire [64-1:0] svtp9g_orl2 = v2k5ixyb1cco74jghjt;
wire [ctu6y0yy1_-1:0]      ovco_g1rr8cl = mhres_bf8ykyi80s;

wire [64-1:0] eaks5rrtzx4;
wire [ctu6y0yy1_-1:0]      qkr7a25rdze;

wire [64-1:0] pw0intormjs1h2x2_69;
i6_4g5fspqlv1svn #(64) zq7zotg5pn5z656ukciuy(svtp9g_orl2, pw0intormjs1h2x2_69);



assign eaks5rrtzx4 =   ({64{f218verzay1lfg_t73r7h}} & pw0intormjs1h2x2_69)
                     | ({64{wvyn3jdt7m5qk570c1zta }} & svtp9g_orl2   )
                     ;

assign qkr7a25rdze = ovco_g1rr8cl;

wire [64-1:0] cvnvrq3lozc;
assign cvnvrq3lozc = (eaks5rrtzx4 << qkr7a25rdze);

assign en2fwj8b2lksbcaz8_f = cvnvrq3lozc;

i6_4g5fspqlv1svn #(64) yt03iszk9clnc02oa6q0m1(cvnvrq3lozc, jhqv9u46f4ilao8a7rqc);

endmodule









































































module aiw2b4qk64vf3344ezyf # (
  parameter ctu6y0yy1_ = 5 
)
(

  
  
  
  



  input  [64-1:0] amgi_rqhtd007,
  input  [64-1:0] otn5ycgat1c9s1a,
  input  [64-1:0] g7tawq8tp6,
  input  [105-1:0] xlkm1ikvsatc2,
  
  
  
  
  output g36_kozc0w4bjtnf,
  output [80-1:0] ileuocpyluq,
  output [80-1:0] yiexcriz0ufmy,
  input  [80-1:0] e231c11ou7ube_b,
  
  
  
  
  output tppbcuxfcn35ghrqja5,
  output iv4pxzd85kko8e8twyro,
  output [64-1:0] ixlv8n_7cgrz2,
  output [64-1:0] gxtsmhtras93dt4g11,
  output [ctu6y0yy1_-1:0]      i8fcutzmv9eer,
  input  [64-1:0] kth4tafeif3978quzt,
  input  [64-1:0] eltrj3g68c3h11e7zli4x0t9,
  input  [64-1:0] u9d99u2san4lbuhbb,
  input  [64-1:0] xlxi2zedzir0xwdjxt,

  
  
  


    
  output [64-1:0] nb3w1rq_ny95rvrt,
  output [64-1:0] dkojj6fim0nxg4jvyafk,
  output vjkz8n6i44pc7o

  );





wire ut6ov1    = xlkm1ikvsatc2[11:11]; 
wire t_5k8fg   = xlkm1ikvsatc2[12:12];
wire dn4ly52z   = xlkm1ikvsatc2[13:13];
wire sz2kkvytoq  = xlkm1ikvsatc2[14:14];
wire uhoire    = xlkm1ikvsatc2[15:15];
wire edo25py4   = xlkm1ikvsatc2[16:16];
wire gnzgoy2_   = xlkm1ikvsatc2[17:17];
wire m2_gkl2  = xlkm1ikvsatc2[18:18];
wire touyo1q    = xlkm1ikvsatc2[19:19];
wire fy8t8148dy   = xlkm1ikvsatc2[20:20];
wire u_l_if   = xlkm1ikvsatc2[21:21];
wire jp3kdt1oe  = xlkm1ikvsatc2[22:22];
wire qchqfra5  = xlkm1ikvsatc2[23:23];
wire ru_hz78 = xlkm1ikvsatc2[24];
wire jnsck9jg4bp = xlkm1ikvsatc2[25:25];
wire l5ydun7   = xlkm1ikvsatc2[26:26];
wire gqnr2s  = xlkm1ikvsatc2[27:27];
wire k_0a102szv0  = xlkm1ikvsatc2[28:28];
wire z09vlclwa = xlkm1ikvsatc2[29:29];
wire uvj5g7_5   = xlkm1ikvsatc2[30:30];
wire u7_kdd  = xlkm1ikvsatc2[31:31];
wire uibivc  = xlkm1ikvsatc2[32:32];
wire mrjkej10vvl0 = xlkm1ikvsatc2[33:33];
wire unlte4n   = xlkm1ikvsatc2[34:34];
wire emldhbp2hfx  = xlkm1ikvsatc2[35:35];
wire m5423_2aw1a  = xlkm1ikvsatc2[36:36];
wire y5f5233zcx = xlkm1ikvsatc2[37:37];
wire f6zwhrtxxt = xlkm1ikvsatc2[38:38];
wire b8qm5m9c4mc= xlkm1ikvsatc2[39];
wire cd1wg_ulmyc9k= xlkm1ikvsatc2[40:40];
wire llv5rm1c   = xlkm1ikvsatc2[47:47];   
wire ruh95m  = xlkm1ikvsatc2[48:48];  
wire l8m8rnx5  = xlkm1ikvsatc2[49:49];  
wire ydvt8avgu = xlkm1ikvsatc2[50:50]; 
wire v5ra1fp   = xlkm1ikvsatc2[51:51];   
wire uu_lqkw  = xlkm1ikvsatc2[52:52];  
wire wnqcbf47  = xlkm1ikvsatc2[53:53];  
wire itn70c49go4u = xlkm1ikvsatc2[54:54]; 
wire k9mgr537   = xlkm1ikvsatc2[55:55];   
wire scsugeqe8ng  = xlkm1ikvsatc2[56:56];  
wire n6kqoj  = xlkm1ikvsatc2[57:57];  
wire j1yir7jdj3x = xlkm1ikvsatc2[58:58]; 
wire qcgre5j0h = xlkm1ikvsatc2[59:59]; 
wire c_fjxrw0ec27= xlkm1ikvsatc2[60:60];



wire go708t    = xlkm1ikvsatc2[41:41];
wire t3xtp_0m8b   = xlkm1ikvsatc2[42:42];
wire fpmfb946  = xlkm1ikvsatc2[43:43];
wire emx9j93ash5 = xlkm1ikvsatc2[44:44];
wire k24cqbg   = xlkm1ikvsatc2[45:45];
wire omx1o91b9q  = xlkm1ikvsatc2[46:46];
wire xy7f1zepm9  = xlkm1ikvsatc2[61:61]; 





wire [5:0] u_tbn73ael9rkr = xlkm1ikvsatc2[10:5];


wire xso8dz60n84ql  = t_5k8fg | sz2kkvytoq | edo25py4 | m2_gkl2 | fy8t8148dy | jp3kdt1oe;
wire sapv8p6do3 = gqnr2s | z09vlclwa | u7_kdd | mrjkej10vvl0 | emldhbp2hfx | y5f5233zcx;
wire ih_s_3uvpxe = ruh95m | ydvt8avgu | uu_lqkw | itn70c49go4u | scsugeqe8ng | j1yir7jdj3x | xy7f1zepm9 | omx1o91b9q;
wire idcimwm2jndo = t3xtp_0m8b;
wire j948ulc40f    = ut6ov1 | dn4ly52z | uhoire | gnzgoy2_ | touyo1q | u_l_if;       
wire mexy1jr    = qchqfra5 | ru_hz78 | jnsck9jg4bp;                       
wire y8xct28c_1   = l5ydun7 | k_0a102szv0 | uvj5g7_5 | uibivc | unlte4n | m5423_2aw1a; 
wire s20eatde5   = f6zwhrtxxt | b8qm5m9c4mc | cd1wg_ulmyc9k;                    
wire lj1p441zbp   = llv5rm1c | l8m8rnx5 | v5ra1fp | wnqcbf47 | k9mgr537 | n6kqoj | k24cqbg; 
wire u22h_8pj   = qcgre5j0h | c_fjxrw0ec27 | fpmfb946 | emx9j93ash5;            

wire nzfb5yi7vj4f   = go708t;                                             
wire j3jhezvx6j   = 1'b0;                                             

wire [5:0] jp97gwmswq0z_wwwa = g7tawq8tp6[6] ? ((g7tawq8tp6[5:0] == 6'b0) ? 6'b111111 : ~g7tawq8tp6[5:0] + 1'b1) :
                              g7tawq8tp6[5:0];
wire [4:0] rh3ck_2qihzfryih3t2xm = g7tawq8tp6[5] ? ((g7tawq8tp6[4:0] == 5'b0) ? 5'b11111 : ~g7tawq8tp6[4:0] + 1'b1) :
                              g7tawq8tp6[4:0];
wire [3:0] nuwrfugjr0r9zj9ij53 = g7tawq8tp6[4] ? ((g7tawq8tp6[3:0] == 4'b0) ? 4'b1111 : ~g7tawq8tp6[3:0] + 1'b1) :
                              g7tawq8tp6[3:0];
wire [2:0] y8gc6wjxhqvx3xo3  = g7tawq8tp6[3] ? ((g7tawq8tp6[2:0] == 3'b0) ? 3'b111 : ~g7tawq8tp6[2:0] + 1'b1) :
                              g7tawq8tp6[2:0];

wire [5:0] ovco_g1rr8cl  = ({6{xso8dz60n84ql}}  & {3'b0, u_tbn73ael9rkr[2:0]})       |
                          ({6{sapv8p6do3}} & {2'b0, u_tbn73ael9rkr[3:0]})       |
                          ({6{ih_s_3uvpxe}} & {1'b0, u_tbn73ael9rkr[4:0]})       |
                          ({6{idcimwm2jndo}} & {      u_tbn73ael9rkr[5:0]})       |
                          ({6{j948ulc40f}}    & {3'b0, g7tawq8tp6[2:0]})         |
                          ({6{mexy1jr}}    & {3'b0, y8gc6wjxhqvx3xo3[2:0]})   |
                          ({6{y8xct28c_1}}   & {2'b0, g7tawq8tp6[3:0]})         |
                          ({6{s20eatde5}}   & {2'b0, nuwrfugjr0r9zj9ij53[3:0]})  |
                          ({6{lj1p441zbp}}   & {1'b0, g7tawq8tp6[4:0]})         |
                          ({6{u22h_8pj}}   & {1'b0, rh3ck_2qihzfryih3t2xm[4:0]})  |
                          ({6{nzfb5yi7vj4f}}   & {      g7tawq8tp6[5:0]})         |
                          ({6{j3jhezvx6j}}   & {      jp97gwmswq0z_wwwa[5:0]})  
                          ;



wire lun9svt1  = jp3kdt1oe | u_l_if | (qchqfra5 | ru_hz78  | jnsck9jg4bp) & ~g7tawq8tp6[3];
wire hr7jjg = y5f5233zcx | m5423_2aw1a | (f6zwhrtxxt | b8qm5m9c4mc | cd1wg_ulmyc9k) & ~g7tawq8tp6[4];
wire uayip3yhv = n6kqoj | j1yir7jdj3x | k24cqbg | omx1o91b9q | ((qcgre5j0h | c_fjxrw0ec27 | fpmfb946 | emx9j93ash5) & ~g7tawq8tp6[5]);
wire wxlzi41w2 = 1'b0;
wire n9mvknsj1brwzi9q3 = k24cqbg | omx1o91b9q | ((fpmfb946 | emx9j93ash5) & ~g7tawq8tp6[5]);
wire wj_jha74 = lun9svt1 | hr7jjg | uayip3yhv | wxlzi41w2;



wire v3eqx9ib0t  = sz2kkvytoq | dn4ly52z | (jnsck9jg4bp & g7tawq8tp6[3]);
wire g85zqyekqm  = m2_gkl2 | gnzgoy2_;
wire cfcw5xnn3i    = v3eqx9ib0t | g85zqyekqm;

wire q54kknz__om8vb = z09vlclwa | k_0a102szv0 | (cd1wg_ulmyc9k & g7tawq8tp6[4]);
wire f0d6_uwmzg = mrjkej10vvl0 | uibivc;
wire j_qce23   = q54kknz__om8vb | f0d6_uwmzg;
wire ahj4h_m1iaa_4x9qgb2fb = xy7f1zepm9 | (emx9j93ash5 & g7tawq8tp6[5]);
wire mxnjtosu3qfa8 = ydvt8avgu | l8m8rnx5 | xy7f1zepm9 | ((c_fjxrw0ec27 | emx9j93ash5) & g7tawq8tp6[5]);
wire tqok3m0mf8 = itn70c49go4u | wnqcbf47;
wire s864qhdj_vmxevu9  = (mxnjtosu3qfa8 & ~ahj4h_m1iaa_4x9qgb2fb) | tqok3m0mf8;
wire xd94m0cezzwq329zknc = ahj4h_m1iaa_4x9qgb2fb;
wire vu42s1b4t3   = mxnjtosu3qfa8 | tqok3m0mf8;
wire oc9vvnc_   = go708t | t3xtp_0m8b;
wire zr9gym5te   = v3eqx9ib0t | q54kknz__om8vb | mxnjtosu3qfa8 | oc9vvnc_;
wire jrdlxbxhql1v   = g85zqyekqm | f0d6_uwmzg | tqok3m0mf8;
wire wl451sp6zo  = cfcw5xnn3i | j_qce23 | vu42s1b4t3 | oc9vvnc_;



wire ok1mzu6  = edo25py4 | m2_gkl2 | uhoire | gnzgoy2_;
wire ru9kq5lf = u7_kdd | mrjkej10vvl0 | uvj5g7_5 | uibivc;
wire scyvyxdqtu4 = uu_lqkw | itn70c49go4u | v5ra1fp | wnqcbf47;
wire s6vixk9hul = 1'b0;
wire tdz9d9   = ok1mzu6 | ru9kq5lf | scyvyxdqtu4 | s6vixk9hul;


wire hc9cj_gw  = t_5k8fg | sz2kkvytoq | ut6ov1 | dn4ly52z | ((qchqfra5 | ru_hz78 | jnsck9jg4bp) & g7tawq8tp6[3]);
wire v_7x_ep_rfu = gqnr2s | z09vlclwa | l5ydun7 | k_0a102szv0 | ((f6zwhrtxxt | b8qm5m9c4mc | cd1wg_ulmyc9k) & g7tawq8tp6[4]);
wire esauilv2r = ruh95m | ydvt8avgu | llv5rm1c | l8m8rnx5 | xy7f1zepm9 | ((qcgre5j0h | c_fjxrw0ec27 | fpmfb946 | emx9j93ash5) & g7tawq8tp6[5]);
wire umogayoopjyhd4x7i = ((fpmfb946 | emx9j93ash5) & g7tawq8tp6[5]);
wire o8ydrzsk = go708t | t3xtp_0m8b;
wire jxe3dht   = hc9cj_gw | v_7x_ep_rfu | esauilv2r | o8ydrzsk;



wire wrer8n1vtx3  = fy8t8148dy | touyo1q | lun9svt1;

wire pajq0f4r = emldhbp2hfx | unlte4n | hr7jjg;

wire rh0exi5f = scsugeqe8ng | k9mgr537 | uayip3yhv;

wire w5rgrbjzguq = wxlzi41w2;
wire onsk4u1y9_e   = wrer8n1vtx3 | pajq0f4r | rh0exi5f | w5rgrbjzguq;

wire mwa0p8uyihgj = ok1mzu6 | hc9cj_gw | wrer8n1vtx3;
wire j7ilfx4t4s = ru9kq5lf | v_7x_ep_rfu | pajq0f4r;
wire jg1_gen5bgn7v4 = scyvyxdqtu4 | esauilv2r | rh0exi5f;
wire lz6cfqxwuxtx = s6vixk9hul | o8ydrzsk | w5rgrbjzguq;




wire [64-1:0] svtp9g_orl2   = amgi_rqhtd007;
wire [64-1:0] kyz24f5u7b6f42w_l = otn5ycgat1c9s1a;
assign tppbcuxfcn35ghrqja5 = jxe3dht | tdz9d9;
assign iv4pxzd85kko8e8twyro = onsk4u1y9_e;
assign ixlv8n_7cgrz2   = svtp9g_orl2;
assign gxtsmhtras93dt4g11 = kyz24f5u7b6f42w_l;
assign i8fcutzmv9eer   = ovco_g1rr8cl;

wire [64-1:0] m2ngrd23vsh;
wire [64-1:0] h6cvnvx_d3lnc1622y;
wire [64-1:0] zmfpztwuj1pzoik;
wire [64-1:0] bgh3d68j138h4ok_r7;
wire [64-1:0] ea1fw5akofqeu;
wire [64-1:0] ey9pskykeottfj5o;
wire [64-1:0] hvo606li;
wire [64-1:0] i7f4ir79mtemf6jp;

assign hvo606li             = (~(64'b0)) >> ovco_g1rr8cl;
assign i7f4ir79mtemf6jp[7:0]   = mwa0p8uyihgj ? hvo606li[63:56] : j7ilfx4t4s ? hvo606li[55:48] : jg1_gen5bgn7v4 ? hvo606li[39:32] : hvo606li[7:0];
assign i7f4ir79mtemf6jp[15:8]  = mwa0p8uyihgj ? hvo606li[63:56] : j7ilfx4t4s ? hvo606li[63:56] : jg1_gen5bgn7v4 ? hvo606li[47:40] : hvo606li[15:8];
assign i7f4ir79mtemf6jp[23:16] = mwa0p8uyihgj ? hvo606li[63:56] : j7ilfx4t4s ? hvo606li[55:48] : jg1_gen5bgn7v4 ? hvo606li[55:48] : hvo606li[23:16];
assign i7f4ir79mtemf6jp[31:24] = mwa0p8uyihgj ? hvo606li[63:56] : j7ilfx4t4s ? hvo606li[63:56] : jg1_gen5bgn7v4 ? hvo606li[63:56] : hvo606li[31:24];
assign i7f4ir79mtemf6jp[39:32] = mwa0p8uyihgj ? hvo606li[63:56] : j7ilfx4t4s ? hvo606li[55:48] : jg1_gen5bgn7v4 ? hvo606li[39:32] : hvo606li[39:32];
assign i7f4ir79mtemf6jp[47:40] = mwa0p8uyihgj ? hvo606li[63:56] : j7ilfx4t4s ? hvo606li[63:56] : jg1_gen5bgn7v4 ? hvo606li[47:40] : hvo606li[47:40];
assign i7f4ir79mtemf6jp[55:48] = mwa0p8uyihgj ? hvo606li[63:56] : j7ilfx4t4s ? hvo606li[55:48] : jg1_gen5bgn7v4 ? hvo606li[55:48] : hvo606li[55:48];
assign i7f4ir79mtemf6jp[63:56] = hvo606li[63:56];


wire [64-1:0] at20953pwlpl_sqg;
wire [64-1:0] zjnb75ihgiwibj67qc_;
assign at20953pwlpl_sqg[63:56] = {8{svtp9g_orl2[63]}};
assign at20953pwlpl_sqg[55:48] = mwa0p8uyihgj ? {8{svtp9g_orl2[55]}} : {8{svtp9g_orl2[63]}};
assign at20953pwlpl_sqg[47:40] = mwa0p8uyihgj ? {8{svtp9g_orl2[47]}} : j7ilfx4t4s ? {8{svtp9g_orl2[47]}} : {8{svtp9g_orl2[63]}};
assign at20953pwlpl_sqg[39:32] = mwa0p8uyihgj ? {8{svtp9g_orl2[39]}} : j7ilfx4t4s ? {8{svtp9g_orl2[47]}} : {8{svtp9g_orl2[63]}};
assign at20953pwlpl_sqg[31:24] = mwa0p8uyihgj ? {8{svtp9g_orl2[31]}} : j7ilfx4t4s ? {8{svtp9g_orl2[31]}} : jg1_gen5bgn7v4 ? {8{svtp9g_orl2[31]}} : {8{svtp9g_orl2[63]}};
assign at20953pwlpl_sqg[23:16] = mwa0p8uyihgj ? {8{svtp9g_orl2[23]}} : j7ilfx4t4s ? {8{svtp9g_orl2[31]}} : jg1_gen5bgn7v4 ? {8{svtp9g_orl2[31]}} : {8{svtp9g_orl2[63]}};
assign at20953pwlpl_sqg[15:8]  = mwa0p8uyihgj ? {8{svtp9g_orl2[15]}} : j7ilfx4t4s ? {8{svtp9g_orl2[15]}} : jg1_gen5bgn7v4 ? {8{svtp9g_orl2[31]}} : {8{svtp9g_orl2[63]}};
assign at20953pwlpl_sqg[7:0]   = mwa0p8uyihgj ? {8{svtp9g_orl2[7]}}  : j7ilfx4t4s ? {8{svtp9g_orl2[15]}} : jg1_gen5bgn7v4 ? {8{svtp9g_orl2[31]}} : {8{svtp9g_orl2[63]}}; 

assign zjnb75ihgiwibj67qc_ = 64'b0;






wire [64-1:0] p00v3vf3lxiy;
i6_4g5fspqlv1svn #(64) s66unx11bxb22phc(i7f4ir79mtemf6jp, p00v3vf3lxiy);

assign m2ngrd23vsh   = p00v3vf3lxiy & u9d99u2san4lbuhbb;
assign h6cvnvx_d3lnc1622y = p00v3vf3lxiy & xlxi2zedzir0xwdjxt;
assign ea1fw5akofqeu   = i7f4ir79mtemf6jp & kth4tafeif3978quzt;
assign ey9pskykeottfj5o = i7f4ir79mtemf6jp & eltrj3g68c3h11e7zli4x0t9;
assign zmfpztwuj1pzoik = ea1fw5akofqeu   | (at20953pwlpl_sqg   & (~i7f4ir79mtemf6jp));
wire [64-1:0] vt3rt5h12hv25u_6 = umogayoopjyhd4x7i ? {{32{zmfpztwuj1pzoik[31]}},zmfpztwuj1pzoik[31:0]} : zmfpztwuj1pzoik;

assign bgh3d68j138h4ok_r7 = ey9pskykeottfj5o | (zjnb75ihgiwibj67qc_ & (~i7f4ir79mtemf6jp));

wire j4qv5sod = jxe3dht | onsk4u1y9_e | tdz9d9; 

























































































localparam yk7 = 2;
localparam m0qq = 4;
localparam dk34z = 8;
wire [dk34z-1:0]         jxuls43sqwa;
wire [dk34z-1:0]         mj1ex47gsgf;
wire [dk34z-1:0]         g3x1whn96j2yq4;
wire [dk34z-1:0]         h12hgjnbituwg32d6;
wire [m0qq-1:0]         romko5ymdrfzzldtl;
wire [m0qq-1:0]         jlhtbk3erojleuz_d;
wire [m0qq-1:0]         fkjq_c0a1s83b0ab8;
wire [m0qq-1:0]         dnq81sp0s_88y0m3um;
wire [yk7-1:0]         zgg2kluk7qvo;
wire [yk7-1:0]         fz268jwgd_u7;


wire                  qup6ol8_fenrj;
wire                  km0c_ztzh4o9u0;
wire [64-1:0] wo3i0oqy69jb7   = {1'b0, i7f4ir79mtemf6jp[64-1:1]};
wire [64-1:0] w18mqmjcabw7wdfre   = ~wo3i0oqy69jb7;
wire [31:0]           xqbsjoxa9pziytk0   = {1'b0, i7f4ir79mtemf6jp[31:1]};
wire [31:0]           gve64r8imfbwkbk   = ~xqbsjoxa9pziytk0;
wire [15:0]           g6h7n2_hzn71eye   = {1'b0, i7f4ir79mtemf6jp[15:1]};
wire [15:0]           asd68nn3ya8thdexs0   = ~g6h7n2_hzn71eye;
wire [7:0]            nopz0l86oit1    = {1'b0, i7f4ir79mtemf6jp[7:1]};
wire [7:0]            seocst8b9xoupi0br    = ~nopz0l86oit1;

gr40tady98ryto733e #(
    .yk7(yk7),
    .m0qq(m0qq),
    .dk34z(dk34z)
) q0jzdszo0hdxo9q0sobo (
	.c5qrwj5sm0vc      ( svtp9g_orl2   ),     
	.of4kpekzgop8    ( kyz24f5u7b6f42w_l ),     
	.l59fhx3o23g9ig ( wo3i0oqy69jb7 ),     
	.p2v9igi9t66348 ( w18mqmjcabw7wdfre ),     
	.utwav9is_83yd6ng0 ( xqbsjoxa9pziytk0 ),     
	.sdmfqus_d4n5v3k ( gve64r8imfbwkbk ),     
	.ghpvhjxwavld6r6r0w2 ( g6h7n2_hzn71eye ),     
	.berx62p9_hc2bfcnyn0 ( asd68nn3ya8thdexs0 ),     
	.ky3ucnc3e8n4c_iz  ( nopz0l86oit1  ),     
	.v98eqhdqs8d1wk_qf2  ( seocst8b9xoupi0br  ),     
	.p2tb25qpyet2a_c    ( qup6ol8_fenrj  ),     
	.wms1mxki5gyfyc    ( km0c_ztzh4o9u0  ),     
	.tkuhwm5tyjr    ( zgg2kluk7qvo  ),     
	.rg1trb_7w92    ( fz268jwgd_u7  ),     
	.a1bp0x22t5vu4q    ( romko5ymdrfzzldtl  ),     
	.rgxbhxlvt61yfzn    ( jlhtbk3erojleuz_d  ),     
	.jpltrmmj8jw4lh_  ( fkjq_c0a1s83b0ab8),     
	.gs2s9lvzd_phhnv  ( dnq81sp0s_88y0m3um),     
	.j694o6frj_680_g     ( jxuls43sqwa   ),     
	.n2nedhasxux7buh     ( mj1ex47gsgf   ),     
	.fnv_7okzmo6y4ne85   ( g3x1whn96j2yq4 ),     
	.u_frczxmkmo88ujnp   ( h12hgjnbituwg32d6 )      
);


genvar i;
wire [64-1:0] p3kyq91_n;
wire [64-1:0] v4o5lfhyjaa;










generate 

for(i=0;i<dk34z;i=i+1) begin: kq32sucrnd_m
    assign p3kyq91_n[i*8+7:i*8]   = jxuls43sqwa[i] ? 8'h7f : mj1ex47gsgf[i] ? 8'h80 : m2ngrd23vsh[i*8+7:i*8];
    assign v4o5lfhyjaa[i*8+7:i*8] = g3x1whn96j2yq4[i] ? 8'h7f : h12hgjnbituwg32d6[i] ? 8'h80 : h6cvnvx_d3lnc1622y[i*8+7:i*8];
end

endgenerate

wire [64-1:0] dsbgxzsgdrjcjt;
wire [64-1:0] szhlof75yeu3;





generate 

for(i=0;i<m0qq;i=i+1) begin: wcwb1wp5fxxpxr5
    assign dsbgxzsgdrjcjt[i*16+15:i*16]   = romko5ymdrfzzldtl[i] ? 16'h7fff : jlhtbk3erojleuz_d[i] ? 16'h8000 : m2ngrd23vsh[i*16+15:i*16];
    assign szhlof75yeu3[i*16+15:i*16] = fkjq_c0a1s83b0ab8[i] ? 16'h7fff : dnq81sp0s_88y0m3um[i] ? 16'h8000 : h6cvnvx_d3lnc1622y[i*16+15:i*16];
end

endgenerate

wire [64-1:0] lhuukyau2oh;


generate 

for(i=0;i<yk7;i=i+1) begin: zu9h8b9119xca
    assign lhuukyau2oh[i*32+31:i*32]   = zgg2kluk7qvo[i] ? 32'h7fffffff : fz268jwgd_u7[i] ? 32'h80000000 : m2ngrd23vsh[i*32+31:i*32];
end

endgenerate






wire [64-1:0] ugh99u1va5po;
wire [64-1:0] kfxwyv6mbdgh;
assign ugh99u1va5po          = lun9svt1 ? p3kyq91_n :
                          hr7jjg ? dsbgxzsgdrjcjt :
                          
                          n9mvknsj1brwzi9q3 ? {{32{lhuukyau2oh[31]}},lhuukyau2oh[31:0]} :
                          lhuukyau2oh;

assign kfxwyv6mbdgh        = lun9svt1 ? v4o5lfhyjaa :
                          szhlof75yeu3;






wire [64:0]   wtfp4gxo7pevz2vwfc7;  
wire [64-1:0] pxpgx5vsyhow3ewy; 

wire [64-1:0] olho7eiv2f6;  



i6_4g5fspqlv1svn #(64) nj6ph6h2wz9g_dimed(hvo606li, pxpgx5vsyhow3ewy);

assign wtfp4gxo7pevz2vwfc7 = {1'b1, pxpgx5vsyhow3ewy};


generate 
	for(i=0; i<64; i=i+1) begin: jshecjs0wfglrht2s1

		assign olho7eiv2f6[i] = (~wtfp4gxo7pevz2vwfc7[i] & wtfp4gxo7pevz2vwfc7[i+1]);
	end
endgenerate





wire [dk34z-1:0] b895nyu5cwm2r;





generate 
for(i=0;i<dk34z;i=i+1) begin: a6kajbrkldyp_toc7db2
    assign b895nyu5cwm2r[i]   = |(svtp9g_orl2[i*8+7:i*8] & olho7eiv2f6[7:0]);
end
endgenerate


wire [m0qq-1:0] z1_x22aynlw60_;





generate 
for(i=0;i<m0qq;i=i+1) begin: kc6qdc5599100y24vlgu2r
    if(i==0) begin: mx6vg27fyr2tkgquyltsu
        assign z1_x22aynlw60_[i]   = (|(svtp9g_orl2[15:8] & olho7eiv2f6[15:8])) | b895nyu5cwm2r[0];
    end
    else begin : iu_rl21c17vnxsn25lmrueb1_o
        assign z1_x22aynlw60_[i]   = |(svtp9g_orl2[i*16+15:i*16] & olho7eiv2f6[15:0]);
    end
end
endgenerate


wire [yk7-1:0] jbq3yelms9pzd4g8v;



generate 
for(i=0;i<yk7;i=i+1) begin: ady9y3x9uhrjm5vu8941
    if(i==0) begin: yahxg3uo3i0saphutiodvuyc
        assign jbq3yelms9pzd4g8v[i]   = (|(svtp9g_orl2[31:16] & olho7eiv2f6[31:16])) | z1_x22aynlw60_[0];
    end
    else begin : rhe103vdbxhzempcvw32bj4k1pv
        assign jbq3yelms9pzd4g8v[i]   = |(svtp9g_orl2[i*32+31:i*32] & olho7eiv2f6[31:0]);
    end
end
endgenerate

wire q4xu8jcd49_rpr;
assign q4xu8jcd49_rpr = (|(svtp9g_orl2[63:32] & olho7eiv2f6[63:32])) | jbq3yelms9pzd4g8v[0];   
























































assign ileuocpyluq =   ({80{v3eqx9ib0t }} & {1'b0, zmfpztwuj1pzoik[63], zmfpztwuj1pzoik[63:56], 1'b0, zmfpztwuj1pzoik[55], zmfpztwuj1pzoik[55:48],
                                                                 1'b0, zmfpztwuj1pzoik[47], zmfpztwuj1pzoik[47:40], 1'b0, zmfpztwuj1pzoik[39], zmfpztwuj1pzoik[39:32], 
                                                                 1'b0, zmfpztwuj1pzoik[31], zmfpztwuj1pzoik[31:24], 1'b0, zmfpztwuj1pzoik[23], zmfpztwuj1pzoik[23:16], 
                                                                 1'b0, zmfpztwuj1pzoik[15], zmfpztwuj1pzoik[15:8], 1'b0, zmfpztwuj1pzoik[7], zmfpztwuj1pzoik[7:0]})
                     | ({80{g85zqyekqm }} & {2'b0, ea1fw5akofqeu[63:56], 2'b0, ea1fw5akofqeu[55:48], 
                                                                 2'b0, ea1fw5akofqeu[47:40], 2'b0, ea1fw5akofqeu[39:32],
                                                                 2'b0, ea1fw5akofqeu[31:24], 2'b0, ea1fw5akofqeu[23:16],
                                                                 2'b0, ea1fw5akofqeu[15:8], 2'b0, ea1fw5akofqeu[7:0]})
                     | ({80{q54kknz__om8vb}} & {3'b0, zmfpztwuj1pzoik[63], zmfpztwuj1pzoik[63:48], 3'b0, zmfpztwuj1pzoik[47], zmfpztwuj1pzoik[47:32],
                                                                 3'b0, zmfpztwuj1pzoik[31], zmfpztwuj1pzoik[31:16], 3'b0, zmfpztwuj1pzoik[15], zmfpztwuj1pzoik[15:0]}) 
                     | ({80{f0d6_uwmzg}} & {4'b0, ea1fw5akofqeu[63:48], 4'b0, ea1fw5akofqeu[47:32],
                                                                 4'b0, ea1fw5akofqeu[31:16], 4'b0, ea1fw5akofqeu[15:0]})
                     | ({80{mxnjtosu3qfa8}} & {7'b0, zmfpztwuj1pzoik[63], zmfpztwuj1pzoik[63:32],
                                                                 7'b0, zmfpztwuj1pzoik[31], zmfpztwuj1pzoik[31:0]}) 
                     | ({80{tqok3m0mf8}} & {8'b0,ea1fw5akofqeu[63:32],
                                                                 8'b0,ea1fw5akofqeu[31:0]}) 
                     | ({80{oc9vvnc_  }} & {15'b0, zmfpztwuj1pzoik[63], zmfpztwuj1pzoik[63:0]}) 
                     ;

assign yiexcriz0ufmy =   ({80{v3eqx9ib0t }} & {9'b0, b895nyu5cwm2r[7], 9'b0, b895nyu5cwm2r[6], 9'b0, b895nyu5cwm2r[5], 9'b0, b895nyu5cwm2r[4],
                                                                 9'b0, b895nyu5cwm2r[3], 9'b0, b895nyu5cwm2r[2], 9'b0, b895nyu5cwm2r[1], 9'b0, b895nyu5cwm2r[0]})
                     | ({80{g85zqyekqm }} & {9'b0, b895nyu5cwm2r[7], 9'b0, b895nyu5cwm2r[6], 9'b0, b895nyu5cwm2r[5], 9'b0, b895nyu5cwm2r[4],
                                                                 9'b0, b895nyu5cwm2r[3], 9'b0, b895nyu5cwm2r[2], 9'b0, b895nyu5cwm2r[1], 9'b0, b895nyu5cwm2r[0]})
                     | ({80{q54kknz__om8vb}} & {19'b0, z1_x22aynlw60_[3], 19'b0, z1_x22aynlw60_[2],
                                                                 19'b0, z1_x22aynlw60_[1], 19'b0, z1_x22aynlw60_[0]})
                     | ({80{f0d6_uwmzg}} & {19'b0, z1_x22aynlw60_[3], 19'b0, z1_x22aynlw60_[2],
                                                                 19'b0, z1_x22aynlw60_[1], 19'b0, z1_x22aynlw60_[0]})
                     | ({80{tqok3m0mf8}} & {39'b0, jbq3yelms9pzd4g8v[1],39'b0, jbq3yelms9pzd4g8v[0]})
                     | ({80{mxnjtosu3qfa8}} & {39'b0, jbq3yelms9pzd4g8v[1],39'b0, jbq3yelms9pzd4g8v[0]})
                     | ({80{oc9vvnc_  }} & {79'b0,q4xu8jcd49_rpr})
                     ;

assign g36_kozc0w4bjtnf = wl451sp6zo;
wire [64-1:0] z8p8nm_hann2w4;

assign z8p8nm_hann2w4 =   ({64{cfcw5xnn3i         }} & {e231c11ou7ube_b[77:70], e231c11ou7ube_b[67:60], e231c11ou7ube_b[57:50], e231c11ou7ube_b[47:40],e231c11ou7ube_b[37:30], e231c11ou7ube_b[27:20], e231c11ou7ube_b[17:10], e231c11ou7ube_b[7:0]})
                   | ({64{j_qce23        }} & {e231c11ou7ube_b[75:60], e231c11ou7ube_b[55:40], e231c11ou7ube_b[35:20], e231c11ou7ube_b[15:0]})
                   | ({64{s864qhdj_vmxevu9   }} & {e231c11ou7ube_b[71:40], e231c11ou7ube_b[31:0]})
                   | ({64{xd94m0cezzwq329zknc}} & {{32{e231c11ou7ube_b[31]}},e231c11ou7ube_b[31:0]})
                   | ({64{oc9vvnc_        }} & {e231c11ou7ube_b[63:0]})
                   ;





assign nb3w1rq_ny95rvrt = wj_jha74 ? ugh99u1va5po :
                         wl451sp6zo ? z8p8nm_hann2w4 : 
                         onsk4u1y9_e ? m2ngrd23vsh :
                         tdz9d9 ? ea1fw5akofqeu :
                         jxe3dht ? vt3rt5h12hv25u_6 : 64'b0;
						   






assign dkojj6fim0nxg4jvyafk = wj_jha74 ? kfxwyv6mbdgh :
                           bgh3d68j138h4ok_r7;


wire [yk7-1:0]         ylcp2s2rb7v6zuhdedv0h = n9mvknsj1brwzi9q3 ? {1'b0,zgg2kluk7qvo[0]} : zgg2kluk7qvo;
wire [yk7-1:0]         ogvd4x9j53t_fac02k = n9mvknsj1brwzi9q3 ? {1'b0,fz268jwgd_u7[0]} : fz268jwgd_u7;
wire ayv97dlbh0ci7olawv8 = lun9svt1 ? |{jxuls43sqwa,mj1ex47gsgf} :
                         hr7jjg ? |{romko5ymdrfzzldtl,jlhtbk3erojleuz_d} :
                         uayip3yhv ? |{ylcp2s2rb7v6zuhdedv0h,ogvd4x9j53t_fac02k} : 1'b0;

wire aoo0whg505i4exav193 = ((lun9svt1 & ru_hz78)   & (|{g3x1whn96j2yq4,h12hgjnbituwg32d6}))
                         | ((hr7jjg & b8qm5m9c4mc) & (|{fkjq_c0a1s83b0ab8,dnq81sp0s_88y0m3um}))
                         ;

assign vjkz8n6i44pc7o = ayv97dlbh0ci7olawv8 | aoo0whg505i4exav193;


endmodule



















module e2pg9lpkkc1p07id6ljjmll1r(
    input [64-1:0] u3sluj7j2sehfsy,
    input [64-1:0] xtl841cb0zo01b1f,
    input [32-1:0] tt2c87mcx6t7l4nazopbi8tufyyx2a,
    input [32-1:0] hexy9i9cx278g_gq1xa85w735098s,
    input [32-1:0] scnc2o0onmfzkunfbqlwf96_dqibfx5,
    input [32-1:0] ofydji25el_rhpy7qm466hp1a414dn,
    input gdebc5b6o6bv57ax1bw,
    input jl5uafxavxn4ffun,
    input b4wi1969mw9n534p,
    input hf3_u19xhtm47jygm346ih5592f,
    input niiot38ff0zsxxncd0u_5fljm__dl, 
    input pm3poaltg6mtmffm_87yhorfj9eort_, 
    input x1kaexv26aa2fd_7nz8w2t,
    output [63:0] usrh37qm6nz8yamj6_h_pmbv5,
    output [63:0] mipc_c8bfwk8khoqgtsj65f1f,
    output [63:0] pm3m6aucefl9oas0vqgwfm,
    output [63:0] yc5f_bw94gu1iari4qpmo269z,
    input fxk_v35ltu7y0_q6aadrtlvrl 
);

  wire [31:0]  kliaw77ijuhmkp7j;
  wire [31:0]  bk1g8ipth5ko58yud6s;
  wire [3:0] xtkz3ys1dkgji1r0whon8;
  wire [3:0] b6duomqhd0n_18tvaktgj;
  wire [7:0] yr4wjk5fwhr8y6330lzj;
  wire [7:0] b5ym7cok4l97ddig8;
  wire [16:0] ap5_59_uagoyagga20;
  wire [16:0] wj_jfjj58w1_mza;
  wire [16:0] mwmtdzhjf5nvx94so_0;
  wire [16:0] ak1454lmtzo468o;
  wire [16:0] k1tqxl_4te89ii72f;
  wire [16:0] hais7_mbqlaihy3f2;
  wire [16:0] uc9d81vxk5l8cw;
  wire [16:0] g_3998bc1nuo4ndc2as;
  wire [16:0] uy4kpukqylvx7x5u2; 
  wire [16:0] i72snoyr81kd29a; 
  wire [16:0] n3gmmegfj9lr61do; 
  wire [16:0] a_ag9c74seh44iszeni; 
  wire [16:0] cl4yicexhcu1m60h;
  wire [16:0] o08jfuwa9jfk_5pzc;
  wire [16:0] qj6t5fq1j9rxgyd0yo;
  wire [16:0] hksrg7y1zckh4trqz6;
  wire [15:0] evyo5rqy4s2hac61[0:4-1];
  wire [15:0] a5wqs01ckyzpd0tmo[0:4-1];
  wire [8:0] ktju422az9_bk1qyi [0:8-1];
  wire [8:0] jhrp4_1ewkw3t1dtpo5 [0:8-1];
  wire [8:0] t71yjbhu_iasb [0:8-1];
  wire [8:0] rfasz6b4hhxtzem [0:8-1];
  wire [7:0] lnsxqgrkkgs3[0:8-1];
  wire [7:0] u2uyjynwthp77[0:8-1];
  wire [15:0] cnaelowqu0ymg[0:8-1];
  wire signed [16:0] k34o2bl_37qo6__jtr0k[0:8-1];
  wire [31:0] qxh8w5u3c745gfsf[0:8-1];
  wire signed [32:0] gp46y0ajdwrqtrvlvj8eep_k[0:8-1];
  assign kliaw77ijuhmkp7j = u3sluj7j2sehfsy[63:32];
  assign bk1g8ipth5ko58yud6s = xtl841cb0zo01b1f[63:32];

  wire [7:0] n18wuasb4ft4w = u3sluj7j2sehfsy[7:0];
  wire [7:0] h0jt4fy_se = u3sluj7j2sehfsy[15:8];
  wire [7:0] vylyasnjvqv = u3sluj7j2sehfsy[23:16];
  wire [7:0] n8w4j2me47 = u3sluj7j2sehfsy[31:24];
  wire [7:0] u9uua39cmmk3gq = xtl841cb0zo01b1f[7:0];
  wire [7:0] jenirtz2ha9qz = xtl841cb0zo01b1f[15:8];
  wire [7:0] sjb6dsw6__h_b4b = xtl841cb0zo01b1f[23:16];
  wire [7:0] fxra2prun_r = xtl841cb0zo01b1f[31:24];

  wire [7:0] iye0fi056owm = kliaw77ijuhmkp7j[7:0];
  wire [7:0] o87ao8ercxs35 = kliaw77ijuhmkp7j[15:8];
  wire [7:0] yzk435hjdqy3 = kliaw77ijuhmkp7j[23:16];
  wire [7:0] nqlvhcmcu10lapc4y = kliaw77ijuhmkp7j[31:24];
  wire [7:0] xqaoliz6jx87j2 = bk1g8ipth5ko58yud6s[7:0];
  wire [7:0] lsl05qsz_96mld3 = bk1g8ipth5ko58yud6s[15:8];
  wire [7:0] xoc_wrb6clt9t = bk1g8ipth5ko58yud6s[23:16];
  wire [7:0] y8skhg2t5444 = bk1g8ipth5ko58yud6s[31:24];

  assign yr4wjk5fwhr8y6330lzj[0] = gdebc5b6o6bv57ax1bw & u3sluj7j2sehfsy[7]   ;
  assign yr4wjk5fwhr8y6330lzj[1] = gdebc5b6o6bv57ax1bw & u3sluj7j2sehfsy[15]  ;
  assign yr4wjk5fwhr8y6330lzj[2] = gdebc5b6o6bv57ax1bw & u3sluj7j2sehfsy[23]  ;
  assign yr4wjk5fwhr8y6330lzj[3] = gdebc5b6o6bv57ax1bw & u3sluj7j2sehfsy[31]  ;
  assign yr4wjk5fwhr8y6330lzj[4] = gdebc5b6o6bv57ax1bw & kliaw77ijuhmkp7j[7] ;
  assign yr4wjk5fwhr8y6330lzj[5] = gdebc5b6o6bv57ax1bw & kliaw77ijuhmkp7j[15];
  assign yr4wjk5fwhr8y6330lzj[6] = gdebc5b6o6bv57ax1bw & kliaw77ijuhmkp7j[23];
  assign yr4wjk5fwhr8y6330lzj[7] = gdebc5b6o6bv57ax1bw & kliaw77ijuhmkp7j[31]; 

  wire  ogcy7b6ipwxp1ihd79x3btg0fkxkd = (~fxk_v35ltu7y0_q6aadrtlvrl) & gdebc5b6o6bv57ax1bw;
  assign b5ym7cok4l97ddig8[0] = ogcy7b6ipwxp1ihd79x3btg0fkxkd & (x1kaexv26aa2fd_7nz8w2t ? xtl841cb0zo01b1f[15] : xtl841cb0zo01b1f[7]);
  assign b5ym7cok4l97ddig8[1] = ogcy7b6ipwxp1ihd79x3btg0fkxkd & (x1kaexv26aa2fd_7nz8w2t ? xtl841cb0zo01b1f[7] : xtl841cb0zo01b1f[15]);
  assign b5ym7cok4l97ddig8[2] = ogcy7b6ipwxp1ihd79x3btg0fkxkd & (x1kaexv26aa2fd_7nz8w2t ? xtl841cb0zo01b1f[31] : xtl841cb0zo01b1f[23]);
  assign b5ym7cok4l97ddig8[3] = ogcy7b6ipwxp1ihd79x3btg0fkxkd & (x1kaexv26aa2fd_7nz8w2t ? xtl841cb0zo01b1f[23] : xtl841cb0zo01b1f[31]);
  assign b5ym7cok4l97ddig8[4] = ogcy7b6ipwxp1ihd79x3btg0fkxkd & (x1kaexv26aa2fd_7nz8w2t ? bk1g8ipth5ko58yud6s[15] : bk1g8ipth5ko58yud6s[7]);
  assign b5ym7cok4l97ddig8[5] = ogcy7b6ipwxp1ihd79x3btg0fkxkd & (x1kaexv26aa2fd_7nz8w2t ? bk1g8ipth5ko58yud6s[7] : bk1g8ipth5ko58yud6s[15]);
  assign b5ym7cok4l97ddig8[6] = ogcy7b6ipwxp1ihd79x3btg0fkxkd & (x1kaexv26aa2fd_7nz8w2t ? bk1g8ipth5ko58yud6s[31] : bk1g8ipth5ko58yud6s[23]);
  assign b5ym7cok4l97ddig8[7] = ogcy7b6ipwxp1ihd79x3btg0fkxkd & (x1kaexv26aa2fd_7nz8w2t ? bk1g8ipth5ko58yud6s[23] : bk1g8ipth5ko58yud6s[31]);
  

  assign xtkz3ys1dkgji1r0whon8[0] = gdebc5b6o6bv57ax1bw & u3sluj7j2sehfsy[15];
  assign xtkz3ys1dkgji1r0whon8[1] = gdebc5b6o6bv57ax1bw & u3sluj7j2sehfsy[31];
  assign xtkz3ys1dkgji1r0whon8[2] = gdebc5b6o6bv57ax1bw & kliaw77ijuhmkp7j[15];
  assign xtkz3ys1dkgji1r0whon8[3] = gdebc5b6o6bv57ax1bw & kliaw77ijuhmkp7j[31];
  assign b6duomqhd0n_18tvaktgj[0] = gdebc5b6o6bv57ax1bw & xtl841cb0zo01b1f[15];
  assign b6duomqhd0n_18tvaktgj[1] = gdebc5b6o6bv57ax1bw & xtl841cb0zo01b1f[31];
  assign b6duomqhd0n_18tvaktgj[2] = gdebc5b6o6bv57ax1bw & bk1g8ipth5ko58yud6s[15];
  assign b6duomqhd0n_18tvaktgj[3] = gdebc5b6o6bv57ax1bw & bk1g8ipth5ko58yud6s[31];

  assign lnsxqgrkkgs3[0] = n18wuasb4ft4w;
  assign lnsxqgrkkgs3[1] = h0jt4fy_se;
  assign lnsxqgrkkgs3[2] = vylyasnjvqv;
  assign lnsxqgrkkgs3[3] = n8w4j2me47;
  assign lnsxqgrkkgs3[4] = iye0fi056owm;
  assign lnsxqgrkkgs3[5] = o87ao8ercxs35;
  assign lnsxqgrkkgs3[6] = yzk435hjdqy3;
  assign lnsxqgrkkgs3[7] = nqlvhcmcu10lapc4y;

  assign u2uyjynwthp77[0] = x1kaexv26aa2fd_7nz8w2t ? jenirtz2ha9qz   : u9uua39cmmk3gq;
  assign u2uyjynwthp77[1] = x1kaexv26aa2fd_7nz8w2t ? u9uua39cmmk3gq   : jenirtz2ha9qz;
  assign u2uyjynwthp77[2] = x1kaexv26aa2fd_7nz8w2t ? fxra2prun_r   : sjb6dsw6__h_b4b;
  assign u2uyjynwthp77[3] = x1kaexv26aa2fd_7nz8w2t ? sjb6dsw6__h_b4b   : fxra2prun_r;
  assign u2uyjynwthp77[4] = x1kaexv26aa2fd_7nz8w2t ? lsl05qsz_96mld3 : xqaoliz6jx87j2;
  assign u2uyjynwthp77[5] = x1kaexv26aa2fd_7nz8w2t ? xqaoliz6jx87j2 : lsl05qsz_96mld3;
  assign u2uyjynwthp77[6] = x1kaexv26aa2fd_7nz8w2t ? y8skhg2t5444 : xoc_wrb6clt9t;
  assign u2uyjynwthp77[7] = x1kaexv26aa2fd_7nz8w2t ? xoc_wrb6clt9t : y8skhg2t5444;

  assign evyo5rqy4s2hac61[0] = u3sluj7j2sehfsy[15:0];
  assign evyo5rqy4s2hac61[1] = u3sluj7j2sehfsy[31:16];
  assign evyo5rqy4s2hac61[2] = u3sluj7j2sehfsy[47:32];
  assign evyo5rqy4s2hac61[3] = u3sluj7j2sehfsy[63:48];
  assign a5wqs01ckyzpd0tmo[0] = xtl841cb0zo01b1f[15:0];
  assign a5wqs01ckyzpd0tmo[1] = xtl841cb0zo01b1f[31:16];
  assign a5wqs01ckyzpd0tmo[2] = xtl841cb0zo01b1f[47:32];
  assign a5wqs01ckyzpd0tmo[3] = xtl841cb0zo01b1f[63:48];

  assign ktju422az9_bk1qyi[0] = {yr4wjk5fwhr8y6330lzj[0],lnsxqgrkkgs3[0]};
  assign ktju422az9_bk1qyi[1] = {yr4wjk5fwhr8y6330lzj[1],lnsxqgrkkgs3[1]};
  assign ktju422az9_bk1qyi[2] = {yr4wjk5fwhr8y6330lzj[2],lnsxqgrkkgs3[2]};
  assign ktju422az9_bk1qyi[3] = {yr4wjk5fwhr8y6330lzj[3],lnsxqgrkkgs3[3]};
  assign ktju422az9_bk1qyi[4] = {yr4wjk5fwhr8y6330lzj[4],lnsxqgrkkgs3[4]};
  assign ktju422az9_bk1qyi[5] = {yr4wjk5fwhr8y6330lzj[5],lnsxqgrkkgs3[5]};
  assign ktju422az9_bk1qyi[6] = {yr4wjk5fwhr8y6330lzj[6],lnsxqgrkkgs3[6]};
  assign ktju422az9_bk1qyi[7] = {yr4wjk5fwhr8y6330lzj[7],lnsxqgrkkgs3[7]};

  assign jhrp4_1ewkw3t1dtpo5[0] = {b5ym7cok4l97ddig8[0],u2uyjynwthp77[0]};
  assign jhrp4_1ewkw3t1dtpo5[1] = {b5ym7cok4l97ddig8[1],u2uyjynwthp77[1]};
  assign jhrp4_1ewkw3t1dtpo5[2] = {b5ym7cok4l97ddig8[2],u2uyjynwthp77[2]};
  assign jhrp4_1ewkw3t1dtpo5[3] = {b5ym7cok4l97ddig8[3],u2uyjynwthp77[3]};
  assign jhrp4_1ewkw3t1dtpo5[4] = {b5ym7cok4l97ddig8[4],u2uyjynwthp77[4]};
  assign jhrp4_1ewkw3t1dtpo5[5] = {b5ym7cok4l97ddig8[5],u2uyjynwthp77[5]};
  assign jhrp4_1ewkw3t1dtpo5[6] = {b5ym7cok4l97ddig8[6],u2uyjynwthp77[6]};
  assign jhrp4_1ewkw3t1dtpo5[7] = {b5ym7cok4l97ddig8[7],u2uyjynwthp77[7]};

  assign t71yjbhu_iasb[0] = ktju422az9_bk1qyi[0];
  assign t71yjbhu_iasb[1] = ktju422az9_bk1qyi[1];
  assign t71yjbhu_iasb[2] = ktju422az9_bk1qyi[2];
  assign t71yjbhu_iasb[3] = ktju422az9_bk1qyi[3];
  assign t71yjbhu_iasb[4] = ktju422az9_bk1qyi[4];
  assign t71yjbhu_iasb[5] = ktju422az9_bk1qyi[5];
  assign t71yjbhu_iasb[6] = ktju422az9_bk1qyi[6];
  assign t71yjbhu_iasb[7] = ktju422az9_bk1qyi[7];
  assign rfasz6b4hhxtzem[0] = jhrp4_1ewkw3t1dtpo5[0];
  assign rfasz6b4hhxtzem[1] = jhrp4_1ewkw3t1dtpo5[1];
  assign rfasz6b4hhxtzem[2] = jhrp4_1ewkw3t1dtpo5[2];
  assign rfasz6b4hhxtzem[3] = jhrp4_1ewkw3t1dtpo5[3];
  assign rfasz6b4hhxtzem[4] = jhrp4_1ewkw3t1dtpo5[4];
  assign rfasz6b4hhxtzem[5] = jhrp4_1ewkw3t1dtpo5[5];
  assign rfasz6b4hhxtzem[6] = jhrp4_1ewkw3t1dtpo5[6];
  assign rfasz6b4hhxtzem[7] = jhrp4_1ewkw3t1dtpo5[7];

  assign ap5_59_uagoyagga20 = ({17{b4wi1969mw9n534p}} & {xtkz3ys1dkgji1r0whon8[0],evyo5rqy4s2hac61[0]})
                        | ({17{hf3_u19xhtm47jygm346ih5592f}} & {(niiot38ff0zsxxncd0u_5fljm__dl & tt2c87mcx6t7l4nazopbi8tufyyx2a[15]),tt2c87mcx6t7l4nazopbi8tufyyx2a[15:0]})
                        ;
  assign uy4kpukqylvx7x5u2 = ({17{b4wi1969mw9n534p & x1kaexv26aa2fd_7nz8w2t}} & {b6duomqhd0n_18tvaktgj[1],a5wqs01ckyzpd0tmo[1]})
                        | ({17{b4wi1969mw9n534p & (~x1kaexv26aa2fd_7nz8w2t)}} & {b6duomqhd0n_18tvaktgj[0],a5wqs01ckyzpd0tmo[0]})
                        | ({17{hf3_u19xhtm47jygm346ih5592f}} & {(niiot38ff0zsxxncd0u_5fljm__dl & hexy9i9cx278g_gq1xa85w735098s[15]),hexy9i9cx278g_gq1xa85w735098s[15:0]})
                        ;

  assign wj_jfjj58w1_mza = ({17{b4wi1969mw9n534p}} & {xtkz3ys1dkgji1r0whon8[1],evyo5rqy4s2hac61[1]})
                        | ({17{pm3poaltg6mtmffm_87yhorfj9eort_}} & {((gdebc5b6o6bv57ax1bw) & tt2c87mcx6t7l4nazopbi8tufyyx2a[31]),tt2c87mcx6t7l4nazopbi8tufyyx2a[31:16]})
                        ;
  assign i72snoyr81kd29a = ({17{b4wi1969mw9n534p & x1kaexv26aa2fd_7nz8w2t}} & {b6duomqhd0n_18tvaktgj[0],a5wqs01ckyzpd0tmo[0]})
                        | ({17{b4wi1969mw9n534p & (~x1kaexv26aa2fd_7nz8w2t)}} & {b6duomqhd0n_18tvaktgj[1],a5wqs01ckyzpd0tmo[1]})
                        | ({17{pm3poaltg6mtmffm_87yhorfj9eort_}} & {1'b0,hexy9i9cx278g_gq1xa85w735098s[15:0]})
                        ;

  assign mwmtdzhjf5nvx94so_0 = ({17{b4wi1969mw9n534p}} & {xtkz3ys1dkgji1r0whon8[2],evyo5rqy4s2hac61[2]})
                        | ({17{pm3poaltg6mtmffm_87yhorfj9eort_}} & {1'b0,tt2c87mcx6t7l4nazopbi8tufyyx2a[15:0]})
                        ;
  assign n3gmmegfj9lr61do = ({17{b4wi1969mw9n534p & x1kaexv26aa2fd_7nz8w2t}} & {b6duomqhd0n_18tvaktgj[3],a5wqs01ckyzpd0tmo[3]})
                        | ({17{b4wi1969mw9n534p & (~x1kaexv26aa2fd_7nz8w2t)}} & {b6duomqhd0n_18tvaktgj[2],a5wqs01ckyzpd0tmo[2]})
                        | ({17{pm3poaltg6mtmffm_87yhorfj9eort_}} & {((gdebc5b6o6bv57ax1bw) & hexy9i9cx278g_gq1xa85w735098s[31]),hexy9i9cx278g_gq1xa85w735098s[31:16]})
                        ;

  assign ak1454lmtzo468o = ({17{b4wi1969mw9n534p}} & {xtkz3ys1dkgji1r0whon8[3],evyo5rqy4s2hac61[3]})
                        | ({17{pm3poaltg6mtmffm_87yhorfj9eort_}} & {((gdebc5b6o6bv57ax1bw) & tt2c87mcx6t7l4nazopbi8tufyyx2a[31]),tt2c87mcx6t7l4nazopbi8tufyyx2a[31:16]})
                        ;
  assign a_ag9c74seh44iszeni = ({17{b4wi1969mw9n534p & x1kaexv26aa2fd_7nz8w2t}} & {b6duomqhd0n_18tvaktgj[2],a5wqs01ckyzpd0tmo[2]})
                        | ({17{b4wi1969mw9n534p & (~x1kaexv26aa2fd_7nz8w2t)}} & {b6duomqhd0n_18tvaktgj[3],a5wqs01ckyzpd0tmo[3]})
                        | ({17{pm3poaltg6mtmffm_87yhorfj9eort_}} & {((gdebc5b6o6bv57ax1bw) & hexy9i9cx278g_gq1xa85w735098s[31]),hexy9i9cx278g_gq1xa85w735098s[31:16]})
                        ;
  assign k1tqxl_4te89ii72f = ({17{pm3poaltg6mtmffm_87yhorfj9eort_}} & {((niiot38ff0zsxxncd0u_5fljm__dl) & scnc2o0onmfzkunfbqlwf96_dqibfx5[15]),scnc2o0onmfzkunfbqlwf96_dqibfx5[15:0]})
                        ;
  assign cl4yicexhcu1m60h = ({17{pm3poaltg6mtmffm_87yhorfj9eort_}} & {((niiot38ff0zsxxncd0u_5fljm__dl) & ofydji25el_rhpy7qm466hp1a414dn[15]),ofydji25el_rhpy7qm466hp1a414dn[15:0]})
                        ;

  assign hais7_mbqlaihy3f2 = ({17{pm3poaltg6mtmffm_87yhorfj9eort_}} & {((gdebc5b6o6bv57ax1bw) & scnc2o0onmfzkunfbqlwf96_dqibfx5[31]),scnc2o0onmfzkunfbqlwf96_dqibfx5[31:16]}) 
                        ;
  assign o08jfuwa9jfk_5pzc = ({17{pm3poaltg6mtmffm_87yhorfj9eort_}} & {1'b0,ofydji25el_rhpy7qm466hp1a414dn[15:0]})
                        ;

  assign uc9d81vxk5l8cw = ({17{pm3poaltg6mtmffm_87yhorfj9eort_}} & {1'b0,scnc2o0onmfzkunfbqlwf96_dqibfx5[15:0]})
                        ;
  assign qj6t5fq1j9rxgyd0yo = ({17{pm3poaltg6mtmffm_87yhorfj9eort_}} & {((gdebc5b6o6bv57ax1bw) & ofydji25el_rhpy7qm466hp1a414dn[31]),ofydji25el_rhpy7qm466hp1a414dn[31:16]})
                        ;

  assign g_3998bc1nuo4ndc2as = ({17{pm3poaltg6mtmffm_87yhorfj9eort_}} & {((gdebc5b6o6bv57ax1bw) & scnc2o0onmfzkunfbqlwf96_dqibfx5[31]),scnc2o0onmfzkunfbqlwf96_dqibfx5[31:16]})
                        ;
  assign hksrg7y1zckh4trqz6 = ({17{pm3poaltg6mtmffm_87yhorfj9eort_}} & {((gdebc5b6o6bv57ax1bw) & ofydji25el_rhpy7qm466hp1a414dn[31]),ofydji25el_rhpy7qm466hp1a414dn[31:16]})
                        ;

  assign k34o2bl_37qo6__jtr0k[0] = $signed(t71yjbhu_iasb[0]) * $signed(rfasz6b4hhxtzem[0]); 
  assign k34o2bl_37qo6__jtr0k[1] = $signed(t71yjbhu_iasb[1]) * $signed(rfasz6b4hhxtzem[1]); 
  assign k34o2bl_37qo6__jtr0k[2] = $signed(t71yjbhu_iasb[2]) * $signed(rfasz6b4hhxtzem[2]); 
  assign k34o2bl_37qo6__jtr0k[3] = $signed(t71yjbhu_iasb[3]) * $signed(rfasz6b4hhxtzem[3]); 
  assign k34o2bl_37qo6__jtr0k[4] = $signed(t71yjbhu_iasb[4]) * $signed(rfasz6b4hhxtzem[4]); 
  assign k34o2bl_37qo6__jtr0k[5] = $signed(t71yjbhu_iasb[5]) * $signed(rfasz6b4hhxtzem[5]); 
  assign k34o2bl_37qo6__jtr0k[6] = $signed(t71yjbhu_iasb[6]) * $signed(rfasz6b4hhxtzem[6]); 
  assign k34o2bl_37qo6__jtr0k[7] = $signed(t71yjbhu_iasb[7]) * $signed(rfasz6b4hhxtzem[7]); 
  assign gp46y0ajdwrqtrvlvj8eep_k[0] = $signed(ap5_59_uagoyagga20) * $signed(uy4kpukqylvx7x5u2);
  assign gp46y0ajdwrqtrvlvj8eep_k[1] = $signed(wj_jfjj58w1_mza) * $signed(i72snoyr81kd29a);
  assign gp46y0ajdwrqtrvlvj8eep_k[2] = $signed(mwmtdzhjf5nvx94so_0) * $signed(n3gmmegfj9lr61do);
  assign gp46y0ajdwrqtrvlvj8eep_k[3] = $signed(ak1454lmtzo468o) * $signed(a_ag9c74seh44iszeni);
  assign gp46y0ajdwrqtrvlvj8eep_k[4] = $signed(k1tqxl_4te89ii72f) * $signed(cl4yicexhcu1m60h);
  assign gp46y0ajdwrqtrvlvj8eep_k[5] = $signed(hais7_mbqlaihy3f2) * $signed(o08jfuwa9jfk_5pzc);
  assign gp46y0ajdwrqtrvlvj8eep_k[6] = $signed(uc9d81vxk5l8cw) * $signed(qj6t5fq1j9rxgyd0yo);
  assign gp46y0ajdwrqtrvlvj8eep_k[7] = $signed(g_3998bc1nuo4ndc2as) * $signed(hksrg7y1zckh4trqz6);

  assign cnaelowqu0ymg[0] = $unsigned(k34o2bl_37qo6__jtr0k[0][15:0]);
  assign cnaelowqu0ymg[1] = $unsigned(k34o2bl_37qo6__jtr0k[1][15:0]);
  assign cnaelowqu0ymg[2] = $unsigned(k34o2bl_37qo6__jtr0k[2][15:0]);
  assign cnaelowqu0ymg[3] = $unsigned(k34o2bl_37qo6__jtr0k[3][15:0]);
  assign cnaelowqu0ymg[4] = $unsigned(k34o2bl_37qo6__jtr0k[4][15:0]);
  assign cnaelowqu0ymg[5] = $unsigned(k34o2bl_37qo6__jtr0k[5][15:0]);
  assign cnaelowqu0ymg[6] = $unsigned(k34o2bl_37qo6__jtr0k[6][15:0]);
  assign cnaelowqu0ymg[7] = $unsigned(k34o2bl_37qo6__jtr0k[7][15:0]);
  assign qxh8w5u3c745gfsf[0] = $unsigned(gp46y0ajdwrqtrvlvj8eep_k[0][31:0]);
  assign qxh8w5u3c745gfsf[1] = $unsigned(gp46y0ajdwrqtrvlvj8eep_k[1][31:0]);
  assign qxh8w5u3c745gfsf[2] = $unsigned(gp46y0ajdwrqtrvlvj8eep_k[2][31:0]);
  assign qxh8w5u3c745gfsf[3] = $unsigned(gp46y0ajdwrqtrvlvj8eep_k[3][31:0]);
  assign qxh8w5u3c745gfsf[4] = $unsigned(gp46y0ajdwrqtrvlvj8eep_k[4][31:0]);
  assign qxh8w5u3c745gfsf[5] = $unsigned(gp46y0ajdwrqtrvlvj8eep_k[5][31:0]);
  assign qxh8w5u3c745gfsf[6] = $unsigned(gp46y0ajdwrqtrvlvj8eep_k[6][31:0]);
  assign qxh8w5u3c745gfsf[7] = $unsigned(gp46y0ajdwrqtrvlvj8eep_k[7][31:0]);
  assign usrh37qm6nz8yamj6_h_pmbv5 = ({64{b4wi1969mw9n534p | hf3_u19xhtm47jygm346ih5592f}} & {qxh8w5u3c745gfsf[1],qxh8w5u3c745gfsf[0]})
                              | ({64{jl5uafxavxn4ffun}} & {cnaelowqu0ymg[3],cnaelowqu0ymg[2],cnaelowqu0ymg[1],cnaelowqu0ymg[0]})
                              ;
  assign mipc_c8bfwk8khoqgtsj65f1f = ({64{b4wi1969mw9n534p | hf3_u19xhtm47jygm346ih5592f}} & {qxh8w5u3c745gfsf[3],qxh8w5u3c745gfsf[2]})
                              | ({64{jl5uafxavxn4ffun}} & {cnaelowqu0ymg[7],cnaelowqu0ymg[6],cnaelowqu0ymg[5],cnaelowqu0ymg[4]})
                              ;
  assign pm3m6aucefl9oas0vqgwfm = ({64{hf3_u19xhtm47jygm346ih5592f}} & {qxh8w5u3c745gfsf[5],qxh8w5u3c745gfsf[4]})
                              ;
  assign yc5f_bw94gu1iari4qpmo269z = ({64{hf3_u19xhtm47jygm346ih5592f}} & {qxh8w5u3c745gfsf[7],qxh8w5u3c745gfsf[6]});

endmodule







































































































module rrxf4gi2j6 #(
   parameter xio4kx7ep1ojwa_r      = 78,
   parameter cmnocc9r2aiw8za       = 8,
   parameter xholqktr732apzsv8d0  = 3
) (
    input                                    es6_9ffb14edb7t,                  
    input                                    mv5to8v6,                       
    
    input                                    ba9r7fnn73020zwu2mxj,              
    input                                    k3n1uuckanw669a,               
    input  [27-1:0]      qfy7pr76nvqld1f,               
    input  [1:0]                             nowfs1y75z9hmhv6r0ppp6vjly,        
    input                                    xtm2ue4np_4lj4a7ik,                        
    input  [26-1:0]    fsxy2ey9lgj3xvg2hw_sqfrgy,         
    input  [64-1:0]                  h5arfbj2deloqqwtp1,              
    input  [64-1:0]                  elgnxkek04s_nuz6z,              
    input                                    gcoematpqzttdb81ozfq3zg1v9,                        
    
    input                                    a9q83azb3dode6qt,

    
    output                                   yvy4oon7f_rsa81003k5snsy28,       
    output [26-1:0]    p761bsjfs381j2b7xfn02m8vbu4u,    
    output [20-1:0]         avdv23oy5gvvj_aozmzn5,         
    output                                   gojz6nraxpmhlx_7ewrhi6di9,        
    output                                   pxjlub1gdgqvcckianojxej7_mt,        
    output                                   ro2z68ba11neqxvjf0uqiz03nt,        
    output                                   ovl08q5ylus9d7r7ckvnrb0,        
    output                                   f6o85b68_amv01vbog6ngjt,        
    output                                   q5guxjr1bjcc5ehbwvbbdz6a__mpjv74z,  
    output                                   qkq4xk9dqb1zawk5qa22ux2h35d9lrg,


    output                                   lrn8i28ncm6vualne3lnezatrmx,        
    output [26-1:0]    d757aw4s0emlk_xndccuz9wrpek3n,     
    output [20-1:0]         ky4b1pzcyo6z1omquzzoj,          
    output                                   stcauj4mexs59diuva_xf1308li,         
    output                                   v_sj7f9mnvn2sgj37k1ave5g,         
    output                                   dce56zk48npvti3u7osyzacy,         
    output                                   dspbo9b1im8onetqwxjnw7,         
    output                                   kf99vegpc45l_wd1vhgluhfo65,         
    output                                   q0kprornbncukpltocigbw9tba03,   
    output                                   w_jjbyn9u5snyb45kcy8r78z6d9iz5, 
    output                                   faamp7iz46_jj1ci8a,             
    
    output                                   v66ux9ovjkzt3jn,                
    output  [27-1:0]     cd3lo77nievm4v3,                 
    output  [1:0]                            rgnht1zljy67subvhyua_,          
    output                                   uy22rssg5uc6vyiti9szp,
    output                                   h8djzt4zbmppcv2_ai,
    
    input                                    nmlix317bu48vgct7x02m7vgn,          
    input                                    s6zb15tq6xjiqgce5nwjcg7be4,     
    input                                    ry0rypry86op3l_hqbwk8pe32ena3e,   
    input  [xio4kx7ep1ojwa_r-1:0]              h4zmq2srkdf5iaeagd8d7i87,           
    input                                    dzo70vq3_1_kyxyiurxy1d20ed,         
    input                                    b0c0o6unssb9h3tgqck870,         

    
    output                                   c2_546oy8pb0vifo,                 
    input                                    gf33atgy,
    input                                    ru_wi,
    input                                    gc4b3kdcan6do88ta_
);

    localparam pse_9oeblmiqo   = 0;
    localparam bixr4rzvy34       = 1;
    localparam kbjnkuh       = 2;
    localparam cgidk92       = 3;
    localparam wh6wd1qdq2       = 4;
    localparam skhfe86rjzr       = 5;
    localparam c6bt4uxhjt76ybdb  = 6;
    localparam ir1y97hv4a9oct4l  = 7;
    localparam pvu039o1s9t1m9x_  = xio4kx7ep1ojwa_r-1;
    localparam obu455a2wnp4vu0  = pvu039o1s9t1m9x_+1-27;
    localparam snj9jgmwt45902 = obu455a2wnp4vu0-1;
    localparam la40sjjy7dga49 = snj9jgmwt45902+1-20;

    localparam rqzr_eaa     = 2'b00;
    localparam eri_rah_b     = 2'b01;
    localparam ib1cruu      = 2'b10;

    localparam b1lh2fnh92    = 2;

    localparam cpuuvz0x4_r5s = cmnocc9r2aiw8za-1;    




    genvar i;
    wire [xio4kx7ep1ojwa_r-1:0]                vsbxpc1qp3j8l [cmnocc9r2aiw8za-1:0];
    wire [cmnocc9r2aiw8za-1:0]                 i25ll1dii3u_d2n76;




    wire pj9rc44fi;
    wire vkm_fyjfzj9 = mv5to8v6 | b0c0o6unssb9h3tgqck870;
  ux607_clkgate u_oq26k57nedglq(
    .clk_in        (gf33atgy                    ),
    .clkgate_bypass(gc4b3kdcan6do88ta_         ),
    .clock_en      (vkm_fyjfzj9                ),
    .clk_out       (pj9rc44fi               )
  );




    wire [cmnocc9r2aiw8za-1:0]                 hw9pzy7xw26mqd67;
    wire [cmnocc9r2aiw8za-1:0]                 hnigkwjr_ezglt;
    wire [cmnocc9r2aiw8za-1:0]                 b7i5j5t_4whk_l2;
    wire [cmnocc9r2aiw8za-1:0]                 fhubgca2c9mrs;
    wire [cmnocc9r2aiw8za-1:0]                 d935qvi2jkbr_6n3;
    wire [cmnocc9r2aiw8za-1:0]                 pjisxg4auax56ugw;
    wire [1:0]                               wpxfw0jit8znrgcnnkq3he [cmnocc9r2aiw8za-1:0];
    wire [20-1:0]           ufhrnwb_tir83f [cmnocc9r2aiw8za-1:0];
    wire [27-1:0]        da5jkvbuwnfukf5p [cmnocc9r2aiw8za-1:0];

    wire [cmnocc9r2aiw8za-1:0]                 wskyn9jef_ao7fnlha;
    wire [cmnocc9r2aiw8za-1:0]                 yo5yfpeiuk3zechv7ry;
    wire [cmnocc9r2aiw8za-1:0]                 a_jrytlfkm3zom4pys8;
    wire [cmnocc9r2aiw8za-1:0]                 oqsatg3u7plwgaxlx8l;
    wire [cmnocc9r2aiw8za-1:0]                 ay8so07buwsbzd75a9;
    wire [cmnocc9r2aiw8za-1:0]                 pssati_l9flmulwcwpa820;
    wire [cmnocc9r2aiw8za-1:0]                 dqb744wwgwrkj8pmzlqz;
    reg  [xholqktr732apzsv8d0-1:0]            z0jov5agimrterpp2_e8sx6cjqcm;

    reg                                      kjhl4o5pi1i5qodyqewx;
    reg                                      bd82a9l7q7af53te0b0x;
    reg                                      vnqlzjx3yo4ma1dwa2;
    reg                                      ie77y48i7vsg8mclm8;
    reg                                      cpznd0fzt2newpz7w_;
    reg [1:0]                                t1xmqfke8fk5mqeub28crervpv9ocj;
    reg [20-1:0]            rtdki0i0xl5hvqfbkj371;


    wire udqn4evfqnp;
    wire eqb83t6;
    wire ku0a1r2r_h4;
    
    wire [39:0]                      bedhx0h5v3ki;
    wire                             utz9xevtl2wu;
    wire                             dfthmessjludvjd;
    wire                             wyfa30n_h0i2;
    wire                             scc4lj1z95m6;
    wire                             wphc19dg0fgz;
    wire                             ll1bfqtizvki9bzaw;
    wire [8:0]                       zft0wp87j7eq42;
    wire [8:0]                       cikk3phit89gu15z;
    wire [8:0]                       j6o83o1mu2mwcb;
    wire [8:0]                       l_hoppaexuxz2i;
    wire [8:0]                       jl48kanv3t6las;
    wire [8:0]                       e1asl5tgtgh8nro7lj;

    
    wire [8:0]         rzau5sna2h7g1xxei_7tzftbc [cmnocc9r2aiw8za-1:0];
    wire [8:0]         v4vyfn9vu7mi1j6qs0fs26f_k [cmnocc9r2aiw8za-1:0];
    wire [8:0]         hirqn5ba89vmhdyygl92c3j3l [cmnocc9r2aiw8za-1:0];
    wire [8:0]         nya00eozpx6ful79iac_0gzz0tl [cmnocc9r2aiw8za-1:0];
    wire [8:0]         fin1gyu2nfqkzd5j_fa1mikanqo5_ [cmnocc9r2aiw8za-1:0];
    wire [8:0]         gnoqp_ppw_9avgq5dlahpxno_1 [cmnocc9r2aiw8za-1:0];

    
    
    
    
    assign
    {  bedhx0h5v3ki[39:30] , ll1bfqtizvki9bzaw,
       bedhx0h5v3ki[29:21] , wphc19dg0fgz,
       bedhx0h5v3ki[20:12] , scc4lj1z95m6,
       bedhx0h5v3ki[11:0]                 } =   {h5arfbj2deloqqwtp1[39:30],1'b1,h5arfbj2deloqqwtp1[29:21],1'b1,h5arfbj2deloqqwtp1[20:12],1'b1,h5arfbj2deloqqwtp1[11:0]} 
                                              + {elgnxkek04s_nuz6z[39:30],1'b0,elgnxkek04s_nuz6z[29:21],1'b0,elgnxkek04s_nuz6z[20:12],1'b0,elgnxkek04s_nuz6z[11:0]}
                                              + {39'b0,gcoematpqzttdb81ozfq3zg1v9};

    assign utz9xevtl2wu = !scc4lj1z95m6;
    assign dfthmessjludvjd = !wphc19dg0fgz;
    assign wyfa30n_h0i2 = !ll1bfqtizvki9bzaw;
    assign zft0wp87j7eq42 = h5arfbj2deloqqwtp1[20:12] ^ elgnxkek04s_nuz6z[20:12];
    assign cikk3phit89gu15z = h5arfbj2deloqqwtp1[29:21] ^ elgnxkek04s_nuz6z[29:21];
    assign j6o83o1mu2mwcb = h5arfbj2deloqqwtp1[38:30] ^ elgnxkek04s_nuz6z[38:30];
    assign l_hoppaexuxz2i = h5arfbj2deloqqwtp1[20:12] & elgnxkek04s_nuz6z[20:12];
    assign jl48kanv3t6las = h5arfbj2deloqqwtp1[29:21] & elgnxkek04s_nuz6z[29:21];
    assign e1asl5tgtgh8nro7lj = h5arfbj2deloqqwtp1[38:30] & elgnxkek04s_nuz6z[38:30];


generate 
    for(i= 0; i<cmnocc9r2aiw8za; i=i+1) begin: n5jg7z9942w5zidr6
        assign hw9pzy7xw26mqd67[i]     = vsbxpc1qp3j8l[i][pse_9oeblmiqo];
        assign hnigkwjr_ezglt[i]         = vsbxpc1qp3j8l[i][bixr4rzvy34];
        assign b7i5j5t_4whk_l2[i]         = vsbxpc1qp3j8l[i][cgidk92];
        assign fhubgca2c9mrs[i]         = vsbxpc1qp3j8l[i][kbjnkuh];
        assign d935qvi2jkbr_6n3[i]         = vsbxpc1qp3j8l[i][wh6wd1qdq2];
        assign pjisxg4auax56ugw[i]         = vsbxpc1qp3j8l[i][skhfe86rjzr];
        assign wpxfw0jit8znrgcnnkq3he[i] = vsbxpc1qp3j8l[i][ir1y97hv4a9oct4l:c6bt4uxhjt76ybdb];
        assign ufhrnwb_tir83f[i]       = vsbxpc1qp3j8l[i][snj9jgmwt45902:la40sjjy7dga49];
        assign da5jkvbuwnfukf5p[i]        = vsbxpc1qp3j8l[i][pvu039o1s9t1m9x_:obu455a2wnp4vu0];
        assign wskyn9jef_ao7fnlha[i]   = wpxfw0jit8znrgcnnkq3he[i] == 2'b00;
        assign yo5yfpeiuk3zechv7ry[i]   = wpxfw0jit8znrgcnnkq3he[i] == 2'b01;
        assign a_jrytlfkm3zom4pys8[i]   = wpxfw0jit8znrgcnnkq3he[i] == 2'b10;

        assign rzau5sna2h7g1xxei_7tzftbc [i] = l_hoppaexuxz2i | (~vsbxpc1qp3j8l[i][obu455a2wnp4vu0 + 0*9 +: 9] & h5arfbj2deloqqwtp1[20:12]) | (~vsbxpc1qp3j8l[i][obu455a2wnp4vu0 + 0*9 +: 9] & elgnxkek04s_nuz6z[20:12]);
        assign hirqn5ba89vmhdyygl92c3j3l [i] = jl48kanv3t6las | (~vsbxpc1qp3j8l[i][obu455a2wnp4vu0 + 1*9 +: 9] & h5arfbj2deloqqwtp1[29:21]) | (~vsbxpc1qp3j8l[i][obu455a2wnp4vu0 + 1*9 +: 9] & elgnxkek04s_nuz6z[29:21]);
        assign fin1gyu2nfqkzd5j_fa1mikanqo5_ [i] = e1asl5tgtgh8nro7lj | (~vsbxpc1qp3j8l[i][obu455a2wnp4vu0 + 2*9 +: 9] & h5arfbj2deloqqwtp1[38:30]) | (~vsbxpc1qp3j8l[i][obu455a2wnp4vu0 + 2*9 +: 9] & elgnxkek04s_nuz6z[38:30]);
        assign v4vyfn9vu7mi1j6qs0fs26f_k   [i] = zft0wp87j7eq42 ^  ~vsbxpc1qp3j8l[i][obu455a2wnp4vu0 + 0*9 +: 9];
        assign nya00eozpx6ful79iac_0gzz0tl   [i] = cikk3phit89gu15z ^  ~vsbxpc1qp3j8l[i][obu455a2wnp4vu0 + 1*9 +: 9];
        assign gnoqp_ppw_9avgq5dlahpxno_1   [i] = j6o83o1mu2mwcb ^  ~vsbxpc1qp3j8l[i][obu455a2wnp4vu0 + 2*9 +: 9];

        assign oqsatg3u7plwgaxlx8l[i]  = &(v4vyfn9vu7mi1j6qs0fs26f_k[i] ^ ({rzau5sna2h7g1xxei_7tzftbc[i][7:0],utz9xevtl2wu}));
        assign ay8so07buwsbzd75a9[i]  = &(nya00eozpx6ful79iac_0gzz0tl[i] ^ ({hirqn5ba89vmhdyygl92c3j3l[i][7:0],dfthmessjludvjd}));
        assign pssati_l9flmulwcwpa820[i]  = &(gnoqp_ppw_9avgq5dlahpxno_1[i] ^ ({fin1gyu2nfqkzd5j_fa1mikanqo5_[i][7:0],wyfa30n_h0i2}));
        assign dqb744wwgwrkj8pmzlqz[i]     = ( 1'b0                 || pssati_l9flmulwcwpa820[i]) &&
                                        ( a_jrytlfkm3zom4pys8[i] || ay8so07buwsbzd75a9[i]) &&
                                        (!wskyn9jef_ao7fnlha[i] || oqsatg3u7plwgaxlx8l[i]) &&
                                          hw9pzy7xw26mqd67[i]
                                        ;
    end
endgenerate

    assign ku0a1r2r_h4 = |dqb744wwgwrkj8pmzlqz;
    assign eqb83t6     =  ku0a1r2r_h4 & k3n1uuckanw669a;
    assign udqn4evfqnp    = ~ku0a1r2r_h4 & k3n1uuckanw669a;


    integer j;
    always @(*) begin: vsxvdv5in4v_1f267wqv_2v
        kjhl4o5pi1i5qodyqewx = 1'b0;
        bd82a9l7q7af53te0b0x = 1'b0;
        vnqlzjx3yo4ma1dwa2 = 1'b0;
        ie77y48i7vsg8mclm8 = 1'b0;
        cpznd0fzt2newpz7w_ = 1'b0;
        t1xmqfke8fk5mqeub28crervpv9ocj = 2'b0;
        rtdki0i0xl5hvqfbkj371 = 20'b0;

        for (j=0; j<cmnocc9r2aiw8za; j=j+1) begin: wio55hb7s7eikmtdkw6
            kjhl4o5pi1i5qodyqewx = kjhl4o5pi1i5qodyqewx | (hnigkwjr_ezglt[j] & dqb744wwgwrkj8pmzlqz[j]);
            bd82a9l7q7af53te0b0x = bd82a9l7q7af53te0b0x | (b7i5j5t_4whk_l2[j] & dqb744wwgwrkj8pmzlqz[j]);
            vnqlzjx3yo4ma1dwa2 = vnqlzjx3yo4ma1dwa2 | (fhubgca2c9mrs[j] & dqb744wwgwrkj8pmzlqz[j]);
            ie77y48i7vsg8mclm8 = ie77y48i7vsg8mclm8 | (d935qvi2jkbr_6n3[j] & dqb744wwgwrkj8pmzlqz[j]);
            cpznd0fzt2newpz7w_ = cpznd0fzt2newpz7w_ | (pjisxg4auax56ugw[j] & dqb744wwgwrkj8pmzlqz[j]);
            t1xmqfke8fk5mqeub28crervpv9ocj = t1xmqfke8fk5mqeub28crervpv9ocj | (wpxfw0jit8znrgcnnkq3he[j] & {2{dqb744wwgwrkj8pmzlqz[j]}});
            rtdki0i0xl5hvqfbkj371 = rtdki0i0xl5hvqfbkj371 | (ufhrnwb_tir83f[j] & {20{dqb744wwgwrkj8pmzlqz[j]}});
        end
    end


    wire                                     twm0b4dd7ahh8f  =    dzo70vq3_1_kyxyiurxy1d20ed;
    wire                                     pubj1y308jtf6 =   (nmlix317bu48vgct7x02m7vgn & s6zb15tq6xjiqgce5nwjcg7be4  )
                                                            | (nmlix317bu48vgct7x02m7vgn & ry0rypry86op3l_hqbwk8pe32ena3e)
                                                            ;
    wire                                     ayqqbzrthvt93;
    wire                                     h624jgnv03hp4iysjt03z = eqb83t6 | twm0b4dd7ahh8f;
    wire                                     dyfajupgyhb37_vdc4elw = (eqb83t6 & ~ba9r7fnn73020zwu2mxj) | (twm0b4dd7ahh8f & ~ayqqbzrthvt93);
    wire                                     kt1oec5u1zomt6rpumj = (eqb83t6 & ba9r7fnn73020zwu2mxj) | (twm0b4dd7ahh8f &ayqqbzrthvt93);

    
    wire [cmnocc9r2aiw8za-1:0]                 cs4v4br38e3kc1mou;
    wire [cmnocc9r2aiw8za-1:0]                 jsb3cun4k6fukeall7w71;
    wire                                     prkeaifroj4g2dpakqjw;

    assign prkeaifroj4g2dpakqjw = h624jgnv03hp4iysjt03z;
    assign jsb3cun4k6fukeall7w71 = eqb83t6 ? dqb744wwgwrkj8pmzlqz : i25ll1dii3u_d2n76;
    ux607_gnrl_dfflr #(cmnocc9r2aiw8za) ijnyeqvww8x_chwcif9vbwi  (prkeaifroj4g2dpakqjw, jsb3cun4k6fukeall7w71, cs4v4br38e3kc1mou, gf33atgy, ru_wi);


    
    
    
    wire                                     k2iq1fadynzw7wzp0l0;
    wire                                     dn8u4c3b3oluzz8r0eta;
    wire                                     jbk57k2cscbog4x7ubvqu;

    assign jbk57k2cscbog4x7ubvqu = dyfajupgyhb37_vdc4elw;
    assign dn8u4c3b3oluzz8r0eta = eqb83t6 ? kjhl4o5pi1i5qodyqewx : h4zmq2srkdf5iaeagd8d7i87[bixr4rzvy34];
    ux607_gnrl_dfflr #(1) hf9ca_zyre50gs_psd0evt  (jbk57k2cscbog4x7ubvqu, dn8u4c3b3oluzz8r0eta, k2iq1fadynzw7wzp0l0, gf33atgy, ru_wi);

    
    wire                                     qgxdl96kyqmm_z6_vqw;
    wire                                     cle1bxl_u4dg0q2yaw;
    wire                                     p8h09lrjceoed7ijl;

    assign p8h09lrjceoed7ijl = dyfajupgyhb37_vdc4elw;
    assign cle1bxl_u4dg0q2yaw = eqb83t6 ? bd82a9l7q7af53te0b0x : h4zmq2srkdf5iaeagd8d7i87[cgidk92];
    ux607_gnrl_dfflr #(1) xnl6hx_a8iif0tvcz2w_c  (p8h09lrjceoed7ijl, cle1bxl_u4dg0q2yaw, qgxdl96kyqmm_z6_vqw, gf33atgy, ru_wi);

    
    wire                                     ffo1jrw6y2afg69e;
    wire                                     p2p7_2l8wvkex1g872t;
    wire                                     l39k5eut92oxksws;

    assign l39k5eut92oxksws = dyfajupgyhb37_vdc4elw;
    assign p2p7_2l8wvkex1g872t = eqb83t6 ? vnqlzjx3yo4ma1dwa2 : h4zmq2srkdf5iaeagd8d7i87[kbjnkuh];
    ux607_gnrl_dfflr #(1) h3sa1r6s9ja_h304xpk_  (l39k5eut92oxksws, p2p7_2l8wvkex1g872t, ffo1jrw6y2afg69e, gf33atgy, ru_wi);

    
    wire                                     fouse5g_ouj8b6we9;
    wire                                     hsc2dee4baq9cemtsh;
    wire                                     za059er_oz19zlqnzecd;

    assign za059er_oz19zlqnzecd = dyfajupgyhb37_vdc4elw;
    assign hsc2dee4baq9cemtsh = eqb83t6 ? ie77y48i7vsg8mclm8 : h4zmq2srkdf5iaeagd8d7i87[wh6wd1qdq2];
    ux607_gnrl_dfflr #(1) yl287_ylvhwaxti2_a8q  (za059er_oz19zlqnzecd, hsc2dee4baq9cemtsh, fouse5g_ouj8b6we9, gf33atgy, ru_wi);

    
    wire                                     u7ojjt008cvz5fxy;
    wire                                     wd2fxreyp_nnvnkip;
    wire                                     nw6lypdp24pr0apqg5z;

    assign nw6lypdp24pr0apqg5z = dyfajupgyhb37_vdc4elw;
    assign wd2fxreyp_nnvnkip = eqb83t6 ? cpznd0fzt2newpz7w_ : h4zmq2srkdf5iaeagd8d7i87[skhfe86rjzr];
    ux607_gnrl_dfflr #(1) j_bj7ds6bpdl9vp91  (nw6lypdp24pr0apqg5z, wd2fxreyp_nnvnkip, u7ojjt008cvz5fxy, gf33atgy, ru_wi);

    
    wire [1:0]                               p9frop7brmle_jm0khe2owdtd;
    wire [1:0]                               icw0skcu8uf8t7hiq4p35nip;
    wire                                     f366i7bawybnunt3kx2nxe9eqxj;

    assign f366i7bawybnunt3kx2nxe9eqxj = dyfajupgyhb37_vdc4elw;
    assign icw0skcu8uf8t7hiq4p35nip = eqb83t6 ? t1xmqfke8fk5mqeub28crervpv9ocj : h4zmq2srkdf5iaeagd8d7i87[ir1y97hv4a9oct4l:c6bt4uxhjt76ybdb];
    ux607_gnrl_dfflr #(2) od6jd8cvvriflfae1d7pdmhh5435  (f366i7bawybnunt3kx2nxe9eqxj, icw0skcu8uf8t7hiq4p35nip, p9frop7brmle_jm0khe2owdtd, gf33atgy, ru_wi);

    
    wire [20-1:0]           w1iqy20cnlpnd5hflpqy_;
    wire [20-1:0]           lm9eg685zlu9y59op9fg_s1;
    wire                                     ytyhsorz5j6gzm_nhv;

    assign ytyhsorz5j6gzm_nhv = dyfajupgyhb37_vdc4elw;
    assign lm9eg685zlu9y59op9fg_s1 = eqb83t6 ? rtdki0i0xl5hvqfbkj371 : h4zmq2srkdf5iaeagd8d7i87[snj9jgmwt45902:la40sjjy7dga49];
    ux607_gnrl_dfflr  #(20) wdeesqqte3f_nz8qfs1yvo0m (ytyhsorz5j6gzm_nhv, lm9eg685zlu9y59op9fg_s1, w1iqy20cnlpnd5hflpqy_, gf33atgy, ru_wi);

    wire [20-1:0]           th4w08jy003d95gfdsuxyi;
    wire                                     kuhud6tga9qt9y77qmkifhs5jbj;
    wire                                     n2aoj5pg0g6om07rzr3l58ngwso;
    wire [20-1:0]           re59d1fkoqi2m9vdfr65;
    wire [20-1:0]           jc2um6ob799jklbpoe;
    wire [27-1:0]        cq30mwyfhqwa;

    assign kuhud6tga9qt9y77qmkifhs5jbj = (p9frop7brmle_jm0khe2owdtd == 2'b00);
    assign n2aoj5pg0g6om07rzr3l58ngwso = (p9frop7brmle_jm0khe2owdtd == 2'b01);
    assign re59d1fkoqi2m9vdfr65    = kuhud6tga9qt9y77qmkifhs5jbj ? {20{1'b1}} :
                                      n2aoj5pg0g6om07rzr3l58ngwso ? {{20-9{1'b1}}, 9'b0} :
                                      {{20-18{1'b1}}, 18'b0};
    assign jc2um6ob799jklbpoe          = {{20-18{1'b0}}, cq30mwyfhqwa[17:0]};

    assign th4w08jy003d95gfdsuxyi = (w1iqy20cnlpnd5hflpqy_ & re59d1fkoqi2m9vdfr65) | (jc2um6ob799jklbpoe & ~re59d1fkoqi2m9vdfr65);
    
    wire [26-1:0]      zmxmooo4wvcx2e65u0o70qz00;
    wire [26-1:0]      p3n0ufpmzb7a3qicbclpwngd9;
    wire                                     xsnqbd8b9xnbarm150g22o410e;
    assign xsnqbd8b9xnbarm150g22o410e = k3n1uuckanw669a & ~ba9r7fnn73020zwu2mxj;
    assign p3n0ufpmzb7a3qicbclpwngd9 = fsxy2ey9lgj3xvg2hw_sqfrgy;
    ux607_gnrl_dfflr  #(26) ts7rvesm28ihiyl8uk79gsl44 (xsnqbd8b9xnbarm150g22o410e, p3n0ufpmzb7a3qicbclpwngd9, zmxmooo4wvcx2e65u0o70qz00, gf33atgy, ru_wi);

    
    
    wire [27-1:0]        t5ylupwx64ytnhyg4;
    wire                                     yqatidd9aw6r9_5;

    assign yqatidd9aw6r9_5     = k3n1uuckanw669a & ~ba9r7fnn73020zwu2mxj;   
    assign t5ylupwx64ytnhyg4  = qfy7pr76nvqld1f;
    ux607_gnrl_dfflr #(27) usdacoa8c57n8ofbge8 (yqatidd9aw6r9_5, t5ylupwx64ytnhyg4, cq30mwyfhqwa, gf33atgy, ru_wi);

    
    
    
    wire                                     yjuujp8x84pgx57z0kn;
    wire                                     g17mb30b8ydiy2ga0;
    wire                                     ziptbtdm6e6gyr15nxbd;

    assign ziptbtdm6e6gyr15nxbd = kt1oec5u1zomt6rpumj;
    assign g17mb30b8ydiy2ga0 = eqb83t6 ? kjhl4o5pi1i5qodyqewx : h4zmq2srkdf5iaeagd8d7i87[bixr4rzvy34];
    ux607_gnrl_dfflr #(1) mxk3af7porwtgsall6sp0  (ziptbtdm6e6gyr15nxbd, g17mb30b8ydiy2ga0, yjuujp8x84pgx57z0kn, gf33atgy, ru_wi);

    
    wire                                     dh2xowtqx9d9mq_icq5;
    wire                                     b2c3p645r_cttxt2;
    wire                                     zbvjr45dj8atgv91;

    assign zbvjr45dj8atgv91 = kt1oec5u1zomt6rpumj;
    assign b2c3p645r_cttxt2 = eqb83t6 ? bd82a9l7q7af53te0b0x : h4zmq2srkdf5iaeagd8d7i87[cgidk92];
    ux607_gnrl_dfflr #(1) tgu98log3buxlt5zerf3wq  (zbvjr45dj8atgv91, b2c3p645r_cttxt2, dh2xowtqx9d9mq_icq5, gf33atgy, ru_wi);

    
    wire                                     yqqbs3_6flcq_idm;
    wire                                     h66ttcu744z0o4wa;
    wire                                     npijj1n86ybscn3j;

    assign npijj1n86ybscn3j = kt1oec5u1zomt6rpumj;
    assign h66ttcu744z0o4wa = eqb83t6 ? vnqlzjx3yo4ma1dwa2 : h4zmq2srkdf5iaeagd8d7i87[kbjnkuh];
    ux607_gnrl_dfflr #(1) ipfuarkjmth_plovtj  (npijj1n86ybscn3j, h66ttcu744z0o4wa, yqqbs3_6flcq_idm, gf33atgy, ru_wi);

    
    wire                                     j5934321vs15d6dj;
    wire                                     dcjcleg3gnq6c423g2;
    wire                                     prpx3mtfb1es78_lwy;

    assign prpx3mtfb1es78_lwy = kt1oec5u1zomt6rpumj;
    assign dcjcleg3gnq6c423g2 = eqb83t6 ? ie77y48i7vsg8mclm8 : h4zmq2srkdf5iaeagd8d7i87[wh6wd1qdq2];
    ux607_gnrl_dfflr #(1) hcculs6s606q3h51v1c7ox  (prpx3mtfb1es78_lwy, dcjcleg3gnq6c423g2, j5934321vs15d6dj, gf33atgy, ru_wi);

    
    wire                                     gx5bpb6ffz6f__05cr;
    wire                                     vf0u0go71y9nioca;
    wire                                     pkug_3q925jjg5cs83;

    assign pkug_3q925jjg5cs83 = kt1oec5u1zomt6rpumj;
    assign vf0u0go71y9nioca = eqb83t6 ? cpznd0fzt2newpz7w_ : h4zmq2srkdf5iaeagd8d7i87[skhfe86rjzr];
    ux607_gnrl_dfflr #(1) jifitnk0rve7h39pjqv_  (pkug_3q925jjg5cs83, vf0u0go71y9nioca, gx5bpb6ffz6f__05cr, gf33atgy, ru_wi);

    
    wire [1:0]                               sjulazmgchq2b9fioxgko8wpms;
    wire [1:0]                               dfofhmtskslyx0k2b042y37_f39;
    wire                                     pl2gg8yglok1lfwovn2g4atvhr;

    assign pl2gg8yglok1lfwovn2g4atvhr = kt1oec5u1zomt6rpumj;
    assign dfofhmtskslyx0k2b042y37_f39 = eqb83t6 ? t1xmqfke8fk5mqeub28crervpv9ocj : h4zmq2srkdf5iaeagd8d7i87[ir1y97hv4a9oct4l:c6bt4uxhjt76ybdb];
    ux607_gnrl_dfflr #(2) rs4wh76_u523z6cd1gs8upp9jh  (pl2gg8yglok1lfwovn2g4atvhr, dfofhmtskslyx0k2b042y37_f39, sjulazmgchq2b9fioxgko8wpms, gf33atgy, ru_wi);

    
    wire [20-1:0]           o79bcp0v2kv7jcot00nz;
    wire [20-1:0]           stbeapnmxvyt2_jx38l;
    wire                                     melwgjj38qq367sojwpgm1;

    assign melwgjj38qq367sojwpgm1 = kt1oec5u1zomt6rpumj;
    assign stbeapnmxvyt2_jx38l = eqb83t6 ? rtdki0i0xl5hvqfbkj371 : h4zmq2srkdf5iaeagd8d7i87[snj9jgmwt45902:la40sjjy7dga49];
    ux607_gnrl_dfflr  #(20) xn9sn9itv7o21t6d1l64a (melwgjj38qq367sojwpgm1, stbeapnmxvyt2_jx38l, o79bcp0v2kv7jcot00nz, gf33atgy, ru_wi);

    wire [20-1:0]           vneu1upjrxltagmeu7x;
    wire                                     qjr88q0o08c1t5yiv63ufl8;
    wire                                     kr53a5tsn6v4ixody_t56uw;
    wire [20-1:0]           uhi4dwn0ol3z96u3r4to8;
    wire [20-1:0]           dgf5fj2vjwhmr5p0;
    wire [27-1:0]        qbo1b11wky6gxke_;

    assign qjr88q0o08c1t5yiv63ufl8 = (sjulazmgchq2b9fioxgko8wpms == 2'b00);
    assign kr53a5tsn6v4ixody_t56uw = (sjulazmgchq2b9fioxgko8wpms == 2'b01);
    assign uhi4dwn0ol3z96u3r4to8    = qjr88q0o08c1t5yiv63ufl8 ? {20{1'b1}} :
                                      kr53a5tsn6v4ixody_t56uw ? {{20-9{1'b1}}, 9'b0} :
                                      {{20-18{1'b1}}, 18'b0};
    assign dgf5fj2vjwhmr5p0          = {{20-18{1'b0}}, qbo1b11wky6gxke_[17:0]};

    assign vneu1upjrxltagmeu7x = (o79bcp0v2kv7jcot00nz & uhi4dwn0ol3z96u3r4to8) | (dgf5fj2vjwhmr5p0 & ~uhi4dwn0ol3z96u3r4to8);
    
    wire [26-1:0]      d6ihhd9s3mwhlwqpcw9o0xq;
    wire [26-1:0]      ywlfdz180iy6ldp7a_sdxf7w;
    wire                                     hkuh1gs9i0pdc628876e9w_kc4g;
    assign hkuh1gs9i0pdc628876e9w_kc4g = k3n1uuckanw669a & ba9r7fnn73020zwu2mxj;
    assign ywlfdz180iy6ldp7a_sdxf7w = fsxy2ey9lgj3xvg2hw_sqfrgy;
    ux607_gnrl_dfflr  #(26) fbphy8n5ea07nnnudjnoa5seqw8 (hkuh1gs9i0pdc628876e9w_kc4g, ywlfdz180iy6ldp7a_sdxf7w, d6ihhd9s3mwhlwqpcw9o0xq, gf33atgy, ru_wi);

    
    
    wire [27-1:0]        p9pe2g4_4tqbrjsr;
    wire                                     ee8bq7w082zv_c;

    assign ee8bq7w082zv_c     = k3n1uuckanw669a & ba9r7fnn73020zwu2mxj;   
    assign p9pe2g4_4tqbrjsr  = qfy7pr76nvqld1f;
    ux607_gnrl_dfflr #(27) n8rwawictg7_6xw (ee8bq7w082zv_c, p9pe2g4_4tqbrjsr, qbo1b11wky6gxke_, gf33atgy, ru_wi);

    
    wire [1:0]                               wdmmpqdswy4kjj3h31ammx;
    wire [1:0]                               ry4hr887uddag55rijdf;
    wire                                     cbho67y3xn6i3qlrzbpii;

    assign cbho67y3xn6i3qlrzbpii     = k3n1uuckanw669a;   
    assign ry4hr887uddag55rijdf  = nowfs1y75z9hmhv6r0ppp6vjly;
    ux607_gnrl_dfflr #(2) x_9qx902y0e8kr2mn2br02u4 (cbho67y3xn6i3qlrzbpii, ry4hr887uddag55rijdf, wdmmpqdswy4kjj3h31ammx, gf33atgy, ru_wi);

    wire                                     zaab503am_hhz0afn;
    wire                                     islvmtohfnuv1yc8mv;
    wire                                     jcmibolyq7z_wmf21lnw;

    assign jcmibolyq7z_wmf21lnw     = k3n1uuckanw669a;   
    assign islvmtohfnuv1yc8mv  = xtm2ue4np_4lj4a7ik;
    ux607_gnrl_dfflr #(1) fmcnqcbrs8xpi3__ca2c (jcmibolyq7z_wmf21lnw, islvmtohfnuv1yc8mv, zaab503am_hhz0afn, gf33atgy, ru_wi);

    
    wire                                     whpmltdnnmuxptumq;
    wire                                     dqbg_iv8botjtanoa;
    wire                                     nhtgbu_4g0hkmbntq;

    assign nhtgbu_4g0hkmbntq    = udqn4evfqnp;   
    assign dqbg_iv8botjtanoa =!a9q83azb3dode6qt;
    ux607_gnrl_dfflr #(1) evditodto8hn21z6 (nhtgbu_4g0hkmbntq, dqbg_iv8botjtanoa, whpmltdnnmuxptumq, gf33atgy, ru_wi);

    
    wire                                     ae0u6lggf97n7el;
    wire                                     elk8xd86q_z1rck7oqh;
    wire                                     msew56fe20a3zu1ts9;
    assign msew56fe20a3zu1ts9     = k3n1uuckanw669a;   
    assign elk8xd86q_z1rck7oqh     = ba9r7fnn73020zwu2mxj;
    ux607_gnrl_dfflr #(1) pmwegl0g474ci7zj50j (msew56fe20a3zu1ts9, elk8xd86q_z1rck7oqh, ae0u6lggf97n7el, gf33atgy, ru_wi);

    assign ayqqbzrthvt93 = ae0u6lggf97n7el;




    wire [xio4kx7ep1ojwa_r-1:0]                unj96xqpx4osi2 [cmnocc9r2aiw8za-1:0];
    wire [cmnocc9r2aiw8za-1:0]                 sgncc5i359h6_b7y9;
generate 
    for(i=0; i<cmnocc9r2aiw8za; i=i+1) begin: mpi9jkoirzo4ev3ab
        assign sgncc5i359h6_b7y9[i] = mv5to8v6 | (twm0b4dd7ahh8f & i25ll1dii3u_d2n76[i]);
        assign unj96xqpx4osi2[i] = mv5to8v6 ? {xio4kx7ep1ojwa_r{1'b0}} : h4zmq2srkdf5iaeagd8d7i87;

        ux607_gnrl_dfflr #(xio4kx7ep1ojwa_r) koqjnfv662ks1 (sgncc5i359h6_b7y9[i], unj96xqpx4osi2[i], vsbxpc1qp3j8l[i], pj9rc44fi, ru_wi);
    end
endgenerate




wire [cpuuvz0x4_r5s-1:0] blk93p1i16xx;
wire xtuu_xtcsg4icbv_ = &hw9pzy7xw26mqd67; 
wire [cpuuvz0x4_r5s-1:0] vs7xk5fv2idvsx3b;
wire [cmnocc9r2aiw8za-1:0] tmtwlbn11k8pot_5kb;
wire [cmnocc9r2aiw8za-1:0] j6u1lgj0jf7udo;
wire [cmnocc9r2aiw8za-1:0] bnrmlmaiin9wudfye9v7j7; 

assign bnrmlmaiin9wudfye9v7j7 =  dqb744wwgwrkj8pmzlqz;

generate
if(cmnocc9r2aiw8za ==16) begin:vt5kaq6
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   

    assign tmtwlbn11k8pot_5kb[0]  = ~blk93p1i16xx[7]  &  ~blk93p1i16xx[3] & ~blk93p1i16xx[1] &  ~blk93p1i16xx[0] & xtuu_xtcsg4icbv_;
    assign tmtwlbn11k8pot_5kb[1]  =  blk93p1i16xx[7]  &  ~blk93p1i16xx[3] & ~blk93p1i16xx[1] &  ~blk93p1i16xx[0] & xtuu_xtcsg4icbv_;
    assign tmtwlbn11k8pot_5kb[2]  = ~blk93p1i16xx[8]  &   blk93p1i16xx[3] & ~blk93p1i16xx[1] &  ~blk93p1i16xx[0] & xtuu_xtcsg4icbv_;
    assign tmtwlbn11k8pot_5kb[3]  =  blk93p1i16xx[8]  &   blk93p1i16xx[3] & ~blk93p1i16xx[1] &  ~blk93p1i16xx[0] & xtuu_xtcsg4icbv_;
    assign tmtwlbn11k8pot_5kb[4]  = ~blk93p1i16xx[9]  &  ~blk93p1i16xx[4] &  blk93p1i16xx[1] &  ~blk93p1i16xx[0] & xtuu_xtcsg4icbv_;
    assign tmtwlbn11k8pot_5kb[5]  =  blk93p1i16xx[9]  &  ~blk93p1i16xx[4] &  blk93p1i16xx[1] &  ~blk93p1i16xx[0] & xtuu_xtcsg4icbv_;
    assign tmtwlbn11k8pot_5kb[6]  = ~blk93p1i16xx[10] &   blk93p1i16xx[4] &  blk93p1i16xx[1] &  ~blk93p1i16xx[0] & xtuu_xtcsg4icbv_;
    assign tmtwlbn11k8pot_5kb[7]  =  blk93p1i16xx[10] &   blk93p1i16xx[4] &  blk93p1i16xx[1] &  ~blk93p1i16xx[0] & xtuu_xtcsg4icbv_;
    assign tmtwlbn11k8pot_5kb[8]  = ~blk93p1i16xx[11] &  ~blk93p1i16xx[5] & ~blk93p1i16xx[2] &   blk93p1i16xx[0] & xtuu_xtcsg4icbv_;
    assign tmtwlbn11k8pot_5kb[9]  =  blk93p1i16xx[11] &  ~blk93p1i16xx[5] & ~blk93p1i16xx[2] &   blk93p1i16xx[0] & xtuu_xtcsg4icbv_;
    assign tmtwlbn11k8pot_5kb[10] = ~blk93p1i16xx[12] &   blk93p1i16xx[5] & ~blk93p1i16xx[2] &   blk93p1i16xx[0] & xtuu_xtcsg4icbv_;
    assign tmtwlbn11k8pot_5kb[11] =  blk93p1i16xx[12] &   blk93p1i16xx[5] & ~blk93p1i16xx[2] &   blk93p1i16xx[0] & xtuu_xtcsg4icbv_;
    assign tmtwlbn11k8pot_5kb[12] = ~blk93p1i16xx[13] &  ~blk93p1i16xx[6] &  blk93p1i16xx[2] &   blk93p1i16xx[0] & xtuu_xtcsg4icbv_;
    assign tmtwlbn11k8pot_5kb[13] =  blk93p1i16xx[13] &  ~blk93p1i16xx[6] &  blk93p1i16xx[2] &   blk93p1i16xx[0] & xtuu_xtcsg4icbv_;
    assign tmtwlbn11k8pot_5kb[14] = ~blk93p1i16xx[14] &   blk93p1i16xx[6] &  blk93p1i16xx[2] &   blk93p1i16xx[0] & xtuu_xtcsg4icbv_;
    assign tmtwlbn11k8pot_5kb[15] =  blk93p1i16xx[14] &   blk93p1i16xx[6] &  blk93p1i16xx[2] &   blk93p1i16xx[0] & xtuu_xtcsg4icbv_;

    assign vs7xk5fv2idvsx3b = ({15{j6u1lgj0jf7udo[0]}} & {blk93p1i16xx[14:8],1'b1,blk93p1i16xx[6:4],1'b1,blk93p1i16xx[2], 2'b11}) |
                             ({15{j6u1lgj0jf7udo[1]}} & {blk93p1i16xx[14:8],1'b0,blk93p1i16xx[6:4],1'b1,blk93p1i16xx[2], 2'b11}) |
                             ({15{j6u1lgj0jf7udo[2]}} & {blk93p1i16xx[14:9],1'b1,blk93p1i16xx[7:4],1'b0,blk93p1i16xx[2], 2'b11}) |
                             ({15{j6u1lgj0jf7udo[3]}} & {blk93p1i16xx[14:9],1'b0,blk93p1i16xx[7:4],1'b0,blk93p1i16xx[2], 2'b11}) |
                             ({15{j6u1lgj0jf7udo[4]}} & {blk93p1i16xx[14:10],1'b1,blk93p1i16xx[8:5],1'b1,blk93p1i16xx[3:2], 2'b01}) |
                             ({15{j6u1lgj0jf7udo[5]}} & {blk93p1i16xx[14:10],1'b0,blk93p1i16xx[8:5],1'b1,blk93p1i16xx[3:2], 2'b01}) |
                             ({15{j6u1lgj0jf7udo[6]}} & {blk93p1i16xx[14:11],1'b1,blk93p1i16xx[9:5],1'b0,blk93p1i16xx[3:2], 2'b01}) |
                             ({15{j6u1lgj0jf7udo[7]}} & {blk93p1i16xx[14:11],1'b0,blk93p1i16xx[9:5],1'b0,blk93p1i16xx[3:2], 2'b01}) |
                             ({15{j6u1lgj0jf7udo[8]}} & {blk93p1i16xx[14:12],1'b1,blk93p1i16xx[10:6],1'b1,blk93p1i16xx[4:3],  1'b1,blk93p1i16xx[1],1'b0}) |
                             ({15{j6u1lgj0jf7udo[9]}} & {blk93p1i16xx[14:12],1'b0,blk93p1i16xx[10:6],1'b1,blk93p1i16xx[4:3],  1'b1,blk93p1i16xx[1],1'b0}) |
                             ({15{j6u1lgj0jf7udo[10]}} & {blk93p1i16xx[14:13],1'b1,blk93p1i16xx[11:6],1'b0,blk93p1i16xx[4:3], 1'b1,blk93p1i16xx[1],1'b0}) |
                             ({15{j6u1lgj0jf7udo[11]}} & {blk93p1i16xx[14:13],1'b0,blk93p1i16xx[11:6],1'b0,blk93p1i16xx[4:3], 1'b1,blk93p1i16xx[1],1'b0}) |
                             ({15{j6u1lgj0jf7udo[12]}} & {blk93p1i16xx[14],1'b1,blk93p1i16xx[12:7],1'b1,blk93p1i16xx[5:3],  1'b0,blk93p1i16xx[1],1'b0}) |
                             ({15{j6u1lgj0jf7udo[13]}} & {blk93p1i16xx[14],1'b0,blk93p1i16xx[12:7],1'b1,blk93p1i16xx[5:3],  1'b0,blk93p1i16xx[1],1'b0}) |
                             ({15{j6u1lgj0jf7udo[14]}} & {1'b1,blk93p1i16xx[13:7],1'b0,blk93p1i16xx[5:3], 1'b0,blk93p1i16xx[1],1'b0}) |
                             ({15{j6u1lgj0jf7udo[15]}} & {1'b0,blk93p1i16xx[13:7],1'b0,blk93p1i16xx[5:3], 1'b0,blk93p1i16xx[1],1'b0});
end
else if(cmnocc9r2aiw8za ==8) begin:g62rpi2e
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   

    assign tmtwlbn11k8pot_5kb[0]  = ~blk93p1i16xx[3] & ~blk93p1i16xx[1] &  ~blk93p1i16xx[0] & xtuu_xtcsg4icbv_;
    assign tmtwlbn11k8pot_5kb[1]  =  blk93p1i16xx[3] & ~blk93p1i16xx[1] &  ~blk93p1i16xx[0] & xtuu_xtcsg4icbv_;
    assign tmtwlbn11k8pot_5kb[2]  = ~blk93p1i16xx[4] &  blk93p1i16xx[1] &  ~blk93p1i16xx[0] & xtuu_xtcsg4icbv_;
    assign tmtwlbn11k8pot_5kb[3]  =  blk93p1i16xx[4] &  blk93p1i16xx[1] &  ~blk93p1i16xx[0] & xtuu_xtcsg4icbv_;
    assign tmtwlbn11k8pot_5kb[4]  = ~blk93p1i16xx[5] & ~blk93p1i16xx[2] &   blk93p1i16xx[0] & xtuu_xtcsg4icbv_;
    assign tmtwlbn11k8pot_5kb[5]  =  blk93p1i16xx[5] & ~blk93p1i16xx[2] &   blk93p1i16xx[0] & xtuu_xtcsg4icbv_;
    assign tmtwlbn11k8pot_5kb[6]  = ~blk93p1i16xx[6] &  blk93p1i16xx[2] &   blk93p1i16xx[0] & xtuu_xtcsg4icbv_;
    assign tmtwlbn11k8pot_5kb[7]  =  blk93p1i16xx[6] &  blk93p1i16xx[2] &   blk93p1i16xx[0] & xtuu_xtcsg4icbv_;

                          

    assign vs7xk5fv2idvsx3b = ({7{j6u1lgj0jf7udo[0]}} & {blk93p1i16xx[6:4],1'b1,blk93p1i16xx[2],2'b11})
                           | ({7{j6u1lgj0jf7udo[1]}} & {blk93p1i16xx[6:4],1'b0,blk93p1i16xx[2],2'b11})
                           | ({7{j6u1lgj0jf7udo[2]}} & {blk93p1i16xx[6:5],1'b1,blk93p1i16xx[3:2],2'b01})
                           | ({7{j6u1lgj0jf7udo[3]}} & {blk93p1i16xx[6:5],1'b0,blk93p1i16xx[3:2],2'b01})
                           | ({7{j6u1lgj0jf7udo[4]}} & {blk93p1i16xx[6],1'b1,blk93p1i16xx[4:3],1'b1,blk93p1i16xx[1],1'b0})
                           | ({7{j6u1lgj0jf7udo[5]}} & {blk93p1i16xx[6],1'b0,blk93p1i16xx[4:3],1'b1,blk93p1i16xx[1],1'b0})
                           | ({7{j6u1lgj0jf7udo[6]}} & {1'b1,blk93p1i16xx[5:3],1'b0,blk93p1i16xx[1],1'b0})
                           | ({7{j6u1lgj0jf7udo[7]}} & {1'b0,blk93p1i16xx[5:3],1'b0,blk93p1i16xx[1],1'b0})
                           ;
end
else begin:g4j8p5
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   

    assign tmtwlbn11k8pot_5kb[0]  =  ~blk93p1i16xx[1] &  ~blk93p1i16xx[0] & xtuu_xtcsg4icbv_;
    assign tmtwlbn11k8pot_5kb[1]  =   blk93p1i16xx[1] &  ~blk93p1i16xx[0] & xtuu_xtcsg4icbv_;
    assign tmtwlbn11k8pot_5kb[2]  =  ~blk93p1i16xx[2] &   blk93p1i16xx[0] & xtuu_xtcsg4icbv_;
    assign tmtwlbn11k8pot_5kb[3]  =   blk93p1i16xx[2] &   blk93p1i16xx[0] & xtuu_xtcsg4icbv_;

                          

    assign vs7xk5fv2idvsx3b = ({3{j6u1lgj0jf7udo[0]}} & {blk93p1i16xx[2],2'b11})
                           | ({3{j6u1lgj0jf7udo[1]}} & {blk93p1i16xx[2],2'b01})
                           | ({3{j6u1lgj0jf7udo[2]}} & {1'b1,blk93p1i16xx[1],1'b0})
                           | ({3{j6u1lgj0jf7udo[3]}} & {1'b0,blk93p1i16xx[1],1'b0})
                           ;
end
endgenerate

assign j6u1lgj0jf7udo = mv5to8v6 ? {cpuuvz0x4_r5s{1'b0}} : 
                      eqb83t6 ? bnrmlmaiin9wudfye9v7j7   : 
                                i25ll1dii3u_d2n76    ;


wire ou029l35_79b7g0uc00638i = (xtuu_xtcsg4icbv_ & h624jgnv03hp4iysjt03z) | mv5to8v6;
ux607_gnrl_dfflr #(cpuuvz0x4_r5s) paca0uqimbbvs4d0n933f(ou029l35_79b7g0uc00638i,vs7xk5fv2idvsx3b,blk93p1i16xx,gf33atgy,ru_wi); 

wire [cmnocc9r2aiw8za-1:0] dc3tx2ejpweplpq8ck1f27 =  {hw9pzy7xw26mqd67[cmnocc9r2aiw8za-2:0],1'b1} ^ hw9pzy7xw26mqd67;
wire [cmnocc9r2aiw8za-1:0] re7qj5c2go8inyaoucg;

generate
for(i=0;i<cmnocc9r2aiw8za;i=i+1) begin:sxq_amt5geudw_mtdr8g2d41y2
    if(i==0) begin
        assign re7qj5c2go8inyaoucg[i] = dc3tx2ejpweplpq8ck1f27[0];
    end
    else begin
        assign re7qj5c2go8inyaoucg[i] = |dc3tx2ejpweplpq8ck1f27[i:0];
    end
end
endgenerate

wire [cmnocc9r2aiw8za-1:0] ridudot9q3ozuzce_05rf = {re7qj5c2go8inyaoucg[cmnocc9r2aiw8za-2:0],1'b0} ^ re7qj5c2go8inyaoucg;



assign i25ll1dii3u_d2n76 = (xtuu_xtcsg4icbv_ ? tmtwlbn11k8pot_5kb : ridudot9q3ozuzce_05rf);












    wire [b1lh2fnh92-1:0]         sat482scl8zle;
    wire [b1lh2fnh92-1:0]         fdr3d671e7dw6;
    wire                         h8ghyl6u7gffe;
    wire [b1lh2fnh92-1:0]         u99tnldu986760c5;
    wire [b1lh2fnh92-1:0]         y5ramxcxkrqsz12gk;
    wire [b1lh2fnh92-1:0]         frmnwpwxl1k1l;
    wire                         wfoen161d4r42bkqp34lj;
    wire                         hln5byq3t_zxwy8c51dq;
    wire                         klef245vk22hxpmozv2gww9;
    wire                         uoozmjtee2uc_8o;
    wire                         ejae6qevtda080dzd5d;

    assign c2_546oy8pb0vifo = (sat482scl8zle == rqzr_eaa);
    assign uoozmjtee2uc_8o = (sat482scl8zle == eri_rah_b);
    assign ejae6qevtda080dzd5d  = (sat482scl8zle == ib1cruu);

    
    assign wfoen161d4r42bkqp34lj = c2_546oy8pb0vifo & k3n1uuckanw669a & ~es6_9ffb14edb7t;
    assign u99tnldu986760c5 = udqn4evfqnp ? eri_rah_b : ib1cruu;

    
    assign hln5byq3t_zxwy8c51dq = uoozmjtee2uc_8o & (nmlix317bu48vgct7x02m7vgn | es6_9ffb14edb7t);  
    assign y5ramxcxkrqsz12gk = es6_9ffb14edb7t ? rqzr_eaa : ib1cruu;

    
    assign klef245vk22hxpmozv2gww9 = ejae6qevtda080dzd5d;
    assign frmnwpwxl1k1l = es6_9ffb14edb7t ? rqzr_eaa : k3n1uuckanw669a ? (udqn4evfqnp ? eri_rah_b : ib1cruu) : rqzr_eaa;

    assign h8ghyl6u7gffe = wfoen161d4r42bkqp34lj | hln5byq3t_zxwy8c51dq | klef245vk22hxpmozv2gww9;
    assign fdr3d671e7dw6 =    ({b1lh2fnh92{wfoen161d4r42bkqp34lj}} & u99tnldu986760c5)
                            | ({b1lh2fnh92{hln5byq3t_zxwy8c51dq}} & y5ramxcxkrqsz12gk)
                            | ({b1lh2fnh92{klef245vk22hxpmozv2gww9 }} & frmnwpwxl1k1l )
                            ; 

    ux607_gnrl_dfflr #(b1lh2fnh92) afp_kqyn5ft8m (h8ghyl6u7gffe, fdr3d671e7dw6, sat482scl8zle, gf33atgy, ru_wi);




    assign v66ux9ovjkzt3jn   = uoozmjtee2uc_8o & ~es6_9ffb14edb7t;        
    assign cd3lo77nievm4v3    = ayqqbzrthvt93 ? qbo1b11wky6gxke_ : cq30mwyfhqwa;
    assign rgnht1zljy67subvhyua_   = wdmmpqdswy4kjj3h31ammx;
    assign uy22rssg5uc6vyiti9szp = zaab503am_hhz0afn;
    assign h8djzt4zbmppcv2_ai  = whpmltdnnmuxptumq;





    wire               nzo__5h79lmu5x9dbyazy0938h;                      
    wire               ses29jmv82l0e_eww3jzpsb;                      
    wire               ngmbrvnel2lq6mrjp0jyzppp_4;                      
    wire               ipgh1v55v5pp5011n59gpe;                     
    wire               lqbbt_n1cietaa6hc0i47jb;                     

    assign nzo__5h79lmu5x9dbyazy0938h = (ejae6qevtda080dzd5d | c2_546oy8pb0vifo) & k3n1uuckanw669a & ~ba9r7fnn73020zwu2mxj;
    assign ses29jmv82l0e_eww3jzpsb = (s6zb15tq6xjiqgce5nwjcg7be4 & nmlix317bu48vgct7x02m7vgn & ~ayqqbzrthvt93)
                                  ;
    assign ngmbrvnel2lq6mrjp0jyzppp_4 = nzo__5h79lmu5x9dbyazy0938h | ses29jmv82l0e_eww3jzpsb;
    assign ipgh1v55v5pp5011n59gpe = (~nzo__5h79lmu5x9dbyazy0938h) | ses29jmv82l0e_eww3jzpsb;
    ux607_gnrl_dfflr #(1) n3zp7o6x09u_njmw10r (ngmbrvnel2lq6mrjp0jyzppp_4, ipgh1v55v5pp5011n59gpe, lqbbt_n1cietaa6hc0i47jb, gf33atgy, ru_wi);


    wire               adesjoqhoke1n_csw_yxx2xa7h;                      
    wire               u93sq9murty2gxf1w2v9jj8n;                      
    wire               u1mvvdo7j8jptrujwrfabsspc3;                      
    wire               k565bn6i9gvgihmxtnggtjyt85;                     
    wire               nmn9es8_uvn_7f62zzi_vpr;                     

    assign adesjoqhoke1n_csw_yxx2xa7h = (ejae6qevtda080dzd5d | c2_546oy8pb0vifo) & k3n1uuckanw669a & ~ba9r7fnn73020zwu2mxj;
    assign u93sq9murty2gxf1w2v9jj8n = ry0rypry86op3l_hqbwk8pe32ena3e & nmlix317bu48vgct7x02m7vgn & ~ayqqbzrthvt93;
    assign u1mvvdo7j8jptrujwrfabsspc3 = adesjoqhoke1n_csw_yxx2xa7h | u93sq9murty2gxf1w2v9jj8n;
    assign k565bn6i9gvgihmxtnggtjyt85 = (~adesjoqhoke1n_csw_yxx2xa7h) | u93sq9murty2gxf1w2v9jj8n;
    ux607_gnrl_dfflr #(1) nul52ts1l0mwtnxu4jbct8 (u1mvvdo7j8jptrujwrfabsspc3, k565bn6i9gvgihmxtnggtjyt85, nmn9es8_uvn_7f62zzi_vpr, gf33atgy, ru_wi);




    wire               yk4jqd47rvpo13t0dhd_;
    wire               g_2hm45kw1umnxddnda3;
    wire               zo4t1c5t6whg1_p90rbh_;
    wire               sc6nxigf9dbzxk0v_7;
    wire               l7rplj2hf9dlnk_qpyn;
    
    assign yk4jqd47rvpo13t0dhd_ = k3n1uuckanw669a & udqn4evfqnp & ~ba9r7fnn73020zwu2mxj;
    
    assign g_2hm45kw1umnxddnda3 = (k3n1uuckanw669a & eqb83t6 & ~ba9r7fnn73020zwu2mxj) | (nmlix317bu48vgct7x02m7vgn & ~ayqqbzrthvt93);
    assign zo4t1c5t6whg1_p90rbh_ = yk4jqd47rvpo13t0dhd_ | g_2hm45kw1umnxddnda3;
    assign sc6nxigf9dbzxk0v_7 = ~yk4jqd47rvpo13t0dhd_ | g_2hm45kw1umnxddnda3;
    ux607_gnrl_dfflr #(1) y047zq9fspxz7yljr6x72v1 (zo4t1c5t6whg1_p90rbh_, sc6nxigf9dbzxk0v_7, l7rplj2hf9dlnk_qpyn, gf33atgy, ru_wi);

    assign yvy4oon7f_rsa81003k5snsy28 = l7rplj2hf9dlnk_qpyn;
    assign p761bsjfs381j2b7xfn02m8vbu4u  = zmxmooo4wvcx2e65u0o70qz00;
    assign avdv23oy5gvvj_aozmzn5   = th4w08jy003d95gfdsuxyi;
    assign gojz6nraxpmhlx_7ewrhi6di9  = k2iq1fadynzw7wzp0l0;
    assign pxjlub1gdgqvcckianojxej7_mt  = qgxdl96kyqmm_z6_vqw;
    assign ro2z68ba11neqxvjf0uqiz03nt  = ffo1jrw6y2afg69e;
    assign ovl08q5ylus9d7r7ckvnrb0  = fouse5g_ouj8b6we9;
    assign f6o85b68_amv01vbog6ngjt  = u7ojjt008cvz5fxy;
    assign q5guxjr1bjcc5ehbwvbbdz6a__mpjv74z = lqbbt_n1cietaa6hc0i47jb;                             
    assign qkq4xk9dqb1zawk5qa22ux2h35d9lrg = nmn9es8_uvn_7f62zzi_vpr;





    wire               ucbsllt7d9tyc15njkiwhpegs_;                      
    wire               g352qqakre74tm_h4n1sppij7w5;                      
    wire               v95zsr2rei3k5ztke6tdg9ixs7;                      
    wire               vre3k7qwvxmnwss3vzxhey7p;                     
    wire               a1zulvh2tq3r0_lavx8cn;                     

    assign ucbsllt7d9tyc15njkiwhpegs_ = (ejae6qevtda080dzd5d | c2_546oy8pb0vifo) & k3n1uuckanw669a & ba9r7fnn73020zwu2mxj;
    assign g352qqakre74tm_h4n1sppij7w5 = (s6zb15tq6xjiqgce5nwjcg7be4 & nmlix317bu48vgct7x02m7vgn & ayqqbzrthvt93)
                                  ;
    assign v95zsr2rei3k5ztke6tdg9ixs7 = ucbsllt7d9tyc15njkiwhpegs_ | g352qqakre74tm_h4n1sppij7w5;
    assign vre3k7qwvxmnwss3vzxhey7p = (~ucbsllt7d9tyc15njkiwhpegs_) | g352qqakre74tm_h4n1sppij7w5;
    ux607_gnrl_dfflr #(1) mlvm0a__xczmu0w6qc9 (v95zsr2rei3k5ztke6tdg9ixs7, vre3k7qwvxmnwss3vzxhey7p, a1zulvh2tq3r0_lavx8cn, gf33atgy, ru_wi);


    wire               aglad6xjso0b32p8z3whesdla;                      
    wire               xzu4f3fnb505lmb6auc5t9f64;                      
    wire               t8e65ahay1g6z2r0i_lol_4q7t6b;                      
    wire               uu6hbhk64bqs07o3fmb224wpb0m9d;                     
    wire               muetr7m8smfwxsmdyvhgus0cl3;                     

    assign aglad6xjso0b32p8z3whesdla = (ejae6qevtda080dzd5d | c2_546oy8pb0vifo) & k3n1uuckanw669a & ba9r7fnn73020zwu2mxj;
    assign xzu4f3fnb505lmb6auc5t9f64 = ry0rypry86op3l_hqbwk8pe32ena3e & nmlix317bu48vgct7x02m7vgn & ayqqbzrthvt93;
    assign t8e65ahay1g6z2r0i_lol_4q7t6b = aglad6xjso0b32p8z3whesdla | xzu4f3fnb505lmb6auc5t9f64;
    assign uu6hbhk64bqs07o3fmb224wpb0m9d = (~aglad6xjso0b32p8z3whesdla) | xzu4f3fnb505lmb6auc5t9f64;
    ux607_gnrl_dfflr #(1) o782d52smt_m23j8iqiy (t8e65ahay1g6z2r0i_lol_4q7t6b, uu6hbhk64bqs07o3fmb224wpb0m9d, muetr7m8smfwxsmdyvhgus0cl3, gf33atgy, ru_wi);




    wire               guz3xjxid2hcav0hcxkre4;
    wire               s9rtarlwi7eqh6dpj681z;
    wire               k_o_qnnj5p7tj3tldttn;
    wire               rb2_q3e8x_m30zvky;
    wire               jzh0gbz_3czq9s33a01;
    
    assign guz3xjxid2hcav0hcxkre4 = k3n1uuckanw669a & udqn4evfqnp & ba9r7fnn73020zwu2mxj;
    
    assign s9rtarlwi7eqh6dpj681z = (k3n1uuckanw669a & eqb83t6 & ba9r7fnn73020zwu2mxj) | (nmlix317bu48vgct7x02m7vgn & ayqqbzrthvt93);
    assign k_o_qnnj5p7tj3tldttn = guz3xjxid2hcav0hcxkre4 | s9rtarlwi7eqh6dpj681z;
    assign rb2_q3e8x_m30zvky = ~guz3xjxid2hcav0hcxkre4 | s9rtarlwi7eqh6dpj681z;
    ux607_gnrl_dfflr #(1) pqorz_p8xpu5jgq97l9ofg (k_o_qnnj5p7tj3tldttn, rb2_q3e8x_m30zvky, jzh0gbz_3czq9s33a01, gf33atgy, ru_wi);

    assign lrn8i28ncm6vualne3lnezatrmx = jzh0gbz_3czq9s33a01;
    assign d757aw4s0emlk_xndccuz9wrpek3n  = d6ihhd9s3mwhlwqpcw9o0xq;
    assign ky4b1pzcyo6z1omquzzoj   = vneu1upjrxltagmeu7x;
    assign stcauj4mexs59diuva_xf1308li  = yjuujp8x84pgx57z0kn;
    assign v_sj7f9mnvn2sgj37k1ave5g  = dh2xowtqx9d9mq_icq5;
    assign dce56zk48npvti3u7osyzacy  = yqqbs3_6flcq_idm;
    assign dspbo9b1im8onetqwxjnw7  = j5934321vs15d6dj;
    assign kf99vegpc45l_wd1vhgluhfo65  = gx5bpb6ffz6f__05cr;
    assign q0kprornbncukpltocigbw9tba03 = a1zulvh2tq3r0_lavx8cn;                             
    assign w_jjbyn9u5snyb45kcy8r78z6d9iz5 = muetr7m8smfwxsmdyvhgus0cl3;

    assign faamp7iz46_jj1ci8a = uoozmjtee2uc_8o;

endmodule























module kho7cvkwdsu6ed90f6_18aax2 #(
   parameter xio4kx7ep1ojwa_r      = 78,
   parameter cmnocc9r2aiw8za       = 8,
   parameter xholqktr732apzsv8d0  = 3
) (
    input                                    es6_9ffb14edb7t,                
    input                                    mv5to8v6,                       
    
    input                                    zh907qs92c1ixb_97gmdepk,               
    input  [27-1:0]      phofig8d5zd_8v9g8,               
    input  [1:0]                             hey6uxy22wzzlom6mekyg2y,        
    input                                    qerr94cedlotaj08239y,
    input  [26-1:0]    js0ml55dtie8qenb4eoj2,         
    input  [64-1:0]                  ticm3jrqt6tjtf6,              
    input  [64-1:0]                  hpaul9bznamp4qkl,              
    input                                    vq7jwn83uus_ac4s4ghf,                        
    
    input                                    gzh3us4_ux10aey,
    output                                   np3fnkgbpsuf8nkgnf,
    
    
    input                                    evji0n54bi8hm_n24uk853qw9c,               
    input  [27-1:0]      s9psy03yyyxh7qrmosmb1,               
    input  [1:0]                             sqkbogq1h4psprgoosl2lmrpj9_,        
    input                                    n5gj_lxl9078ky9b2zawd0,
    input  [26-1:0]    b0fkq6hghv6az5l_j1j2c12imdd6,         
    input  [64-1:0]                  argq10f3h723e0jtlrdbu53,              
    input  [64-1:0]                  e7iar94ylidlt25a9g9n,              
    input                                    qj6kqe1holct34gfb0q9p9a04_alrzg,                        
    
    input                                    bmkssziw1_8am7ea6dv,
    output                                   xefc2nul9m648jueckdrui_l,

    
    input                                    hpk3eafyque5ubt_c62flnny,        
    input  [27-1:0]      sfezv1xz2ghvo8pkt,               
    input  [1:0]                             vagaza053272juvmo59v8w20s,        
    input                                    rzf45534z36ejq96260,
    input  [26-1:0]    frzfsbt7hp3n4aj3zvvumnh0s,         
    input  [64-1:0]                  zkuxqezrmlhyyjjgx,              
    input  [64-1:0]                  u3h5tvu1g2q93141j9o,              
    input                                    pjh0wad7t_5du3cync_0c,                        
    
    input                                    wmkgrgf631pbq,
    output                                   oyq1p3qa2iffjuqns0jkgg,
    
    
    output                                   c9k79dqw2z4f63_8lcp4w,        
    output [26-1:0]    ly39gmn8_bufgxi162s47mj5md,     
    output [20-1:0]         u6f8hwzstewuo7nl0iywamw,          
    output                                   owio9cfz6lmpk7katn_gtlo9,         
    output                                   dna64e9sa3ona8c40stq,         
    output                                   yqonk7rjhe328d_deg1,         
    output                                   fvuwaqmgv_r72l8z4ys0lq59,         
    output                                   x5_495u23v2cqjqs7nx9m3s,         
    output                                   qvfjqeg7co1udtegoqx2t09jmc,   
    output                                   m6_yvtzjevmj_c4bel_9vu0kkk_t, 

    
    output                                   woq47beoqkpu1um82nv58l1u_hyj4,        
    output [26-1:0]    a1r66jlym5w100htq8lfn_o0rapdf5s,     
    output [20-1:0]         trt0bnwhmoe0r7apy2x_p9hltd,          
    output                                   wqjorkypks0nndgahingvyvil3dvqo,         
    output                                   obokll126527kg6wlw1t6vfh8,         
    output                                   msh4030y2dhqf78kyckys0c2ue0ic,         
    output                                   oebo4piph5o2byr1030bgmb0ye31c6,         
    output                                   tlmtrlht_1gsijvzms1twiewyym,         
    output                                   ez_fxjs3_wlsve__62ua9tqsfa6k89twfir,   
    output                                   p3nsxkqv6seglstz4ge77tdjcngbig0w30rq, 

    
    output                                   qjw2q0j88rjr42lautsqnca,             
    output [26-1:0]    imkm56ujne9v4m6n08w1yf5622,          
    output [20-1:0]         txk1r9aiq_7l2nkw101w_,               
    output                                   ih4hmwugasiodbx5da9_40kx,              
    output                                   x5vjq7mshfwr0h3q514t7mhdt,              
    output                                   qrxtk7e03100_uwkx73sg7,              
    output                                   i7qiq2q9c6hbeful9qu9lb,              
    output                                   yr0s3skqk7cdqflsrbsxg9znu,              
    output                                   adqieke11qo0elfz93hlouwjc0,        
    output                                   w93gdpnnxuydy53eu0s9nxw7xdct7,      

    
    output                                   v66ux9ovjkzt3jn,                
    output  [27-1:0]     cd3lo77nievm4v3,                 
    output  [1:0]                            rgnht1zljy67subvhyua_,          
    output                                   uy22rssg5uc6vyiti9szp,
    output                                   h8djzt4zbmppcv2_ai,
    
    input                                    nmlix317bu48vgct7x02m7vgn,          
    input                                    s6zb15tq6xjiqgce5nwjcg7be4,     
    input                                    ry0rypry86op3l_hqbwk8pe32ena3e,   
    input  [xio4kx7ep1ojwa_r-1:0]              h4zmq2srkdf5iaeagd8d7i87,           
    input                                    dzo70vq3_1_kyxyiurxy1d20ed,         
    input                                    b0c0o6unssb9h3tgqck870,         

    
    output                                   dlygovkaje808pt5_j,                

    
    output                                   c2_546oy8pb0vifo,                 
    input                                    gf33atgy,
    input                                    ru_wi,
    input                                    gc4b3kdcan6do88ta_

);
    wire                                    zn1ks63jnkl4aagnf5ts4ehf; 
    wire  [27-1:0]      lt7tkehfruirbj6stb8ad;
    wire  [1:0]                             vqqsie8bta17asuq1620f3jovdi;
    wire                                    f2wl4y7js12216tnckhdq4qk; 
    wire  [26-1:0]    xzg_tk3qveh7zx8huonb_byrat0k;
    wire  [64-1:0]                  oh96mndsu3cfphpbstk0d3ium; 
    wire  [64-1:0]                  uos9rm9ew98djscgrglaktns;
    wire                                    d57mx4mrtntzzh0eqigojjkjeu;
    wire                                    etn63vnhji57t5oya0fq;
    
    
    
    
    
    
    
    
    
    
    
    
    
    wire                                    rbkv5037v6_ob752blhmqgiaspp;
    wire [26-1:0]     z2wp12c5wlqm2okygg1d0cjllle785;
    wire [20-1:0]          zd199nz1tppq5s3f96i5gs8;
    wire                                    c_yreeadd7fpcjinm5jg9oe;
    wire                                    j856hmn7dn85lwratlc4dk5m;
    wire                                    opis286s9rlfwc1ofmp51q9z3jk;
    wire                                    bkqfcp8pnecu5sgn9_7f_qrgcz;
    wire                                    krwq_tqmkurqot6778_u9r;
    wire                                    a9meb4mfh189f6ja8vgs0186lc5ivx9;
    wire                                    m6xa8a1m1yyfrzyaiiwwu_u71spkil;
    wire                                    dss_r3_bg6s44_cm333fe2f2am;
    wire                                    bnr3veh8i8ec4b_97h5t3c_7gebhn;
    wire                                    uj_wg22_2r4rkzrihrkdd;

    
    
    assign np3fnkgbpsuf8nkgnf       = !dss_r3_bg6s44_cm333fe2f2am && !evji0n54bi8hm_n24uk853qw9c && !hpk3eafyque5ubt_c62flnny;
    assign oyq1p3qa2iffjuqns0jkgg      = !dss_r3_bg6s44_cm333fe2f2am && !evji0n54bi8hm_n24uk853qw9c;
    assign xefc2nul9m648jueckdrui_l = !dss_r3_bg6s44_cm333fe2f2am;

    assign zn1ks63jnkl4aagnf5ts4ehf        = zh907qs92c1ixb_97gmdepk && np3fnkgbpsuf8nkgnf || evji0n54bi8hm_n24uk853qw9c && xefc2nul9m648jueckdrui_l || hpk3eafyque5ubt_c62flnny && oyq1p3qa2iffjuqns0jkgg;
    assign lt7tkehfruirbj6stb8ad        = evji0n54bi8hm_n24uk853qw9c? s9psy03yyyxh7qrmosmb1        : hpk3eafyque5ubt_c62flnny? sfezv1xz2ghvo8pkt        :  phofig8d5zd_8v9g8        ;
    assign vqqsie8bta17asuq1620f3jovdi = evji0n54bi8hm_n24uk853qw9c? sqkbogq1h4psprgoosl2lmrpj9_ : hpk3eafyque5ubt_c62flnny? vagaza053272juvmo59v8w20s :  hey6uxy22wzzlom6mekyg2y ;
    assign f2wl4y7js12216tnckhdq4qk     = evji0n54bi8hm_n24uk853qw9c? n5gj_lxl9078ky9b2zawd0     : hpk3eafyque5ubt_c62flnny? rzf45534z36ejq96260     :  qerr94cedlotaj08239y     ;
    assign xzg_tk3qveh7zx8huonb_byrat0k  = evji0n54bi8hm_n24uk853qw9c? b0fkq6hghv6az5l_j1j2c12imdd6  : hpk3eafyque5ubt_c62flnny? frzfsbt7hp3n4aj3zvvumnh0s  :  js0ml55dtie8qenb4eoj2  ;
    assign oh96mndsu3cfphpbstk0d3ium       = evji0n54bi8hm_n24uk853qw9c? argq10f3h723e0jtlrdbu53       : hpk3eafyque5ubt_c62flnny? zkuxqezrmlhyyjjgx       :  ticm3jrqt6tjtf6       ; 
    assign uos9rm9ew98djscgrglaktns       = evji0n54bi8hm_n24uk853qw9c? e7iar94ylidlt25a9g9n       : hpk3eafyque5ubt_c62flnny? u3h5tvu1g2q93141j9o       :  hpaul9bznamp4qkl       ;
    assign d57mx4mrtntzzh0eqigojjkjeu = evji0n54bi8hm_n24uk853qw9c? qj6kqe1holct34gfb0q9p9a04_alrzg : hpk3eafyque5ubt_c62flnny? pjh0wad7t_5du3cync_0c :  vq7jwn83uus_ac4s4ghf ;
    assign etn63vnhji57t5oya0fq         = evji0n54bi8hm_n24uk853qw9c? bmkssziw1_8am7ea6dv         : hpk3eafyque5ubt_c62flnny? wmkgrgf631pbq         :  gzh3us4_ux10aey         ;
    assign uj_wg22_2r4rkzrihrkdd       = (evji0n54bi8hm_n24uk853qw9c | hpk3eafyque5ubt_c62flnny)   ;
    wire   ni4jijvnr8sd190kgotesti2q4d6a   =  zn1ks63jnkl4aagnf5ts4ehf & uj_wg22_2r4rkzrihrkdd; 
    wire   rxs_xr0gl6z95j50100lmn7lfbbo   = evji0n54bi8hm_n24uk853qw9c;
    ux607_gnrl_dffl #(1) pvjg2spuu_vlcyc7b5qrxos60s9z1 (ni4jijvnr8sd190kgotesti2q4d6a, rxs_xr0gl6z95j50100lmn7lfbbo, bnr3veh8i8ec4b_97h5t3c_7gebhn, gf33atgy, ru_wi);

    
    
    
    
    
    
    
    
    
    
    
    
    
    

    assign woq47beoqkpu1um82nv58l1u_hyj4         =  bnr3veh8i8ec4b_97h5t3c_7gebhn && rbkv5037v6_ob752blhmqgiaspp ;
    assign a1r66jlym5w100htq8lfn_o0rapdf5s      =  z2wp12c5wlqm2okygg1d0cjllle785                  ;
    assign trt0bnwhmoe0r7apy2x_p9hltd           =  zd199nz1tppq5s3f96i5gs8                       ;
    assign wqjorkypks0nndgahingvyvil3dvqo          =  c_yreeadd7fpcjinm5jg9oe                      ;
    assign obokll126527kg6wlw1t6vfh8          =  j856hmn7dn85lwratlc4dk5m                      ;
    assign msh4030y2dhqf78kyckys0c2ue0ic          =  opis286s9rlfwc1ofmp51q9z3jk                      ;
    assign oebo4piph5o2byr1030bgmb0ye31c6          =  bkqfcp8pnecu5sgn9_7f_qrgcz                      ;
    assign tlmtrlht_1gsijvzms1twiewyym          =  krwq_tqmkurqot6778_u9r                      ;
    assign ez_fxjs3_wlsve__62ua9tqsfa6k89twfir    =  a9meb4mfh189f6ja8vgs0186lc5ivx9                ;
    assign p3nsxkqv6seglstz4ge77tdjcngbig0w30rq  =  m6xa8a1m1yyfrzyaiiwwu_u71spkil              ;

    assign qjw2q0j88rjr42lautsqnca         =  !bnr3veh8i8ec4b_97h5t3c_7gebhn && rbkv5037v6_ob752blhmqgiaspp ;
    assign imkm56ujne9v4m6n08w1yf5622      =  z2wp12c5wlqm2okygg1d0cjllle785                  ;
    assign txk1r9aiq_7l2nkw101w_           =  zd199nz1tppq5s3f96i5gs8                       ;
    assign ih4hmwugasiodbx5da9_40kx          =  c_yreeadd7fpcjinm5jg9oe                      ;
    assign x5vjq7mshfwr0h3q514t7mhdt          =  j856hmn7dn85lwratlc4dk5m                      ;
    assign qrxtk7e03100_uwkx73sg7          =  opis286s9rlfwc1ofmp51q9z3jk                      ;
    assign i7qiq2q9c6hbeful9qu9lb          =  bkqfcp8pnecu5sgn9_7f_qrgcz                      ;
    assign yr0s3skqk7cdqflsrbsxg9znu          =  krwq_tqmkurqot6778_u9r                      ;
    assign adqieke11qo0elfz93hlouwjc0    =  a9meb4mfh189f6ja8vgs0186lc5ivx9                ;
    assign w93gdpnnxuydy53eu0s9nxw7xdct7  =  m6xa8a1m1yyfrzyaiiwwu_u71spkil              ;

    
    wire p5q87c1_052rxw0fd;
    ux607_gnrl_dffr #(1) o2hkz4toqzq9567pgsr (es6_9ffb14edb7t, p5q87c1_052rxw0fd, gf33atgy, ru_wi);

    assign dlygovkaje808pt5_j = dss_r3_bg6s44_cm333fe2f2am;

    rrxf4gi2j6 #(
       .xio4kx7ep1ojwa_r     (xio4kx7ep1ojwa_r    ),
       .cmnocc9r2aiw8za      (cmnocc9r2aiw8za     ),
       .xholqktr732apzsv8d0 (xholqktr732apzsv8d0)
    ) qp7tor58p55 (
       .es6_9ffb14edb7t                     (es6_9ffb14edb7t                  ),   
       .mv5to8v6                          (mv5to8v6                       ),                       
       .ba9r7fnn73020zwu2mxj                 (uj_wg22_2r4rkzrihrkdd          ),   
       .k3n1uuckanw669a                  (zn1ks63jnkl4aagnf5ts4ehf           ),               
       .qfy7pr76nvqld1f                  (lt7tkehfruirbj6stb8ad           ),               
       .nowfs1y75z9hmhv6r0ppp6vjly           (vqqsie8bta17asuq1620f3jovdi    ),               
       .xtm2ue4np_4lj4a7ik               (f2wl4y7js12216tnckhdq4qk        ),               
       .fsxy2ey9lgj3xvg2hw_sqfrgy            (xzg_tk3qveh7zx8huonb_byrat0k     ),         
       .h5arfbj2deloqqwtp1                 (oh96mndsu3cfphpbstk0d3ium          ),              
       .elgnxkek04s_nuz6z                 (uos9rm9ew98djscgrglaktns          ),              
       .gcoematpqzttdb81ozfq3zg1v9           (d57mx4mrtntzzh0eqigojjkjeu    ),        
       .a9q83azb3dode6qt                   (etn63vnhji57t5oya0fq            ),
       .yvy4oon7f_rsa81003k5snsy28          (c9k79dqw2z4f63_8lcp4w          ),        
       .p761bsjfs381j2b7xfn02m8vbu4u       (ly39gmn8_bufgxi162s47mj5md       ),     
       .avdv23oy5gvvj_aozmzn5            (u6f8hwzstewuo7nl0iywamw            ),          
       .gojz6nraxpmhlx_7ewrhi6di9           (owio9cfz6lmpk7katn_gtlo9           ),         
       .pxjlub1gdgqvcckianojxej7_mt           (dna64e9sa3ona8c40stq           ),         
       .ro2z68ba11neqxvjf0uqiz03nt           (yqonk7rjhe328d_deg1           ),         
       .ovl08q5ylus9d7r7ckvnrb0           (fvuwaqmgv_r72l8z4ys0lq59           ),         
       .f6o85b68_amv01vbog6ngjt           (x5_495u23v2cqjqs7nx9m3s           ),         
       .q5guxjr1bjcc5ehbwvbbdz6a__mpjv74z     (qvfjqeg7co1udtegoqx2t09jmc     ),   
       .qkq4xk9dqb1zawk5qa22ux2h35d9lrg   (m6_yvtzjevmj_c4bel_9vu0kkk_t   ), 
       .lrn8i28ncm6vualne3lnezatrmx          (rbkv5037v6_ob752blhmqgiaspp       ),        
       .d757aw4s0emlk_xndccuz9wrpek3n       (z2wp12c5wlqm2okygg1d0cjllle785    ),     
       .ky4b1pzcyo6z1omquzzoj            (zd199nz1tppq5s3f96i5gs8         ),          
       .stcauj4mexs59diuva_xf1308li           (c_yreeadd7fpcjinm5jg9oe        ),         
       .v_sj7f9mnvn2sgj37k1ave5g           (j856hmn7dn85lwratlc4dk5m        ),         
       .dce56zk48npvti3u7osyzacy           (opis286s9rlfwc1ofmp51q9z3jk        ),         
       .dspbo9b1im8onetqwxjnw7           (bkqfcp8pnecu5sgn9_7f_qrgcz        ),         
       .kf99vegpc45l_wd1vhgluhfo65           (krwq_tqmkurqot6778_u9r        ),         
       .q0kprornbncukpltocigbw9tba03     (a9meb4mfh189f6ja8vgs0186lc5ivx9  ),   
       .w_jjbyn9u5snyb45kcy8r78z6d9iz5   (m6xa8a1m1yyfrzyaiiwwu_u71spkil), 

       .faamp7iz46_jj1ci8a                (dss_r3_bg6s44_cm333fe2f2am        ),             
       .v66ux9ovjkzt3jn                   (v66ux9ovjkzt3jn               ),                
       .cd3lo77nievm4v3                    (cd3lo77nievm4v3                ),                 
       .rgnht1zljy67subvhyua_             (rgnht1zljy67subvhyua_         ),                 
       .uy22rssg5uc6vyiti9szp                 (uy22rssg5uc6vyiti9szp             ),                 
       .h8djzt4zbmppcv2_ai                  (h8djzt4zbmppcv2_ai              ),
       .nmlix317bu48vgct7x02m7vgn             (nmlix317bu48vgct7x02m7vgn         ),          
       .s6zb15tq6xjiqgce5nwjcg7be4        (s6zb15tq6xjiqgce5nwjcg7be4    ),     
       .ry0rypry86op3l_hqbwk8pe32ena3e      (ry0rypry86op3l_hqbwk8pe32ena3e  ),   
       .h4zmq2srkdf5iaeagd8d7i87              (h4zmq2srkdf5iaeagd8d7i87          ),           
       .dzo70vq3_1_kyxyiurxy1d20ed            (dzo70vq3_1_kyxyiurxy1d20ed        ),         
       .b0c0o6unssb9h3tgqck870            (b0c0o6unssb9h3tgqck870        ),         
       .c2_546oy8pb0vifo                  (c2_546oy8pb0vifo              ),               
       .gf33atgy                              (gf33atgy                          ),
       .ru_wi                            (ru_wi                        ),
       .gc4b3kdcan6do88ta_                   (gc4b3kdcan6do88ta_               )
    );
    
endmodule 





















module cqpjxz2qb247thego6htwvkw_aiu (
  
  input                                   f_8ecse5wf0jrndlozy2070bja,        
  input [26-1:0]    e4sprh35cvfb6sw6lnskyaga91,
  input                                   qrvtg_49_dmoggu94orq0,         
  input                                   iocew24g1qos_gvi3_r3uoqfdf,         
  input                                   qh_y92pv7dp1us9t5wxdmm57,         
  input                                   cznjry8adajzgi6gkmyr830m_u,         
  input                                   ugixcggahb26m1glzpuqvpq,         
  input                                   vbpz6tidsg3o93kih6nmamlyg9wmr1zz,   
  input                                   j2dtuvq0m4iir947lery9tpxqwhjj2g3, 
  
  input                                   wzqcq7ug3_gv3tuf0o,
  
  input                                   ng5gq72xr47fw8fztwfo8hw, 
  input [1:0]                             cmyy3ooatm0bn2s6fv8_r, 
  input                                   ckgybqpbvuzwgxv1ixd_6rpf,
  input                                   nguthky_k_yqsf8fa9btry1,
  input [1:0]                             w30ye15yns15,
  input                                   jyl_xsaj6z1u9wndwpi,
  input                                   idg19n7mm21jtb,
  
  output                                  o_4mw1alrjmdzl,
  output                                  nkjxsm02z2_q5_0_,
  
  input     gf33atgy,
  input     ru_wi
);
  wire       r541xuss17h9n9b; 
  wire       uhp_6lt6thhcwq; 
  wire       jyfluwl_ll; 
  wire       ouumoo1sk096;
  wire       qwbsekhtca5zlfo9x;
  wire       s5nurokljqe_w91_yp;
  wire       kmwjyiszj2ya;
  wire       sout20o1pphwqv;
  wire       s9_82_tp66v;

  assign kmwjyiszj2ya      =   (ckgybqpbvuzwgxv1ixd_6rpf && qrvtg_49_dmoggu94orq0)
                         ||  iocew24g1qos_gvi3_r3uoqfdf
                         ;
  assign sout20o1pphwqv     =  ((w30ye15yns15 == 2'b00)                                                           && !idg19n7mm21jtb)          
                         ||((w30ye15yns15 == 2'b11) && ng5gq72xr47fw8fztwfo8hw && (cmyy3ooatm0bn2s6fv8_r == 2'b00) && !idg19n7mm21jtb)          
                         ||((w30ye15yns15 == 2'b11) && ng5gq72xr47fw8fztwfo8hw && (cmyy3ooatm0bn2s6fv8_r == 2'b00) && !idg19n7mm21jtb)          
                         ||(idg19n7mm21jtb && jyl_xsaj6z1u9wndwpi && ng5gq72xr47fw8fztwfo8hw && (cmyy3ooatm0bn2s6fv8_r == 2'b00))                
                         ;
  assign s9_82_tp66v     =  ((w30ye15yns15 == 2'b01)                                                           && !idg19n7mm21jtb)          
                         ||((w30ye15yns15 == 2'b11) && ng5gq72xr47fw8fztwfo8hw && (cmyy3ooatm0bn2s6fv8_r == 2'b01) && !idg19n7mm21jtb)          
                         ||(idg19n7mm21jtb && jyl_xsaj6z1u9wndwpi && ng5gq72xr47fw8fztwfo8hw && (cmyy3ooatm0bn2s6fv8_r == 2'b01))                
                         ;
  assign s5nurokljqe_w91_yp =   (e4sprh35cvfb6sw6lnskyaga91 != {26{1'b1}})
                         && (e4sprh35cvfb6sw6lnskyaga91 != {26{1'b0}})
                         ;
  assign r541xuss17h9n9b     = !wzqcq7ug3_gv3tuf0o && !kmwjyiszj2ya && (sout20o1pphwqv || s9_82_tp66v);
  assign uhp_6lt6thhcwq     =  wzqcq7ug3_gv3tuf0o && !cznjry8adajzgi6gkmyr830m_u && (sout20o1pphwqv || s9_82_tp66v);
  assign jyfluwl_ll     =  wzqcq7ug3_gv3tuf0o && !qh_y92pv7dp1us9t5wxdmm57 && (sout20o1pphwqv || s9_82_tp66v);
  assign ouumoo1sk096   =  sout20o1pphwqv         && !ugixcggahb26m1glzpuqvpq;
  assign qwbsekhtca5zlfo9x   =  s9_82_tp66v         &&  ugixcggahb26m1glzpuqvpq && !nguthky_k_yqsf8fa9btry1;

  assign nkjxsm02z2_q5_0_ = f_8ecse5wf0jrndlozy2070bja && j2dtuvq0m4iir947lery9tpxqwhjj2g3;
  
  wire j0qe7qal7faiwm5se = j2dtuvq0m4iir947lery9tpxqwhjj2g3
                          ;

  assign o_4mw1alrjmdzl   = f_8ecse5wf0jrndlozy2070bja && 
                         (vbpz6tidsg3o93kih6nmamlyg9wmr1zz           ||
                          r541xuss17h9n9b   && !j0qe7qal7faiwm5se    ||
                          uhp_6lt6thhcwq   && !j0qe7qal7faiwm5se    ||
                          jyfluwl_ll   && !j0qe7qal7faiwm5se    ||
                          ouumoo1sk096 && !j0qe7qal7faiwm5se    ||
                          qwbsekhtca5zlfo9x && !j0qe7qal7faiwm5se    ||
                          s5nurokljqe_w91_yp)
                          ;

endmodule






















module xqy0kx72ozzh4s06ej(

  input sxvvsxtbhyvt,

  
  
  
  
  
  
  
  
  
  

  input                        rm1dxjejhq7dh3q5m,
  input                        rvr30vvllni,
  output                       oa95jvzldxkjxnka5,
  output [32-1:0]   hjbzyjew4g2fmth4l66ng8,
  output                       dl59edtk0_9k5jd65gxp,
  output                       unzbnfwje52jxr_9yt38_bmn,
  output                       qtcuhd18j5hjtx41o9tjmv0cm434,
  output                       srphqbnx3w67orxkuwvoz,
  output                       jbju6a9hecf_f8kg2bsz4,
  input                        w66c528fqa9qnfz1btjnm,

  
  
  
  
  input                        badsf4ksbp3k6p_p5hnj2i,
  output                       ed4kcy8s9nrisftgx_q,
  input                        xhpc6eofokpbnya1h3s117_2,
  input  [32-1:0]   bdqo1tgw2_bpi2e8alini, 
  input                        jp5nha2l14e7kx2jzpke, 
  input  [64-1:0]    a4a48egkdkec8d9b_9, 
  input  [8-1:0]    xwfmltfzahuj4qfn4qf2, 
  input  [1:0]                 ggxoqcj7ytp1a4pjf7ee,
  input  [4-1:0]oq9b5zfhza9yvdoj,
  input                        l3c127qdc9a2mfc13,
  input                        zdpamqgv7ddf1n3x5t2q,
  input                        wpsukhyqhl92dzoam7cm,
  input                        v3oo69y614hgiemyyld,
  input                        vy1zc0f0lrbzkonj3v,
  input                        uxlldm0w_h7kicit8gvhqv2,
  input                        yvu98r_7ji4o250r_u, 
  input                        o21b8ypt1xiu5ml63d,

  input      l_giy79jkzkxy7j  ,
  input      cw9xa748nw    ,
  input      x1huhi29x9mco   ,

  input      fpo04urqz74     ,
  input      a2i6e7_7    ,
  input      cque110xwd150_ ,
  input      m705cbtazx7y  ,
  input      etp831o_vh94  ,
  input      w3p1po3pu   ,
  input      nxy2oljfg0lssc  ,
  input      n2s7mr_zvl9k  ,
  input      mzwwsw0h6m1  ,
  input      lydg_n0cr655 ,
  input      tb62wswspbytv ,
  input  [64-1:0]      jttn_e63nm4n4lm9, 

  input      jgah5jfw    ,

  
  input  [1:0]                st2zalpx0uf, 
  input                       ni01kj42oob2x, 
  input                       ah8kjlmvnaxzbi, 
  input  [1:0]                w30ye15yns15,
  
  input                        vdtkg4_jnsbu0p8wqnasmncdouhwmk,
  input  [64-1:0] wqbvx_uqjrfzj8cjke712tpq, 
  input                        dll7vburbug9zho0oh3rpr0pnjnnh,
  
  
  output                                  evji0n54bi8hm_n24uk853qw9c,               
  output  [27-1:0]    s9psy03yyyxh7qrmosmb1,               
  output  [1:0]                           sqkbogq1h4psprgoosl2lmrpj9_,        
  output                                  n5gj_lxl9078ky9b2zawd0,                        
  output  [26-1:0]  b0fkq6hghv6az5l_j1j2c12imdd6,         
  output  [64-1:0]                argq10f3h723e0jtlrdbu53,              
  output  [64-1:0]                e7iar94ylidlt25a9g9n,              
  output                                  qj6kqe1holct34gfb0q9p9a04_alrzg,                        
  
  output                                  bmkssziw1_8am7ea6dv,
  input                                   xefc2nul9m648jueckdrui_l,
  
  input                                   woq47beoqkpu1um82nv58l1u_hyj4,       
  input [26-1:0]    a1r66jlym5w100htq8lfn_o0rapdf5s,    
  input [20-1:0]         trt0bnwhmoe0r7apy2x_p9hltd,         
  input                                   wqjorkypks0nndgahingvyvil3dvqo,        
  input                                   obokll126527kg6wlw1t6vfh8,        
  input                                   msh4030y2dhqf78kyckys0c2ue0ic,        
  input                                   oebo4piph5o2byr1030bgmb0ye31c6,        
  input                                   tlmtrlht_1gsijvzms1twiewyym,        
  input                                   ez_fxjs3_wlsve__62ua9tqsfa6k89twfir,  
  input                                   p3nsxkqv6seglstz4ge77tdjcngbig0w30rq,


  output     xmbe_e4vm6ofjbn7lq ,


  
  
  
  
  output                       aht5xalx865dt9ymg6t4,
  input                        zjmbnwsbyle24ayly67,
  output [32-1:0]   icfwo5l56zab795f, 
  output                       n78yvkhg0miifi58, 
  output [64-1:0]    wu02k99r_ok2kjj4u119us, 
  output [8-1:0]    ccwk4o03vlem_hqcccf1g6, 
  output                       yx2bhxvyxmxjggxrsrr833, 
  output                       qe64ftxd03f_vqrd2sd,
  output                       b36sriu021vdo_ujif8,
  output [1:0]                 ltx9lurd9p2ivmnufrgrw,
  output [4-1:0]o1gawztvzi0onzitk,
  output                       lr02cqs6anj9gvr45kv,
  output                       z6ncd60zcel8m99zg6v,
  output                       st9_is6howar7iysonyyhk,
  output                       o8407eu9fhzcuymr2a4,
  output                       t3ubula_wguy1a2tut1_e,
  output                       ukl6eat4ng6xala4y597l2i,
  output                       w3yoivbzacxwr95dw,
  output                       qsw59ks9jxcsmmh,

  
  input                        s4dz24kz7cxir4hxtt,
  output                       epoc75xqnuvcqziu_9i55h,
  input                        w0vagcfu1v7wkym9f  ,
  input                        sjx2nupt4_7eb6_metse,
  input  [64-1:0]    gxo5tf4bea2gsq4yyn,

  
  
  
  output                         jugi02ecegnos3, 
  input                          rxjuugktc38un, 
  output [64-1:0]        h8wu7unf_ixmxfeh, 
  output [4 -1:0] kdpgigzs75vcc1d,
  output                         coohnlu_ri , 
  output                         x6uy7s6mcepqq2j527jtxk, 
  output                         igo49dpz9ealh4h13a, 
  output                         ks33bi5hojtg0te9bl7, 
  output [64 -1:0]  dwet7q3ucodidho7qxlw,
  output [64   -1:0]  p_p6yt19xmgqbfsn0y,
  output                         k5h5ux92dlz_nn0,
  output                         e6uinbhqc8o7iylg7d,

  output j2_lz0mpsxf4xotgqf1ngx,
  output hcugdkhp9szims1nk8rhakn,
  output dw2ygdedledlm7ps830qgbwonu,

  output ygvgcd3cyi2ipiz53hbsp,

  input  gf33atgy,
  input  ru_wi
  );

  
  wire jrhs989pgz0z8or09 = aht5xalx865dt9ymg6t4 & zjmbnwsbyle24ayly67;
  wire b5b1bdkf9u8xkel6mtmr = s4dz24kz7cxir4hxtt & epoc75xqnuvcqziu_9i55h;
  wire wh1vvvsvv8tc2elyruo93 = badsf4ksbp3k6p_p5hnj2i & ed4kcy8s9nrisftgx_q;
  wire                            csz9svan7w77t2lrv3uyj__;
  wire                            hklxc4qx7d75xvdr5e3x9;
  wire                            d34m6fs9h9d3zali7nxf8ogkumrusqb; 
  wire                            eht8nc5zc5sdbpe9nqr67jeju;
  wire                            f8ouikbgg2hqwm8g;
  wire                            dvqdxyi_ja1x2; 
  wire                            chhrgp_9_w35oxb; 
  wire                            eub1wmkjoekn;
  wire [20-1:0]  ikiluasjdq;

  wire wfoen161d4r42bkqp34lj;

  wire jsrfd8uzrbk =   wfoen161d4r42bkqp34lj;


  wire qndyhstqm8pvl   ;
  wire qj_5hjk5ts  ;
  wire qhbdaf2fmdi6ba ;
  wire y0nv37yd84l    ;
  wire ai2cjirv   ;
  wire euomkrkdp_x2p16;
  wire qdiehi55s8izv5y ;
  wire hksju1a__h21 ;
  wire yod75j20uh  ;
  wire v_zd2akdl84 ;
  wire u1npc4m1kjg ;
  wire ybfhwehnrx61b8 ;
  wire ed7pawk0e32us153;
  wire gg2d7pi35s036m89;

  wire encgymm9xrq0    ;

  wire [8-1:0]   x90uy0klprtqdcq;
  wire [64-1:0]      m6uirg1k2s6vd_m8; 
  wire [64-1:0]      fn5e7uint162p6axap1i1t9; 
  wire [64-1:0]      i200dby;
  wire [64-1:0]      trgbsbj;

  wire  [1:0]                 t6rn2o8trm4jaor9u9i2  ;
  wire  [4-1:0]adng7z_1b3srxoxai1rm  ;
  wire                        deonbdggc2hhsqq88 ;
  wire                        av4ep8dz4xawf95kyr8j ;
  wire                        jomllj1p1gxavhm9n ;
  wire                        ynqlvklp9ljiaqdpo ;
  wire                        pf428il3xdc1fkqtfv706k;
  wire                        fjk5178vaf1h3l5q9_p;
  wire                        zelwmbvyieb_h56;

  wire iy42niqez8r3zkja;

  
  assign d34m6fs9h9d3zali7nxf8ogkumrusqb = bdqo1tgw2_bpi2e8alini[12]; 
  assign eub1wmkjoekn = woq47beoqkpu1um82nv58l1u_hyj4;
  ux607_gnrl_dfflr #(1) wsx8rptuz8iyk6fgyl3g    (jsrfd8uzrbk, d34m6fs9h9d3zali7nxf8ogkumrusqb   , dvqdxyi_ja1x2   , gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1) tcq5mbpnrhb6kzt2cvlkssp_q  (jsrfd8uzrbk, vdtkg4_jnsbu0p8wqnasmncdouhwmk  , f8ouikbgg2hqwm8g  , gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1) t60u_0c7cp_57ro5xi04luqq  (jsrfd8uzrbk, dll7vburbug9zho0oh3rpr0pnjnnh  , chhrgp_9_w35oxb  , gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(20) ibsy8l1yu6may (eub1wmkjoekn, trt0bnwhmoe0r7apy2x_p9hltd, ikiluasjdq, gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1) z1qfjjaszmb2783w    (jsrfd8uzrbk, cw9xa748nw   , qndyhstqm8pvl   , gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1) gzwa10p9yk65rh71yx6f   (jsrfd8uzrbk, x1huhi29x9mco  , qj_5hjk5ts  , gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1) wo83l2v4t1v07ry1zo3s6  (jsrfd8uzrbk, l_giy79jkzkxy7j , qhbdaf2fmdi6ba , gf33atgy, ru_wi);  
  ux607_gnrl_dfflr #(1) md1ifh3d8py1h56     (jsrfd8uzrbk, fpo04urqz74    , y0nv37yd84l    , gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1) dy5ak0hpmcgvgi0r_v    (jsrfd8uzrbk, a2i6e7_7   , ai2cjirv   , gf33atgy, ru_wi); 
  ux607_gnrl_dfflr #(1) sks7bnt1aj6vx9933i_sdq (jsrfd8uzrbk, cque110xwd150_, euomkrkdp_x2p16, gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1) pdlhgmq0g7btxa0bhwrd4  (jsrfd8uzrbk, m705cbtazx7y , qdiehi55s8izv5y , gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1) e4qa_0k8y_7u6sopmxktt  (jsrfd8uzrbk, etp831o_vh94 , hksju1a__h21 , gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1) ekms38r37uyeado   (jsrfd8uzrbk, w3p1po3pu  , yod75j20uh  , gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1) fmz_bmvjqfw8ucwwh9pl  (jsrfd8uzrbk, nxy2oljfg0lssc , v_zd2akdl84 , gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1) n_fu9g6owj0qv0kzao1  (jsrfd8uzrbk, n2s7mr_zvl9k , u1npc4m1kjg , gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1) gmv83k9yaz5_zpmyskv1u  (jsrfd8uzrbk, mzwwsw0h6m1 , ybfhwehnrx61b8 , gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1) y5sl7wkq6r_wxs0q8gw (jsrfd8uzrbk, lydg_n0cr655, ed7pawk0e32us153, gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1) x3hfzwaxvt0aacrevbvn28 (jsrfd8uzrbk, tb62wswspbytv, gg2d7pi35s036m89, gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(64) izhiohxizdwojpabgz (jsrfd8uzrbk, jttn_e63nm4n4lm9, i200dby, gf33atgy, ru_wi);

  ux607_gnrl_dfflr #(1) j449e15lx5c_bho     (jsrfd8uzrbk, jgah5jfw    , encgymm9xrq0    , gf33atgy, ru_wi);

  assign trgbsbj = 64'b0;

  ux607_gnrl_dfflr #(2)                zl8aommdo7h602bjqoinwun5   (jsrfd8uzrbk, ggxoqcj7ytp1a4pjf7ee  , t6rn2o8trm4jaor9u9i2  , gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(4) lwg1fzfftyxh5o8bdm0o1i9i   (jsrfd8uzrbk, oq9b5zfhza9yvdoj  , adng7z_1b3srxoxai1rm  , gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1)                ho3dhs8lfbhe8fqmea38o6em1f  (jsrfd8uzrbk, l3c127qdc9a2mfc13 , deonbdggc2hhsqq88 , gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1)                gbxjtu8vxe9taovdwcvo2wsl7cfh  (jsrfd8uzrbk, zdpamqgv7ddf1n3x5t2q , av4ep8dz4xawf95kyr8j , gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1)                ukaaags0cf1ocz_h_9l2ofgkj  (jsrfd8uzrbk, wpsukhyqhl92dzoam7cm , jomllj1p1gxavhm9n , gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1)                a1pl79t6s9oyybwmlwyphuutdb  (jsrfd8uzrbk, v3oo69y614hgiemyyld , ynqlvklp9ljiaqdpo , gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1)                rx4tekg7wpcv2tkaspi588ju (jsrfd8uzrbk, vy1zc0f0lrbzkonj3v, pf428il3xdc1fkqtfv706k, gf33atgy, ru_wi);
  
  
  
  

  ux607_gnrl_dfflr #(1) xporzza3a2f8nolqrdfws7 (jsrfd8uzrbk, rvr30vvllni, iy42niqez8r3zkja, gf33atgy, ru_wi);


  wire gqljc8mgip  = (t6rn2o8trm4jaor9u9i2 == 2'b00);
  wire glc7xaf_upxku  = (t6rn2o8trm4jaor9u9i2 == 2'b01);
  wire d74326txgko0  = (t6rn2o8trm4jaor9u9i2 == 2'b10);
  wire cfe949_7aiw  = (t6rn2o8trm4jaor9u9i2 == 2'b11);

  wire lgf34_8i5f2254 = (l_giy79jkzkxy7j & cw9xa748nw) ;
  wire u9y07o_n2vgf1zk = (l_giy79jkzkxy7j & x1huhi29x9mco) ;
  wire ldn2go4l40668ayimy = (lgf34_8i5f2254 | u9y07o_n2vgf1zk);
 
  wire ijk5d1s_9m5n = (qhbdaf2fmdi6ba & qndyhstqm8pvl) ;
  wire qxeco0b4xvxw1v = (qhbdaf2fmdi6ba & qj_5hjk5ts) ;
  wire lgnnlckl1qq6psb = (ijk5d1s_9m5n | qxeco0b4xvxw1v);

  wire lkrl_gk1f715er9ueo;

     
  wire [64-1:0] tp6hfcjxcyp899mpksjl;
  wire [64-1:0] f4ds8dbk9kk_ic_;
  wire oso3fj0gx6pnvjni;
  wire xl9r7gr7wciuv2d00b ;
  wire htcsb0affil7c6q ;
  wire vrqdq7uwxf99gj_7  ;
  wire jqgtsdtxss_uios07 ;
  wire hn2h_gkqinydwsdg_i3 ;
  wire re8hncw6m47hrh6 ;
  wire tshku7fgpiu2j7ugwjj9;
  wire arc8ztjel_qlz3xfw0ya;
  wire dukom1hk2mc9i6m4;
  wire [64-1:0] ttgsydregi0kgoj_z;

     
  wire e__67e1k5hdb4ctnr;
  wire [64-1:0] jay_5c6ndpwhj0vqzv;
  wire [64-1:0] kn6tx97_rw9w0v;

  wire nc_3q2q5fz4e2;
  wire [64-1:0] a5y809wbv8w1d0;
  wire [64-1:0] l0vxn4vg6wd;










  localparam fnk0axwxfk4kr8z = 6;

  wire gsoquod_6th_uva;
  wire [fnk0axwxfk4kr8z-1:0] brgdc0amsvlnwf_2j;
  wire [fnk0axwxfk4kr8z-1:0] rc887zv55nqt;

  
  localparam i3mg661fq9njsp5b = 6'd0;
  
  localparam v_qy6klyvlpd9v  = 6'd1 + 6'd32;
  
  localparam elevjtxw8s86z  = 6'd2 + 6'd32;
  
  
  localparam r10y29zxz4oiu3wd  = 6'd3 + 6'd32;
  
  localparam w7jie_pve8zo265khr8  = 6'd4 + 6'd32;
  
  localparam zj40kikmdbcd575xl7lmss  = 6'd5 + 6'd32;
  
  localparam fvtdvg067g05k  = 6'd6 + 6'd32;
  
  localparam m9bvbk39_2zfrkcpc  = 6'd7 + 6'd32;
  
  localparam sr0ftn45dhialfn  = 6'd8 + 6'd32;
  
  localparam d0ga83_71diabio74osj0  = 6'd9 + 6'd32;
  
  localparam p0veyq__3ajbausg2h  = 6'd10 + 6'd32;
  
  localparam x8jj4nrwgh_5270b_ftdv0  = 6'd11 + 6'd32;
  
  localparam saah2jpqh8i05  = 6'd12 + 6'd32;
  
  localparam gippr9ch9ni48cz3e47n  = 6'd13 + 6'd32;
  
  localparam zqlr7fq_zdgau_fa1r  = 6'd14 + 6'd32;
  
  localparam ar4t4ajioitfe1gtru35r  = 6'd15 + 6'd32;
  
  localparam eusn96ps48lsd4p  = 6'd16 + 6'd32;
  localparam zjl6he1ayeuql_m_f    = 6'd17 + 6'd32;
  localparam m3aw6280mg3tu3ht0567 = 6'd18 + 6'd32;
  localparam h_kmmziwjubh_5825       = 6'd19 + 6'd32;
  
   
  
 
  wire [fnk0axwxfk4kr8z-1:0] u99tnldu986760c5   ;
  wire [fnk0axwxfk4kr8z-1:0] g9natvym5lqakd    ;
  wire [fnk0axwxfk4kr8z-1:0] qyw9w17wm01o0ibqri8;
  wire [fnk0axwxfk4kr8z-1:0] evn7vmlv0q87c    ;
  wire [fnk0axwxfk4kr8z-1:0] gyiivu76k6m_fi   ;
  wire [fnk0axwxfk4kr8z-1:0] w9wl5ox_pnuvzp     ;
  wire [fnk0axwxfk4kr8z-1:0] zu_l0qkgxjl8mlhw ;
  wire [fnk0axwxfk4kr8z-1:0] lzbc5hwhr2m0yxt  ; 
  wire [fnk0axwxfk4kr8z-1:0] etqkl_z3d5k_z3n1fr;
  wire [fnk0axwxfk4kr8z-1:0] yqwi1z4q7s0wriam8    ;
  wire [fnk0axwxfk4kr8z-1:0] g897ues2orwmfihybd;
  wire [fnk0axwxfk4kr8z-1:0] skmlitjb4kdramm    ;
  wire [fnk0axwxfk4kr8z-1:0] uv3o5o9wdyyhfp16ijtnst;
  wire [fnk0axwxfk4kr8z-1:0] c9v_t190cck33l9    ;
  wire [fnk0axwxfk4kr8z-1:0] anh_5y93ex8mfy8zqs4h;
  wire [fnk0axwxfk4kr8z-1:0] i41gux5i8cqjqp    ;
  wire [fnk0axwxfk4kr8z-1:0] v_nz7nezxqthl8mkc;
  wire [fnk0axwxfk4kr8z-1:0] dxqq9l9bv3v20jsdv    ;
  wire [fnk0axwxfk4kr8z-1:0] h5chs70629xcwrlur;
  wire [fnk0axwxfk4kr8z-1:0] auqrmggnbde5eb    ;

  wire oz66a4n0vakndgbkbj6ds      ;
  wire odvuoxdd_64egspdavi73jis74  ;
  wire z5xqhvuiqp_g510lj8      ;
  wire j98f_s869qm5bv_dhgbcim3     ;
  wire wtgeux804w78dcd92swmjz7a5    ;
  wire uwnli3a8y85_7gsqwb41d_   ;
  wire d2jegnujjeil20nht       ;
  wire zhuuhqdkyc6hr6he7stv5znjx3  ;
  wire b3s6npyd8da8fvpsu220ds      ;
  wire y27w4xcfx550bp04w6gr_ajr  ;
  wire duwii2jt5_0jetur15      ;
  wire ec34822n58n2jw42xoah940pd0m  ;
  wire djr037wb0rw8_ncab24vw      ;
  wire vscb6v0pa774vboyiiyxrfi3  ;
  wire kco4m_q5nhe0zxzcdxs88f      ;
  wire hxcw2yhpp4okeev3i1vp5rb  ;
  wire cg32iijl_44n51ppdlmca5p      ;
  wire ppml1670rwlohninqy2rv7xxl  ;
  wire s1561otgi027k9i6kmmlis      ;

  
  
  assign lkrl_gk1f715er9ueo    = !rc887zv55nqt[fnk0axwxfk4kr8z-1];
  wire   jgn947pmmcm9a77iuey     = (rc887zv55nqt == v_qy6klyvlpd9v    );
  wire   exn_cjm859bpb9zsghqr97  = (rc887zv55nqt == w7jie_pve8zo265khr8 ) & y0nv37yd84l;
  wire   dwmx63ax2_grri9q93qee = (rc887zv55nqt == w7jie_pve8zo265khr8);
  wire   k8wf2zd3daqs6q     = (rc887zv55nqt == elevjtxw8s86z    );
  wire   f1g98h1x6en1kemv1    = (rc887zv55nqt == r10y29zxz4oiu3wd    );
  wire   ee10pomiu8s7j7cn   = (rc887zv55nqt == zjl6he1ayeuql_m_f   );
  wire   t_o74lk4v_gxtrgop  = (rc887zv55nqt == m3aw6280mg3tu3ht0567);
  wire   is1to20_e01hc6      = (rc887zv55nqt == h_kmmziwjubh_5825      );
  wire   uk63nhcynwa_qtvrcek = (rc887zv55nqt == zj40kikmdbcd575xl7lmss);
  wire   yj737cz9t7gtb5     = (rc887zv55nqt == fvtdvg067g05k    );
  wire   umzor0sgk1r994nu3crx = (rc887zv55nqt == m9bvbk39_2zfrkcpc);
  wire   j3kfdsg0_toqfbv     = (rc887zv55nqt == sr0ftn45dhialfn    );
  wire   n43zel0f3h8f58krco8e = (rc887zv55nqt == d0ga83_71diabio74osj0);
  wire   dqkpvm9nx9kxryogn4     = (rc887zv55nqt == p0veyq__3ajbausg2h    );
  wire   rfes318a1jw5dtuzpbz2 = (rc887zv55nqt == x8jj4nrwgh_5270b_ftdv0);
  wire   d8f8tm6xf5hsinl8hf     = (rc887zv55nqt == saah2jpqh8i05    );
  wire   kgdwxspbwxi691glel5lgi6 = (rc887zv55nqt == gippr9ch9ni48cz3e47n);
  wire   oykqs2v1rwtrvt     = (rc887zv55nqt == zqlr7fq_zdgau_fa1r    );
  wire   lfm_3bqoo7ge6c9h9n_pse = (rc887zv55nqt == ar4t4ajioitfe1gtru35r);
  wire   hp16ita0zzndtl     = (rc887zv55nqt == eusn96ps48lsd4p    );


  wire [32-1:0] e4fbsnfdv8r;                       
  wire gdd8t8qjjaat37;
  wire oumac8m72aija2;
  wire kn_paijjp96y5sarclpoabo = &ggxoqcj7ytp1a4pjf7ee[1:0];
  wire f5ilaqqrs54pats = (e4fbsnfdv8r == bdqo1tgw2_bpi2e8alini) & gdd8t8qjjaat37 & !(oumac8m72aija2^kn_paijjp96y5sarclpoabo);  
  wire atqy1kayf2l1l2i = f5ilaqqrs54pats & gdd8t8qjjaat37 & x1huhi29x9mco & a2i6e7_7;   
  wire syokr6jqxk89zy8h = ((~f5ilaqqrs54pats) | (~gdd8t8qjjaat37)) & x1huhi29x9mco & a2i6e7_7;   

  
      
          
          
          
          
          
          
          
          
  wire x02_xmql777k8126zub0dp =    ( 1'b0  
                                 | fpo04urqz74
                                 | a2i6e7_7     
                                 | ldn2go4l40668ayimy
                                 );
  assign wfoen161d4r42bkqp34lj = lkrl_gk1f715er9ueo & x02_xmql777k8126zub0dp 
                               & (jrhs989pgz0z8or09
                                  | (syokr6jqxk89zy8h & wh1vvvsvv8tc2elyruo93)  
                               );
  assign u99tnldu986760c5      = 
                               a2i6e7_7 ? ((atqy1kayf2l1l2i | cw9xa748nw) ? elevjtxw8s86z : r10y29zxz4oiu3wd) :
                               v_qy6klyvlpd9v;
  assign wtgeux804w78dcd92swmjz7a5 = ee10pomiu8s7j7cn && xefc2nul9m648jueckdrui_l;
  assign lzbc5hwhr2m0yxt = m3aw6280mg3tu3ht0567;
  assign uwnli3a8y85_7gsqwb41d_ = t_o74lk4v_gxtrgop & woq47beoqkpu1um82nv58l1u_hyj4;
  assign zu_l0qkgxjl8mlhw = h_kmmziwjubh_5825;
  assign d2jegnujjeil20nht = is1to20_e01hc6;
  
  assign w9wl5ox_pnuvzp = w7jie_pve8zo265khr8;

      
          
  assign oz66a4n0vakndgbkbj6ds = jgn947pmmcm9a77iuey & b5b1bdkf9u8xkel6mtmr;
  assign g9natvym5lqakd      = 
                (
              
              
                  lgnnlckl1qq6psb ?  (w0vagcfu1v7wkym9f ? r10y29zxz4oiu3wd : chhrgp_9_w35oxb ? zjl6he1ayeuql_m_f : w7jie_pve8zo265khr8) :
                 
                  (y0nv37yd84l) ? w7jie_pve8zo265khr8 :  
                  v_qy6klyvlpd9v
                );
            
  wire  vij3v0mhh5pmf2niajrtl;
  wire  x2n1derqad2ie59_pd542m;
  wire  yzrjop7pz8lqhpmcv2wfbrz_u;
  wire [64-1:0] clur09du62kjid;
  wire xy7mzrc3a5aq_a; 
  wire oq9g104cbco28bc35hbhw = (clur09du62kjid[2:0] == 3'b000) & chhrgp_9_w35oxb; 
  wire de5wl59a329ve2vf4kqilfp8cr = oq9g104cbco28bc35hbhw & xy7mzrc3a5aq_a; 
      
  assign odvuoxdd_64egspdavi73jis74 = dwmx63ax2_grri9q93qee & (zjmbnwsbyle24ayly67 | vij3v0mhh5pmf2niajrtl | x2n1derqad2ie59_pd542m | yzrjop7pz8lqhpmcv2wfbrz_u | de5wl59a329ve2vf4kqilfp8cr);
              
  assign qyw9w17wm01o0ibqri8      = (vij3v0mhh5pmf2niajrtl | x2n1derqad2ie59_pd542m | yzrjop7pz8lqhpmcv2wfbrz_u | de5wl59a329ve2vf4kqilfp8cr) ? r10y29zxz4oiu3wd : elevjtxw8s86z;
  
      
          
  assign z5xqhvuiqp_g510lj8 = k8wf2zd3daqs6q & b5b1bdkf9u8xkel6mtmr;
  assign evn7vmlv0q87c      = 
                (
              
              
                  (lgnnlckl1qq6psb & (d74326txgko0 || cfe949_7aiw) ) ?  (w0vagcfu1v7wkym9f ? r10y29zxz4oiu3wd : zj40kikmdbcd575xl7lmss) : 
                
                  r10y29zxz4oiu3wd 
                );

  
  assign zhuuhqdkyc6hr6he7stv5znjx3 = uk63nhcynwa_qtvrcek & (zjmbnwsbyle24ayly67 | vij3v0mhh5pmf2niajrtl | x2n1derqad2ie59_pd542m | yzrjop7pz8lqhpmcv2wfbrz_u | de5wl59a329ve2vf4kqilfp8cr);
              
  assign etqkl_z3d5k_z3n1fr      = (vij3v0mhh5pmf2niajrtl | x2n1derqad2ie59_pd542m | yzrjop7pz8lqhpmcv2wfbrz_u | de5wl59a329ve2vf4kqilfp8cr) ? r10y29zxz4oiu3wd : fvtdvg067g05k;

  
          
  assign b3s6npyd8da8fvpsu220ds = yj737cz9t7gtb5 & b5b1bdkf9u8xkel6mtmr;
  assign yqwi1z4q7s0wriam8      =                                
                (
              
              
                  (w0vagcfu1v7wkym9f ? r10y29zxz4oiu3wd : m9bvbk39_2zfrkcpc)
                );

  
  assign y27w4xcfx550bp04w6gr_ajr = umzor0sgk1r994nu3crx & (zjmbnwsbyle24ayly67 | vij3v0mhh5pmf2niajrtl | x2n1derqad2ie59_pd542m | yzrjop7pz8lqhpmcv2wfbrz_u | de5wl59a329ve2vf4kqilfp8cr);
              
  assign g897ues2orwmfihybd      = (vij3v0mhh5pmf2niajrtl | x2n1derqad2ie59_pd542m | yzrjop7pz8lqhpmcv2wfbrz_u | de5wl59a329ve2vf4kqilfp8cr) ? r10y29zxz4oiu3wd : sr0ftn45dhialfn;

  
          
  assign duwii2jt5_0jetur15 = j3kfdsg0_toqfbv & b5b1bdkf9u8xkel6mtmr;
  assign skmlitjb4kdramm      =                                
                (
                  (lgnnlckl1qq6psb & cfe949_7aiw) ?  (w0vagcfu1v7wkym9f ? r10y29zxz4oiu3wd : d0ga83_71diabio74osj0) : 
                  r10y29zxz4oiu3wd 
                );

  assign ec34822n58n2jw42xoah940pd0m = n43zel0f3h8f58krco8e & (zjmbnwsbyle24ayly67 | vij3v0mhh5pmf2niajrtl | x2n1derqad2ie59_pd542m | yzrjop7pz8lqhpmcv2wfbrz_u | de5wl59a329ve2vf4kqilfp8cr);
  assign uv3o5o9wdyyhfp16ijtnst      = (vij3v0mhh5pmf2niajrtl | x2n1derqad2ie59_pd542m | yzrjop7pz8lqhpmcv2wfbrz_u | de5wl59a329ve2vf4kqilfp8cr) ? r10y29zxz4oiu3wd : p0veyq__3ajbausg2h;
  assign djr037wb0rw8_ncab24vw = dqkpvm9nx9kxryogn4 & b5b1bdkf9u8xkel6mtmr;
  assign c9v_t190cck33l9      = w0vagcfu1v7wkym9f ? r10y29zxz4oiu3wd : x8jj4nrwgh_5270b_ftdv0;

  assign vscb6v0pa774vboyiiyxrfi3 = rfes318a1jw5dtuzpbz2 & (zjmbnwsbyle24ayly67 | vij3v0mhh5pmf2niajrtl | x2n1derqad2ie59_pd542m | yzrjop7pz8lqhpmcv2wfbrz_u | de5wl59a329ve2vf4kqilfp8cr);
  assign anh_5y93ex8mfy8zqs4h      = (vij3v0mhh5pmf2niajrtl | x2n1derqad2ie59_pd542m | yzrjop7pz8lqhpmcv2wfbrz_u | de5wl59a329ve2vf4kqilfp8cr) ? r10y29zxz4oiu3wd : saah2jpqh8i05;
  assign kco4m_q5nhe0zxzcdxs88f = d8f8tm6xf5hsinl8hf & b5b1bdkf9u8xkel6mtmr;
  assign i41gux5i8cqjqp      = w0vagcfu1v7wkym9f ? r10y29zxz4oiu3wd : gippr9ch9ni48cz3e47n;

  assign hxcw2yhpp4okeev3i1vp5rb = kgdwxspbwxi691glel5lgi6 & (zjmbnwsbyle24ayly67 | vij3v0mhh5pmf2niajrtl | x2n1derqad2ie59_pd542m | yzrjop7pz8lqhpmcv2wfbrz_u | de5wl59a329ve2vf4kqilfp8cr);
  assign v_nz7nezxqthl8mkc      = (vij3v0mhh5pmf2niajrtl | x2n1derqad2ie59_pd542m | yzrjop7pz8lqhpmcv2wfbrz_u | de5wl59a329ve2vf4kqilfp8cr) ? r10y29zxz4oiu3wd : zqlr7fq_zdgau_fa1r;
  assign cg32iijl_44n51ppdlmca5p = oykqs2v1rwtrvt & b5b1bdkf9u8xkel6mtmr;
  assign dxqq9l9bv3v20jsdv      = w0vagcfu1v7wkym9f ? r10y29zxz4oiu3wd : ar4t4ajioitfe1gtru35r;

  assign ppml1670rwlohninqy2rv7xxl = lfm_3bqoo7ge6c9h9n_pse & (zjmbnwsbyle24ayly67 | vij3v0mhh5pmf2niajrtl | x2n1derqad2ie59_pd542m | yzrjop7pz8lqhpmcv2wfbrz_u | de5wl59a329ve2vf4kqilfp8cr);
  assign h5chs70629xcwrlur      = (vij3v0mhh5pmf2niajrtl | x2n1derqad2ie59_pd542m | yzrjop7pz8lqhpmcv2wfbrz_u | de5wl59a329ve2vf4kqilfp8cr) ? r10y29zxz4oiu3wd : eusn96ps48lsd4p;
  assign s1561otgi027k9i6kmmlis = hp16ita0zzndtl & b5b1bdkf9u8xkel6mtmr;
  assign auqrmggnbde5eb      = r10y29zxz4oiu3wd;
  
    
          
              
              
  wire y691hsyucyt;
  wire weqk4hvu3gan052;
  wire fznp6w7g_ncdmns_q;
  wire dsk0idxv2xoskrfgzv91rnwzo;
  assign weqk4hvu3gan052 = j98f_s869qm5bv_dhgbcim3 || wfoen161d4r42bkqp34lj;
  assign fznp6w7g_ncdmns_q = syokr6jqxk89zy8h && lkrl_gk1f715er9ueo;
  assign dsk0idxv2xoskrfgzv91rnwzo = y691hsyucyt ? !xhpc6eofokpbnya1h3s117_2 : 1'b1;
  
  ux607_gnrl_dfflr #(1) kqk1ikhuss_i1a (weqk4hvu3gan052, fznp6w7g_ncdmns_q, y691hsyucyt, gf33atgy, ru_wi);
  
  assign j98f_s869qm5bv_dhgbcim3 = f1g98h1x6en1kemv1 & dsk0idxv2xoskrfgzv91rnwzo & rxjuugktc38un;
  assign gyiivu76k6m_fi      = i3mg661fq9njsp5b;





    
  assign gsoquod_6th_uva = 1'b0 
            | wfoen161d4r42bkqp34lj 
            | oz66a4n0vakndgbkbj6ds  
            | wtgeux804w78dcd92swmjz7a5  
            | uwnli3a8y85_7gsqwb41d_  
            | d2jegnujjeil20nht  
            | odvuoxdd_64egspdavi73jis74 
            | z5xqhvuiqp_g510lj8   
            | j98f_s869qm5bv_dhgbcim3 
            | zhuuhqdkyc6hr6he7stv5znjx3 
            | b3s6npyd8da8fvpsu220ds   
            | y27w4xcfx550bp04w6gr_ajr 
            | duwii2jt5_0jetur15 
            | ec34822n58n2jw42xoah940pd0m 
            | vscb6v0pa774vboyiiyxrfi3 
            | hxcw2yhpp4okeev3i1vp5rb 
            | ppml1670rwlohninqy2rv7xxl 
            | djr037wb0rw8_ncab24vw 
            | kco4m_q5nhe0zxzcdxs88f 
            | cg32iijl_44n51ppdlmca5p 
            | s1561otgi027k9i6kmmlis 
          ;

  
  assign brgdc0amsvlnwf_2j = 
              ({fnk0axwxfk4kr8z{1'b0}})
            | ({fnk0axwxfk4kr8z{wfoen161d4r42bkqp34lj   }} & u99tnldu986760c5   )
            | ({fnk0axwxfk4kr8z{oz66a4n0vakndgbkbj6ds    }} & g9natvym5lqakd    )
            | ({fnk0axwxfk4kr8z{odvuoxdd_64egspdavi73jis74}} & qyw9w17wm01o0ibqri8)
            | ({fnk0axwxfk4kr8z{z5xqhvuiqp_g510lj8    }} & evn7vmlv0q87c    )
            | ({fnk0axwxfk4kr8z{j98f_s869qm5bv_dhgbcim3   }} & gyiivu76k6m_fi   )
            | ({fnk0axwxfk4kr8z{wtgeux804w78dcd92swmjz7a5  }} & lzbc5hwhr2m0yxt  )
            | ({fnk0axwxfk4kr8z{uwnli3a8y85_7gsqwb41d_ }} & zu_l0qkgxjl8mlhw )
            | ({fnk0axwxfk4kr8z{d2jegnujjeil20nht     }} & w9wl5ox_pnuvzp     )
            | ({fnk0axwxfk4kr8z{zhuuhqdkyc6hr6he7stv5znjx3}} & etqkl_z3d5k_z3n1fr)
            | ({fnk0axwxfk4kr8z{b3s6npyd8da8fvpsu220ds    }} & yqwi1z4q7s0wriam8    )
            | ({fnk0axwxfk4kr8z{y27w4xcfx550bp04w6gr_ajr}} & g897ues2orwmfihybd)
            | ({fnk0axwxfk4kr8z{duwii2jt5_0jetur15    }} & skmlitjb4kdramm    )
            | ({fnk0axwxfk4kr8z{ec34822n58n2jw42xoah940pd0m}} & uv3o5o9wdyyhfp16ijtnst)
            | ({fnk0axwxfk4kr8z{vscb6v0pa774vboyiiyxrfi3}} & anh_5y93ex8mfy8zqs4h)
            | ({fnk0axwxfk4kr8z{hxcw2yhpp4okeev3i1vp5rb}} & v_nz7nezxqthl8mkc)
            | ({fnk0axwxfk4kr8z{ppml1670rwlohninqy2rv7xxl}} & h5chs70629xcwrlur)
            | ({fnk0axwxfk4kr8z{djr037wb0rw8_ncab24vw    }} & c9v_t190cck33l9    )
            | ({fnk0axwxfk4kr8z{kco4m_q5nhe0zxzcdxs88f    }} & i41gux5i8cqjqp    )
            | ({fnk0axwxfk4kr8z{cg32iijl_44n51ppdlmca5p    }} & dxqq9l9bv3v20jsdv    )
            | ({fnk0axwxfk4kr8z{s1561otgi027k9i6kmmlis    }} & auqrmggnbde5eb    )
              ;


  ux607_gnrl_dfflr #(fnk0axwxfk4kr8z) qo3f12wu71_4hg0af7 (gsoquod_6th_uva, brgdc0amsvlnwf_2j, rc887zv55nqt, gf33atgy, ru_wi);

  wire jgsfpfezq31q01b2w0in = gsoquod_6th_uva & (brgdc0amsvlnwf_2j == v_qy6klyvlpd9v);
  wire c2q6lda5ak6w6cr45iz_q4 = gsoquod_6th_uva & (brgdc0amsvlnwf_2j == r10y29zxz4oiu3wd);

  wire ncd2vzr5v7ahxaqgb = f1g98h1x6en1kemv1 & dsk0idxv2xoskrfgzv91rnwzo;
  wire ly9og56m3h2etesc4bxfxm = j98f_s869qm5bv_dhgbcim3;



  assign j2_lz0mpsxf4xotgqf1ngx = ((~lkrl_gk1f715er9ueo) | badsf4ksbp3k6p_p5hnj2i);

  
  wire ixsuwxurdtzqx2q1h = gsoquod_6th_uva;
  wire diopbpeh9cwbka2_ey = (brgdc0amsvlnwf_2j != i3mg661fq9njsp5b);
  wire ta_47w4l6age6uy;
  wire x1hlyprlmbf5iq1uax;

  ux607_gnrl_dfflr #(1) eqs_nld6yjpb8x7d9lr (gsoquod_6th_uva, diopbpeh9cwbka2_ey, ta_47w4l6age6uy, gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1) txqv6vrcabwp618nb3p_10b (gsoquod_6th_uva, diopbpeh9cwbka2_ey, x1hlyprlmbf5iq1uax, gf33atgy, ru_wi);

  assign hcugdkhp9szims1nk8rhakn = ta_47w4l6age6uy;
  assign dw2ygdedledlm7ps830qgbwonu = x1hlyprlmbf5iq1uax;
  
  
  
  wire q4zlija4136s_s9d;
  wire [64-1:0] aafyam17vrqz;
  wire [64-1:0] h3p0wpn_ah;
  wire zbyyzobw24m3mrvv0l;
  wire laa1t5iskus82m9g;
  wire omyw5_07_btxhfwq;

  wire k_ieqlp1d1jh734g;
  wire [64-1:0] famxn7sdgfd7riib4i6;
  
  wire dfdmudd4z4p = jgn947pmmcm9a77iuey & y0nv37yd84l;
  wire ke43_l21ebj7w = k8wf2zd3daqs6q & y0nv37yd84l;

  wire swiq3rmoa0huticg4f2z = a2i6e7_7 & cw9xa748nw & wfoen161d4r42bkqp34lj;
  wire vk_o92k7vyx0f84e4tjfbl = syokr6jqxk89zy8h & wfoen161d4r42bkqp34lj;
  wire l2kas5gsiruf5xw6z_b = k8wf2zd3daqs6q & ai2cjirv & qndyhstqm8pvl;
  wire aus6tfj37uprs0ut91l = k8wf2zd3daqs6q & ai2cjirv & qj_5hjk5ts;


  wire uwe7v51c63wk_yn2thuaw = lgf34_8i5f2254 & wfoen161d4r42bkqp34lj;
  wire tvnalus6r57_3jx4uxpz   = u9y07o_n2vgf1zk   & wfoen161d4r42bkqp34lj;
  wire prkdsv0vdtofmvtx16okku = ldn2go4l40668ayimy & wfoen161d4r42bkqp34lj;
  wire m6ssh2_3bt1uudxdqps7jc54qj = ldn2go4l40668ayimy & lkrl_gk1f715er9ueo;
  wire zw_spwk8rmb88ctbzxs_bwwa3c   = u9y07o_n2vgf1zk   & lkrl_gk1f715er9ueo; 
  wire xhaudj8i3rv = ( jgn947pmmcm9a77iuey 
                        | k8wf2zd3daqs6q
                        | yj737cz9t7gtb5
                        | j3kfdsg0_toqfbv
                        | dqkpvm9nx9kxryogn4
                        | d8f8tm6xf5hsinl8hf
                        | oykqs2v1rwtrvt
                        | hp16ita0zzndtl
                        );
  wire eqvc72yrtjp8tx0zny = xhaudj8i3rv & ijk5d1s_9m5n;
  wire tiyz26xe8652bejo2976li = xhaudj8i3rv & lgnnlckl1qq6psb;



                 
  
  wire [8-1:0] d45di3rfd8m8oxlob = 
                                  ({8{(clur09du62kjid[2:0] == 3'b000)}} & gxo5tf4bea2gsq4yyn[7:0])      
                                | ({8{(clur09du62kjid[2:0] == 3'b001)}} & gxo5tf4bea2gsq4yyn[15:8])      
                                | ({8{(clur09du62kjid[2:0] == 3'b010)}} & gxo5tf4bea2gsq4yyn[23:16])      
                                | ({8{(clur09du62kjid[2:0] == 3'b011)}} & gxo5tf4bea2gsq4yyn[31:24])      
                                | ({8{(clur09du62kjid[2:0] == 3'b100)}} & gxo5tf4bea2gsq4yyn[39:32])      
                                | ({8{(clur09du62kjid[2:0] == 3'b101)}} & gxo5tf4bea2gsq4yyn[47:40])      
                                | ({8{(clur09du62kjid[2:0] == 3'b110)}} & gxo5tf4bea2gsq4yyn[55:48])      
                                | ({8{(clur09du62kjid[2:0] == 3'b111)}} & gxo5tf4bea2gsq4yyn[63:56])      
                                ;
  wire [64-1:0] pbm3dgk9csubydfkemlll = {8{d45di3rfd8m8oxlob}};
  
  
  
  
  
  
  
  
  

  wire [64-1:0] p4bzwo27__g97d = 
            ({64{jgn947pmmcm9a77iuey}} & 64'h0000_00FF)
          | ({64{k8wf2zd3daqs6q}} & 64'h0000_FF00)
          | ({64{yj737cz9t7gtb5}} & 64'h00FF_0000)
          | ({64{j3kfdsg0_toqfbv}} & 64'hFF00_0000)
          | ({64{dqkpvm9nx9kxryogn4}} & 64'h0000_00FF_0000_0000)
          | ({64{d8f8tm6xf5hsinl8hf}} & 64'h0000_FF00_0000_0000)
          | ({64{oykqs2v1rwtrvt}} & 64'h00FF_0000_0000_0000)
          | ({64{hp16ita0zzndtl}} & 64'hFF00_0000_0000_0000)
          ;


  wire [64-1:0] kk4oak80apbqjpua8czd8pxn = ((h3p0wpn_ah & (~p4bzwo27__g97d)) | (pbm3dgk9csubydfkemlll[64-1:0] & p4bzwo27__g97d));


  wire jjzjfxy52faix = (glc7xaf_upxku  &   deonbdggc2hhsqq88);
  wire plecoe0fogguy  = (glc7xaf_upxku  & (~deonbdggc2hhsqq88));
  wire idkjxjm61isg = (d74326txgko0  &   deonbdggc2hhsqq88);
  wire zif3xp2n85v1  = (d74326txgko0  & (~deonbdggc2hhsqq88)) & (~encgymm9xrq0);
  wire gjuvgwnbequ57 = (d74326txgko0  & (~deonbdggc2hhsqq88)) & ( encgymm9xrq0);
  wire zyrfrwzdmuy  =  cfe949_7aiw;

  wire [64-1:0] uii11g83mbu8xigaa55 = 64'b0
          | ({64{jjzjfxy52faix}} & {{64-16{          1'b0}}, h3p0wpn_ah[15:0]})
          | ({64{plecoe0fogguy }} & {{64-16{h3p0wpn_ah[15]}}, h3p0wpn_ah[15:0]}) 
          | ({64{idkjxjm61isg}} & {{64-32{          1'b0}}, h3p0wpn_ah[31:0]})
          | ({64{zif3xp2n85v1 }} & {{64-32{h3p0wpn_ah[31]}}, h3p0wpn_ah[31:0]})
          | ({64{gjuvgwnbequ57}} & {{64-32{          1'b1}}, h3p0wpn_ah[31:0]})
          | ({64{zyrfrwzdmuy }} & {                                 h3p0wpn_ah      })
          ;


  assign q4zlija4136s_s9d = (
                   1'b0
                   | (b5b1bdkf9u8xkel6mtmr & dfdmudd4z4p) 
                   
                   | vk_o92k7vyx0f84e4tjfbl                    
                   | (b5b1bdkf9u8xkel6mtmr & l2kas5gsiruf5xw6z_b) 
                   | (b5b1bdkf9u8xkel6mtmr & aus6tfj37uprs0ut91l) 
                   | tvnalus6r57_3jx4uxpz
                   | (b5b1bdkf9u8xkel6mtmr & eqvc72yrtjp8tx0zny) 
                   );

  assign aafyam17vrqz = 
              {64{1'b0}}
            | ({64{dfdmudd4z4p        }} & fn5e7uint162p6axap1i1t9[64-1:0])
            
            | ({64{vk_o92k7vyx0f84e4tjfbl}} & 64'h1)            
            | ({64{l2kas5gsiruf5xw6z_b   }} & fn5e7uint162p6axap1i1t9[64-1:0])
            | ({64{aus6tfj37uprs0ut91l   }} & 64'h0)            
            | ({64{zw_spwk8rmb88ctbzxs_bwwa3c}} & a4a48egkdkec8d9b_9[64-1:0])
            | ({64{eqvc72yrtjp8tx0zny}} & kk4oak80apbqjpua8czd8pxn)
            ;
 

  assign zbyyzobw24m3mrvv0l = 1'b0 
                   | (b5b1bdkf9u8xkel6mtmr & dfdmudd4z4p) 
                   | (b5b1bdkf9u8xkel6mtmr & ke43_l21ebj7w) 
                   | vk_o92k7vyx0f84e4tjfbl                             
                   | (b5b1bdkf9u8xkel6mtmr & l2kas5gsiruf5xw6z_b)
                   | (b5b1bdkf9u8xkel6mtmr & aus6tfj37uprs0ut91l)
                   | (b5b1bdkf9u8xkel6mtmr & tiyz26xe8652bejo2976li) 
         ;

  assign laa1t5iskus82m9g = 1'b0 
            | (dfdmudd4z4p           & w0vagcfu1v7wkym9f)
            | (ke43_l21ebj7w           & (w0vagcfu1v7wkym9f | omyw5_07_btxhfwq))
            | (vk_o92k7vyx0f84e4tjfbl   & 1'b0)           
            | (l2kas5gsiruf5xw6z_b      & w0vagcfu1v7wkym9f)
            | (aus6tfj37uprs0ut91l      & w0vagcfu1v7wkym9f)
            | (tiyz26xe8652bejo2976li   & w0vagcfu1v7wkym9f) 
         ;


  wire pdt4373c_z67vejmh = swiq3rmoa0huticg4f2z;                        
  wire gh0ee01r3ez3xi31 = (wh1vvvsvv8tc2elyruo93 & ~pdt4373c_z67vejmh)      
                       | (l2kas5gsiruf5xw6z_b & w0vagcfu1v7wkym9f)
					   ;
  wire o6b354_5y5bidwlagt = pdt4373c_z67vejmh |  gh0ee01r3ez3xi31;
  wire h_m3swnk1wvddoekta = pdt4373c_z67vejmh | ~gh0ee01r3ez3xi31;
  wire i5zwrqgdlu506t8 = pdt4373c_z67vejmh;
  
  
  assign e__67e1k5hdb4ctnr = q4zlija4136s_s9d;
  assign jay_5c6ndpwhj0vqzv = aafyam17vrqz;
  assign h3p0wpn_ah    = kn6tx97_rw9w0v;

  
  ux607_gnrl_dfflr #(1) sobaz4rsptel5wvuxaj4hpnheg (zbyyzobw24m3mrvv0l, laa1t5iskus82m9g, omyw5_07_btxhfwq, gf33atgy, ru_wi);


  wire r9y8upslfevdvznk53cw;      
  wire hd4oskx3f3ljlt7dh1b515f =   c2q6lda5ak6w6cr45iz_q4 
                             ;
  wire xr82kspf8yl7mns9yxa4 = 
                               1'b0
                             | (dwmx63ax2_grri9q93qee  & c2q6lda5ak6w6cr45iz_q4 & vij3v0mhh5pmf2niajrtl)
                             | (uk63nhcynwa_qtvrcek  & c2q6lda5ak6w6cr45iz_q4 & vij3v0mhh5pmf2niajrtl)
                             | (umzor0sgk1r994nu3crx  & c2q6lda5ak6w6cr45iz_q4 & vij3v0mhh5pmf2niajrtl)
                             | (n43zel0f3h8f58krco8e  & c2q6lda5ak6w6cr45iz_q4 & vij3v0mhh5pmf2niajrtl)
                             | (rfes318a1jw5dtuzpbz2  & c2q6lda5ak6w6cr45iz_q4 & vij3v0mhh5pmf2niajrtl)
                             | (kgdwxspbwxi691glel5lgi6  & c2q6lda5ak6w6cr45iz_q4 & vij3v0mhh5pmf2niajrtl)
                             | (lfm_3bqoo7ge6c9h9n_pse  & c2q6lda5ak6w6cr45iz_q4 & vij3v0mhh5pmf2niajrtl)
                             ;

  ux607_gnrl_dfflr #(1) i22p6rl565jmmhscw2x93426gxz1 (hd4oskx3f3ljlt7dh1b515f, xr82kspf8yl7mns9yxa4, r9y8upslfevdvznk53cw, gf33atgy, ru_wi);

  wire rdbfve_zy3rsium8rq7uj;      
  wire ocwtw05k197_ekfhymxl3_9c =   c2q6lda5ak6w6cr45iz_q4 
                             ;
  wire y578z9gcc5q8hmox0rvm7 = 
                               1'b0
                             | (dwmx63ax2_grri9q93qee  & c2q6lda5ak6w6cr45iz_q4 & x2n1derqad2ie59_pd542m)
                             | (uk63nhcynwa_qtvrcek  & c2q6lda5ak6w6cr45iz_q4 & x2n1derqad2ie59_pd542m)
                             | (umzor0sgk1r994nu3crx  & c2q6lda5ak6w6cr45iz_q4 & x2n1derqad2ie59_pd542m)
                             ;

  ux607_gnrl_dfflr #(1) d6hoed6k6qq49pe6isxuk6_f8sqmdq (ocwtw05k197_ekfhymxl3_9c, y578z9gcc5q8hmox0rvm7, rdbfve_zy3rsium8rq7uj, gf33atgy, ru_wi);

  wire cp18rjpfmjtvgxyp9a;      
  wire ca0h4znd_tvixumg9zke =   c2q6lda5ak6w6cr45iz_q4 
                             ;
  wire cw3bqsbjf_ydogfz82w = 
                               1'b0
                             | (dwmx63ax2_grri9q93qee  & c2q6lda5ak6w6cr45iz_q4 & yzrjop7pz8lqhpmcv2wfbrz_u)
                             | (uk63nhcynwa_qtvrcek  & c2q6lda5ak6w6cr45iz_q4 & yzrjop7pz8lqhpmcv2wfbrz_u)
                             | (umzor0sgk1r994nu3crx  & c2q6lda5ak6w6cr45iz_q4 & yzrjop7pz8lqhpmcv2wfbrz_u)
                             ;

  ux607_gnrl_dfflr #(1) prakd4c7am1m1lxzl16118idv154m (ca0h4znd_tvixumg9zke, cw3bqsbjf_ydogfz82w, cp18rjpfmjtvgxyp9a, gf33atgy, ru_wi);

  ux607_gnrl_dfflr #(1) zx2z7v6c_8vbc6h7kak (o6b354_5y5bidwlagt, h_m3swnk1wvddoekta, gdd8t8qjjaat37, gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1) lupsep2x2zk_aqp8_ (i5zwrqgdlu506t8, kn_paijjp96y5sarclpoabo, oumac8m72aija2, gf33atgy, ru_wi);
  
  
  
  wire g_4x7gokhlckvss_y4g4fk14u = (prkdsv0vdtofmvtx16okku)
                              | ( (  jgn947pmmcm9a77iuey 
                                   | k8wf2zd3daqs6q
                                   | yj737cz9t7gtb5
                                   | j3kfdsg0_toqfbv
                                   | dqkpvm9nx9kxryogn4
                                   | d8f8tm6xf5hsinl8hf
                                   | oykqs2v1rwtrvt
                                   | hp16ita0zzndtl
                                   ) 
                                   & lgnnlckl1qq6psb & b5b1bdkf9u8xkel6mtmr & (~w0vagcfu1v7wkym9f)
                                 );
  
  wire r8u3n7sxmz6ig = fpo04urqz74 & wfoen161d4r42bkqp34lj;
  wire tg6dl6cdzg8cdxg93 = a2i6e7_7 & wfoen161d4r42bkqp34lj;
  wire goefkr663a4o90wdkcs60017huc9e = de5wl59a329ve2vf4kqilfp8cr & (
                                                                 dwmx63ax2_grri9q93qee
                                                               | uk63nhcynwa_qtvrcek
                                                               | umzor0sgk1r994nu3crx
                                                               | n43zel0f3h8f58krco8e
                                                               | rfes318a1jw5dtuzpbz2
                                                               | kgdwxspbwxi691glel5lgi6
                                                               | lfm_3bqoo7ge6c9h9n_pse
                                                              );
  assign k_ieqlp1d1jh734g = 1'b0 
             | r8u3n7sxmz6ig     
             | tg6dl6cdzg8cdxg93        
           | g_4x7gokhlckvss_y4g4fk14u
         
           | goefkr663a4o90wdkcs60017huc9e
         ;
  assign famxn7sdgfd7riib4i6 = (
                           prkdsv0vdtofmvtx16okku   
                          | r8u3n7sxmz6ig
                          | tg6dl6cdzg8cdxg93    
                          ) ? bdqo1tgw2_bpi2e8alini : 
                           ttgsydregi0kgoj_z; 
  
  
  assign nc_3q2q5fz4e2   = k_ieqlp1d1jh734g;
  assign a5y809wbv8w1d0   = famxn7sdgfd7riib4i6;
  assign clur09du62kjid = l0vxn4vg6wd;
  assign e4fbsnfdv8r = clur09du62kjid[32-1:0];    


  
  assign xl9r7gr7wciuv2d00b  = 1'b0
                           | (exn_cjm859bpb9zsghqr97 & qdiehi55s8izv5y)
                           | (lgnnlckl1qq6psb & (jgn947pmmcm9a77iuey  
                                              | k8wf2zd3daqs6q 
                                              | yj737cz9t7gtb5 
                                              | j3kfdsg0_toqfbv 
                                              | dqkpvm9nx9kxryogn4 
                                              | d8f8tm6xf5hsinl8hf 
                                              | oykqs2v1rwtrvt 
                                              | hp16ita0zzndtl 
                                              ) 
                             )
                           | (ee10pomiu8s7j7cn)            
                           | (goefkr663a4o90wdkcs60017huc9e)
                           
                           ;

  assign tp6hfcjxcyp899mpksjl =  
                            exn_cjm859bpb9zsghqr97 ? h3p0wpn_ah :
                           ee10pomiu8s7j7cn            ? {wqbvx_uqjrfzj8cjke712tpq[64-1:12],12'h0} : 
                           goefkr663a4o90wdkcs60017huc9e ? {wqbvx_uqjrfzj8cjke712tpq[64-1:12],12'h0} :
                           m6ssh2_3bt1uudxdqps7jc54qj ? wqbvx_uqjrfzj8cjke712tpq : clur09du62kjid 
                     ;

  assign f4ds8dbk9kk_ic_ =  
                            exn_cjm859bpb9zsghqr97 ? i200dby :
                           ee10pomiu8s7j7cn            ? 64'h1000 : 
                           goefkr663a4o90wdkcs60017huc9e ? 64'h1000 :
                            64'd1 
                     ;

  assign oso3fj0gx6pnvjni =  euomkrkdp_x2p16;
  assign htcsb0affil7c6q  =  hksju1a__h21 ;
  assign vrqdq7uwxf99gj_7   =  yod75j20uh  ;
  assign jqgtsdtxss_uios07  =  v_zd2akdl84 ;
  assign hn2h_gkqinydwsdg_i3  =  u1npc4m1kjg ;
  assign re8hncw6m47hrh6  =  ybfhwehnrx61b8 ;
  assign tshku7fgpiu2j7ugwjj9 =  ed7pawk0e32us153;
  assign arc8ztjel_qlz3xfw0ya =  gg2d7pi35s036m89;
  assign dukom1hk2mc9i6m4   =  cfe949_7aiw || 
                              ~y0nv37yd84l
                            ;





  assign ed4kcy8s9nrisftgx_q =   (lkrl_gk1f715er9ueo & zjmbnwsbyle24ayly67);
  
  


  assign jugi02ecegnos3 = 
        ncd2vzr5v7ahxaqgb 
      ;

  
  assign h8wu7unf_ixmxfeh = {64{1'b0 }}
                    | ({64{ijk5d1s_9m5n }} & uii11g83mbu8xigaa55)
                    | ({64{qxeco0b4xvxw1v }} & 64'b0 )
                    | ({64{y0nv37yd84l      }} & h3p0wpn_ah    ) 
                    | ({64{ai2cjirv     }} & h3p0wpn_ah    ) 
       ;
  

  
  
  
  
  
  
  
  
  
  
  
  

  wire yoop58jcvoblafgy3pvb2bxf;
  wire x79p6ptdcs3v1b_ri0qmwfye;
  wire sc7qvopbyz8bul4k_h_57;
  wire sl4tlevefghkwtcz94e4u87ss8;
  wire pc2lfcg8w9met4at0tga_8g;
  wire ycrhycedz35gkapfocflviq = 1'b0;
  wire ih29gu5ovqcto6pzh = 1'b0;

  assign {x79p6ptdcs3v1b_ri0qmwfye, sc7qvopbyz8bul4k_h_57, pc2lfcg8w9met4at0tga_8g, sl4tlevefghkwtcz94e4u87ss8} = (4'b0 
                      | ({4{lgnnlckl1qq6psb  }} & {omyw5_07_btxhfwq, r9y8upslfevdvznk53cw, rdbfve_zy3rsium8rq7uj, cp18rjpfmjtvgxyp9a})
                      | ({4{y0nv37yd84l         }} & {omyw5_07_btxhfwq, 3'b0})
                      | ({4{ai2cjirv        }} & {omyw5_07_btxhfwq, 3'b0}) 
                      )
                ;

   assign kdpgigzs75vcc1d  = adng7z_1b3srxoxai1rm;
   assign coohnlu_ri   = x79p6ptdcs3v1b_ri0qmwfye | sc7qvopbyz8bul4k_h_57 | ycrhycedz35gkapfocflviq | ih29gu5ovqcto6pzh
                        |ks33bi5hojtg0te9bl7   | eht8nc5zc5sdbpe9nqr67jeju
                         ;
   assign igo49dpz9ealh4h13a   = (sc7qvopbyz8bul4k_h_57 & ~yoop58jcvoblafgy3pvb2bxf)
                               | eht8nc5zc5sdbpe9nqr67jeju
                               ;
   assign x6uy7s6mcepqq2j527jtxk   = coohnlu_ri;

   assign dwet7q3ucodidho7qxlw = (lgnnlckl1qq6psb 
                                | y0nv37yd84l
                                | ai2cjirv
							   ) ? clur09du62kjid[64-1:0] : 64'b0;
   assign k5h5ux92dlz_nn0    = qndyhstqm8pvl;
   assign e6uinbhqc8o7iylg7d = qj_5hjk5ts 
                           | y0nv37yd84l
                           ;
   assign p_p6yt19xmgqbfsn0y    = trgbsbj;



  

  assign epoc75xqnuvcqziu_9i55h = 
        1'b1;


  

  assign qsw59ks9jxcsmmh   = o21b8ypt1xiu5ml63d | (~lkrl_gk1f715er9ueo);       
  assign aht5xalx865dt9ymg6t4 = lkrl_gk1f715er9ueo ?
                            (
                             (atqy1kayf2l1l2i | cw9xa748nw | ~a2i6e7_7) & 
                             badsf4ksbp3k6p_p5hnj2i ) :       
                            ((  dwmx63ax2_grri9q93qee
                             | uk63nhcynwa_qtvrcek
                             | umzor0sgk1r994nu3crx
                             | n43zel0f3h8f58krco8e
                             | rfes318a1jw5dtuzpbz2
                             | kgdwxspbwxi691glel5lgi6
                             | lfm_3bqoo7ge6c9h9n_pse
                             | exn_cjm859bpb9zsghqr97       
                            ) & (~(vij3v0mhh5pmf2niajrtl | x2n1derqad2ie59_pd542m | yzrjop7pz8lqhpmcv2wfbrz_u | de5wl59a329ve2vf4kqilfp8cr)))
                            ;
  assign icfwo5l56zab795f[11:0] = (~lkrl_gk1f715er9ueo) ? clur09du62kjid[11:0] :
                                                       bdqo1tgw2_bpi2e8alini[11:0] ;
  assign icfwo5l56zab795f[32-1:12] = (lkrl_gk1f715er9ueo) ?                       bdqo1tgw2_bpi2e8alini[32-1:12]                  :
                                                  (f8ouikbgg2hqwm8g | ~chhrgp_9_w35oxb) ?      clur09du62kjid[32-1:12]                  :
                                                  
                                                  (dvqdxyi_ja1x2 == clur09du62kjid[12]) ?      clur09du62kjid[32-1:12]                  : 
                                                                                            {{32-32{1'b0}},ikiluasjdq}  
                                                  ;


  assign n78yvkhg0miifi58 = (~lkrl_gk1f715er9ueo) ?
          (
            (lgnnlckl1qq6psb & (qndyhstqm8pvl ? 1'b1 : 1'b0)) 
          | (y0nv37yd84l & ( exn_cjm859bpb9zsghqr97 ? 1'b0 : 1'b1))  
          ) : (jp5nha2l14e7kx2jzpke 
          | fpo04urqz74
              )
          ;
  
  
  wire [32-1:0] e98zc_xde8d =  
                           (f8ouikbgg2hqwm8g | ~chhrgp_9_w35oxb) ?      clur09du62kjid[32-1:0]                  :
                           (dvqdxyi_ja1x2 == clur09du62kjid[12]) ?      clur09du62kjid[32-1:0]                  : 
                                                                     {{32-32{1'b0}},ikiluasjdq,clur09du62kjid[11:0]}; 

  wire naka2ay4mdl;
  wire fs1tpvbf2pxudth;
  wire aqs966d99ig8;

  assign naka2ay4mdl                = w66c528fqa9qnfz1btjnm;
  assign hjbzyjew4g2fmth4l66ng8        = e98zc_xde8d[32-1:0];
  assign dl59edtk0_9k5jd65gxp        = qndyhstqm8pvl;
  assign unzbnfwje52jxr_9yt38_bmn       = qj_5hjk5ts;
  assign qtcuhd18j5hjtx41o9tjmv0cm434  = iy42niqez8r3zkja;
  assign srphqbnx3w67orxkuwvoz       = av4ep8dz4xawf95kyr8j;
  assign jbju6a9hecf_f8kg2bsz4       = ynqlvklp9ljiaqdpo;
  
  wire a62b800xjy4edxn_4s8fzk4wgk       = gsoquod_6th_uva & ldn2go4l40668ayimy & (brgdc0amsvlnwf_2j == v_qy6klyvlpd9v); 
  wire pt2d6wjovqmzmmlp43nczy       = gsoquod_6th_uva & (brgdc0amsvlnwf_2j == r10y29zxz4oiu3wd);                 
  wire n59x0nhz5fq5sl52r8zohz12f2       = a62b800xjy4edxn_4s8fzk4wgk | pt2d6wjovqmzmmlp43nczy;
  wire jbh66pmg85o58n2u5jsyhti       = a62b800xjy4edxn_4s8fzk4wgk & (~pt2d6wjovqmzmmlp43nczy);
  ux607_gnrl_dfflr #(1) htrrsmwdvzobd0ds20onffnv(n59x0nhz5fq5sl52r8zohz12f2, jbh66pmg85o58n2u5jsyhti, oa95jvzldxkjxnka5, gf33atgy, ru_wi);































  assign aqs966d99ig8 =   1'b0; 
  assign fs1tpvbf2pxudth =   1'b0; 

  assign vij3v0mhh5pmf2niajrtl =   1'b0 
                                 | (naka2ay4mdl & lgnnlckl1qq6psb) 
                                 ; 

  assign x2n1derqad2ie59_pd542m =   1'b0 
                                 | (aqs966d99ig8 & lgnnlckl1qq6psb) 
                                 ; 

  assign yzrjop7pz8lqhpmcv2wfbrz_u =   1'b0 
                                 | (fs1tpvbf2pxudth & lgnnlckl1qq6psb) 
                                 ; 


  
  
  wc2lipjaiimwuy7fx9zp32mr  lbpbwc1x5lhcs71rg3inpdi1d2xu(
     .e98zc_xde8d   (e98zc_xde8d            ),
     .lms849k     (zelwmbvyieb_h56    ),  
     .dhzk00cwbk (fjk5178vaf1h3l5q9_p)
  );



  cqpjxz2qb247thego6htwvkw_aiu lpcbtkgnuc86ae4xr8g1d9jqhojv_j(
  .f_8ecse5wf0jrndlozy2070bja                       (woq47beoqkpu1um82nv58l1u_hyj4       ),        
  .e4sprh35cvfb6sw6lnskyaga91                    (a1r66jlym5w100htq8lfn_o0rapdf5s    ),
  .qrvtg_49_dmoggu94orq0                        (wqjorkypks0nndgahingvyvil3dvqo        ),         
  .iocew24g1qos_gvi3_r3uoqfdf                        (obokll126527kg6wlw1t6vfh8        ),         
  .qh_y92pv7dp1us9t5wxdmm57                        (msh4030y2dhqf78kyckys0c2ue0ic        ),         
  .cznjry8adajzgi6gkmyr830m_u                        (oebo4piph5o2byr1030bgmb0ye31c6        ),         
  .ugixcggahb26m1glzpuqvpq                        (tlmtrlht_1gsijvzms1twiewyym        ),         
  .vbpz6tidsg3o93kih6nmamlyg9wmr1zz                  (ez_fxjs3_wlsve__62ua9tqsfa6k89twfir  ),   
  .j2dtuvq0m4iir947lery9tpxqwhjj2g3                (p3nsxkqv6seglstz4ge77tdjcngbig0w30rq), 
  .wzqcq7ug3_gv3tuf0o                           (qj_5hjk5ts    ),
  .ng5gq72xr47fw8fztwfo8hw                         (rm1dxjejhq7dh3q5m ), 
  .cmyy3ooatm0bn2s6fv8_r                          (st2zalpx0uf ), 
  .ckgybqpbvuzwgxv1ixd_6rpf                          (ni01kj42oob2x ),
  .nguthky_k_yqsf8fa9btry1                          (ah8kjlmvnaxzbi ),
  .w30ye15yns15                                     (w30ye15yns15 ),
  .jyl_xsaj6z1u9wndwpi                               (sxvvsxtbhyvt ),

  .idg19n7mm21jtb                                  (ynqlvklp9ljiaqdpo ), 
  .o_4mw1alrjmdzl                                 (csz9svan7w77t2lrv3uyj__),
  .nkjxsm02z2_q5_0_                               (hklxc4qx7d75xvdr5e3x9),
  .gf33atgy    (gf33atgy),
  .ru_wi  (ru_wi)
);

  wire fsgnwimjaxqsp7mcuzwf =   csz9svan7w77t2lrv3uyj__ 
                              | hklxc4qx7d75xvdr5e3x9
                              ;
  wire u8glpkklmtu79t083uk6 = lkrl_gk1f715er9ueo | (t_o74lk4v_gxtrgop & woq47beoqkpu1um82nv58l1u_hyj4); 
  wire t3u7iqj1320a4klcqvg09h = lkrl_gk1f715er9ueo ? 1'b0 : fsgnwimjaxqsp7mcuzwf;
  ux607_gnrl_dfflr #(1)   bizlzn55dt3s8lm276267  (u8glpkklmtu79t083uk6,   t3u7iqj1320a4klcqvg09h,   xy7mzrc3a5aq_a, gf33atgy, ru_wi);

  wire bcdn7gznvbqy4hwxscq = lkrl_gk1f715er9ueo | (t_o74lk4v_gxtrgop & woq47beoqkpu1um82nv58l1u_hyj4);
  wire fh9md012gjtyq1oqynef = lkrl_gk1f715er9ueo ? 1'b0 : csz9svan7w77t2lrv3uyj__;
  wire plfnby2dsepbcecrm;
  ux607_gnrl_dfflr #(1)   ag4jxw01msfs0tyj94x3ey1  (bcdn7gznvbqy4hwxscq,   fh9md012gjtyq1oqynef,   plfnby2dsepbcecrm, gf33atgy, ru_wi);

  wire a7zsjlt7lcl8i8olvtf13 = lkrl_gk1f715er9ueo | (t_o74lk4v_gxtrgop & woq47beoqkpu1um82nv58l1u_hyj4);
  wire m1w7hn98n_6_e762y7tjfa = lkrl_gk1f715er9ueo ? 1'b0 : hklxc4qx7d75xvdr5e3x9;
  wire uz6ebmyjnb1u6gootqxy;
  ux607_gnrl_dfflr #(1)   bnilmx6b1gdztiqt742eo8s3uo  (a7zsjlt7lcl8i8olvtf13,   m1w7hn98n_6_e762y7tjfa,   uz6ebmyjnb1u6gootqxy, gf33atgy, ru_wi);




  wire [64-1:0] nx737mdnbv2dflgkm = 
            ({64{lkrl_gk1f715er9ueo}}     & {8{a4a48egkdkec8d9b_9[ 7: 0]}})
          | ({64{dwmx63ax2_grri9q93qee }} & {8{h3p0wpn_ah[15: 8]}}) 
          | ({64{uk63nhcynwa_qtvrcek }} & {8{h3p0wpn_ah[23:16]}}) 
          | ({64{umzor0sgk1r994nu3crx }} & {8{h3p0wpn_ah[31:24]}})
          | ({64{n43zel0f3h8f58krco8e }} & {8{h3p0wpn_ah[39:32]}})
          | ({64{rfes318a1jw5dtuzpbz2 }} & {8{h3p0wpn_ah[47:40]}})
          | ({64{kgdwxspbwxi691glel5lgi6 }} & {8{h3p0wpn_ah[55:48]}})
          | ({64{lfm_3bqoo7ge6c9h9n_pse }} & {8{h3p0wpn_ah[63:56]}})
          ;

  
  
  
  wire [8-1:0] j1qtcyjbuw9dkt5px3 = 8'b00000001 << icfwo5l56zab795f[2:0];
  
          
  
  assign x90uy0klprtqdcq[3:0]   = {4{cfe949_7aiw |!clur09du62kjid[2]}};
  assign x90uy0klprtqdcq[7:4]   = {4{cfe949_7aiw | clur09du62kjid[2]}};
  assign m6uirg1k2s6vd_m8[31:0]  = ttgsydregi0kgoj_z[31:0];
  assign m6uirg1k2s6vd_m8[63:32] =
                         cfe949_7aiw ? ttgsydregi0kgoj_z[63:32] : 
                         ttgsydregi0kgoj_z[31:0];
  assign fn5e7uint162p6axap1i1t9 =      
                          cfe949_7aiw ? gxo5tf4bea2gsq4yyn                   :
                                  clur09du62kjid[2] ? {{32{gxo5tf4bea2gsq4yyn[63]}} , gxo5tf4bea2gsq4yyn[63:32]}  :
                                                    {{32{gxo5tf4bea2gsq4yyn[31]}} , gxo5tf4bea2gsq4yyn[31: 0]}
                                                  ;
  
  
  
  
  

  assign wu02k99r_ok2kjj4u119us = (~lkrl_gk1f715er9ueo) ? (     
      (y0nv37yd84l & exn_cjm859bpb9zsghqr97) ? m6uirg1k2s6vd_m8:  
      qxeco0b4xvxw1v ? nx737mdnbv2dflgkm :
      64'b0)
      : u9y07o_n2vgf1zk ? nx737mdnbv2dflgkm  
          : a4a48egkdkec8d9b_9;

  assign ccwk4o03vlem_hqcccf1g6 = (~lkrl_gk1f715er9ueo) ? (
         
      y0nv37yd84l ? x90uy0klprtqdcq :
      qxeco0b4xvxw1v ? j1qtcyjbuw9dkt5px3 :
      8'b0)
      : u9y07o_n2vgf1zk ? j1qtcyjbuw9dkt5px3  
      : xwfmltfzahuj4qfn4qf2;


  assign yx2bhxvyxmxjggxrsrr833 =
                             ldn2go4l40668ayimy |
                             fpo04urqz74        |
                             a2i6e7_7       |
                                (~lkrl_gk1f715er9ueo);
  
  
  assign qe64ftxd03f_vqrd2sd     = (~lkrl_gk1f715er9ueo) ? (
                   1'b0 
             ) : (
                   fpo04urqz74
                 
			 );
  assign xmbe_e4vm6ofjbn7lq = (oz66a4n0vakndgbkbj6ds & y0nv37yd84l & w0vagcfu1v7wkym9f & b5b1bdkf9u8xkel6mtmr)     
                          | (l2kas5gsiruf5xw6z_b & w0vagcfu1v7wkym9f & b5b1bdkf9u8xkel6mtmr)                    
                          | (syokr6jqxk89zy8h & wh1vvvsvv8tc2elyruo93);                   
                                                                                   
                                                                                   
																				   
																				   
  assign b36sriu021vdo_ujif8     = 
              1'b0;

  assign o1gawztvzi0onzitk     = (~lkrl_gk1f715er9ueo) ? adng7z_1b3srxoxai1rm : oq9b5zfhza9yvdoj;
  assign lr02cqs6anj9gvr45kv    = (~lkrl_gk1f715er9ueo) ? deonbdggc2hhsqq88 : l3c127qdc9a2mfc13;

  assign ltx9lurd9p2ivmnufrgrw     = (~lkrl_gk1f715er9ueo) ? (
                lgnnlckl1qq6psb  ? 2'b0  :
                t6rn2o8trm4jaor9u9i2 ) :
                  
                  
                l_giy79jkzkxy7j ? 2'b0 : 
                ggxoqcj7ytp1a4pjf7ee; 

  assign z6ncd60zcel8m99zg6v     = (~lkrl_gk1f715er9ueo) ? av4ep8dz4xawf95kyr8j  : zdpamqgv7ddf1n3x5t2q ;
  assign st9_is6howar7iysonyyhk     = (~lkrl_gk1f715er9ueo) ? jomllj1p1gxavhm9n  : wpsukhyqhl92dzoam7cm ;
  assign o8407eu9fhzcuymr2a4     = (~lkrl_gk1f715er9ueo) ? ynqlvklp9ljiaqdpo  : v3oo69y614hgiemyyld ;
  assign t3ubula_wguy1a2tut1_e    = (~lkrl_gk1f715er9ueo) ? pf428il3xdc1fkqtfv706k : vy1zc0f0lrbzkonj3v;
  assign ukl6eat4ng6xala4y597l2i    = (~lkrl_gk1f715er9ueo) ? fjk5178vaf1h3l5q9_p : uxlldm0w_h7kicit8gvhqv2;
  assign w3yoivbzacxwr95dw        = (~lkrl_gk1f715er9ueo) ? zelwmbvyieb_h56     : yvu98r_7ji4o250r_u;
                                 


    wn2t_67c13cwq1_8a6 hnddk5wg7l5nzt535efo(
      .ktu3yhilgxp         (1'b0      ),    
      .odfbwv2n0hmkh9n2v     (1'b0      ),
      .vqqbidi8kkzgxc0qls     (1'b0      ),
      .ujg_tx8c5t9t0ddsmq     (1'b0      ),
      .xxf9gqnuyu__15_t1u     (1'b0      ),
      .f4uqn8qf5ljfnqy     (1'b0      ),
      .k0kxgs4dhk1hf26ky3     (1'b0      ),
      .ngw96h2ls51cor4      (1'b0      ),
      .cj5vhekber5gw1509m86     (1'b0      ),
      .zouaj0qk3vke9quhfiqz     (1'b0      ),
      .u3s5vk_sv9c1gjjto    (1'b0      ),
      .pm7lg8nzlruwwz9t29i     (1'b0      ),
      .tffp7jbfj_acgbf_htp    (1'b0      ),
      .mbmpk0lgl7bqaq0m7j    (1'b0      ),
      .fkbmt37lnc1cbn6h7f5q    (1'b0      ),
      .uhs5rs3m1apmo4oj3c7    (1'b0      ),
      .hkzo9ego93d08t8igz2    (1'b0      ),
      .so01tnkdju7vnwezjvi     (64'b0  ),
      .hxad9091n05p_gjjo4     (64'b0  ),
      .uk0gax2bf5vv97rrbosr     (),
           
      .fv0c5k6cjre         (1'b0           ),
      .bm6cerfr_1bou52muqp     (64'b0  ),
      .tz3kfmltx71a5i0tmaln     (64'b0  ),
      .b9asx2rffq8fclg3_q  (1'b0),
      .m1dubsueroj_o4i9hhxf  (1'b0),
      .vupdzhdsf5tcdbcy3br3  (1'b0),
      .rzgzqvqbgh3abztkqck  (1'b0),
      .n9_mxfs9poavrerrqf3ps (1'b0),
      .a8ql4znkrbh_gj7cnnwc2j (1'b0),
      .tz95dh49670qhxle1     (1'b0),
      .ehhimwdiwsd20nyinnomx (),
      .todxu2rm67fxk1x8y_tl4 (),
             
      .yvw7xod98x7         (1'b1           ),
      .tp6hfcjxcyp899mpksjl     (tp6hfcjxcyp899mpksjl       ),
      .f4ds8dbk9kk_ic_     (f4ds8dbk9kk_ic_       ),
      .oso3fj0gx6pnvjni    (oso3fj0gx6pnvjni      ),
      .xl9r7gr7wciuv2d00b     (xl9r7gr7wciuv2d00b       ),
      .htcsb0affil7c6q     (htcsb0affil7c6q       ),
      .vrqdq7uwxf99gj_7      (vrqdq7uwxf99gj_7        ),
      .jqgtsdtxss_uios07     (jqgtsdtxss_uios07       ),
      .hn2h_gkqinydwsdg_i3     (hn2h_gkqinydwsdg_i3       ),
      .re8hncw6m47hrh6     (re8hncw6m47hrh6       ),
      .tshku7fgpiu2j7ugwjj9    (tshku7fgpiu2j7ugwjj9      ),
      .arc8ztjel_qlz3xfw0ya    (arc8ztjel_qlz3xfw0ya      ),
      .dukom1hk2mc9i6m4      (dukom1hk2mc9i6m4        ),
      .ttgsydregi0kgoj_z     (ttgsydregi0kgoj_z       ),

      .e__67e1k5hdb4ctnr    (e__67e1k5hdb4ctnr),
      .jay_5c6ndpwhj0vqzv    (jay_5c6ndpwhj0vqzv),
      .kn6tx97_rw9w0v      (kn6tx97_rw9w0v  ),
                                      
      .nc_3q2q5fz4e2    (nc_3q2q5fz4e2),
      .a5y809wbv8w1d0    (a5y809wbv8w1d0),
      .l0vxn4vg6wd      (l0vxn4vg6wd  ),

      .hgdur8q6gk2ak91b         (1'b0),    
      .r_aei1gc7v37oo9dghv     (1'b0),    
      .d1_eg4gq3uyxdyycybx     (1'b0),    
      .od3rbv8xxz65lrcy     (64'b0),
      .du4qneuo7c4380bw33j     (64'b0),
      .m2s376x2ngd1fz27iofg3yf1 (),
      .f2mrhq1ax6cmfmtx_l5 (),


      .gf33atgy                 (gf33atgy  ),
      .ru_wi               (ru_wi) 
    );


  assign ygvgcd3cyi2ipiz53hbsp = f1g98h1x6en1kemv1;

  assign evji0n54bi8hm_n24uk853qw9c = ee10pomiu8s7j7cn; 
  assign argq10f3h723e0jtlrdbu53       = wqbvx_uqjrfzj8cjke712tpq;
  assign e7iar94ylidlt25a9g9n       = 64'h1000;
  assign qj6kqe1holct34gfb0q9p9a04_alrzg = 1'b0;
  
  assign b0fkq6hghv6az5l_j1j2c12imdd6  = ttgsydregi0kgoj_z[26+27+12-1-1:27+12-1]; 
  assign s9psy03yyyxh7qrmosmb1        = ttgsydregi0kgoj_z[27+12-1:12];                                                     
  assign sqkbogq1h4psprgoosl2lmrpj9_ = {1'b0,wpsukhyqhl92dzoam7cm};
  assign n5gj_lxl9078ky9b2zawd0     = v3oo69y614hgiemyyld;
  assign bmkssziw1_8am7ea6dv         = !jp5nha2l14e7kx2jzpke;
  wire k4rf2zte9ksefekc13puv39a6s = goefkr663a4o90wdkcs60017huc9e | lkrl_gk1f715er9ueo; 
  wire r6cco2stxdjs0ffk5nptnc6r = lkrl_gk1f715er9ueo ? 1'b0 : plfnby2dsepbcecrm;
  wire pmlxiv6_r35q6q5iu1ncmeq4fh = lkrl_gk1f715er9ueo ? 1'b0 : uz6ebmyjnb1u6gootqxy & ~plfnby2dsepbcecrm;
  wire nkf3hnu4g29m_xl6txc7c6omt0xen8 = lkrl_gk1f715er9ueo ? 1'b0 : xy7mzrc3a5aq_a;
  ux607_gnrl_dfflr #(1)   e0zu4xhqo8lcie6hx2         (k4rf2zte9ksefekc13puv39a6s, r6cco2stxdjs0ffk5nptnc6r,        ks33bi5hojtg0te9bl7, gf33atgy, ru_wi); 
  ux607_gnrl_dfflr #(1)   fhpk06uh5268ifmcgjjw3zc4o       (k4rf2zte9ksefekc13puv39a6s, pmlxiv6_r35q6q5iu1ncmeq4fh,      eht8nc5zc5sdbpe9nqr67jeju, gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1)   fdm_ztcnmldfqhpxsn7pc       (k4rf2zte9ksefekc13puv39a6s, nkf3hnu4g29m_xl6txc7c6omt0xen8,      yoop58jcvoblafgy3pvb2bxf, gf33atgy, ru_wi);

endmodule                                      


























module tkyketfhrvq0gmush9p8_myoe (

  input exltui35irvvmodu205vw,

  input [64-1:0] vyxop00ua6vr ,  
  input [64-1:0] p6rw9no76a3m ,  
  input [64-1:0] zowrmckfhx7k5 ,
  input [64-1:0] tvh1llq2i3_y ,  
  input [64-1:0] hfsmpma3 ,

  input sxvvsxtbhyvt,
  input  [64*4-1:0] azll7rq5fab5ou,
  input  [64*4-1:0] n6a0r_0zddzrme8,

  input [8*32-1:0] pcr4upio7_tx37, 
  input [8*1-1:0] uzklqlncpqqm1rav,
  input [8*1-1:0] ortueunvnkx_l5m_j,
  input [8*1-1:0] hwuhtb7ucto_utk56,
  input [8*2-1:0] i1env2kmns7qvvuuc,
  input [8*1-1:0] g3s3vpafvy3i,


  input  rm1dxjejhq7dh3q5m,
  input  rvr30vvllni,
  input  z1cj655u31,
  


  input f29yand0_mv30jc6grvj6, 


  input  [64-1:0] ibc9r3db5iet7,
  input                   h7pglrrhtu6x34l5a21ern,


  
  
  
  
  
  
  
  
  
  
  
  
  
  

  
  
  
  
  

  
  
  
  
  input                                vs6ryzcr0bwqs5so,
  input [32-1:0]               j25ub196dc_agl8oovaex4,
  input                                pi2nokcm8qf7och7l4g,
  input                                c0i0hs5tz64_ce5f0z,
  input                                dmzdczrqcueolg3dzufj_by5rmf,
  input                                a1sqko6fok9qzpbtyuw0,
  input                                bquohubxiv2rsayn62v,
  output                               kqyojh1maxy0x834htg,


  
  
  
  
  input                                oa95jvzldxkjxnka5,
  input [32-1:0]               hjbzyjew4g2fmth4l66ng8,
  input                                dl59edtk0_9k5jd65gxp,
  input                                unzbnfwje52jxr_9yt38_bmn,
  input                                qtcuhd18j5hjtx41o9tjmv0cm434,
  input                                srphqbnx3w67orxkuwvoz,
  input                                jbju6a9hecf_f8kg2bsz4,
  output                               w66c528fqa9qnfz1btjnm,






  input                                q9d7ens0ettrow,

  input                                fl5uzx8oymfa, 
  output                               ypn14jlxvbvoxkesp, 
  input  [48-1:0]     gyb1vfnsiaxnp,
  input  [4-1:0]        elf4ijc6zyn02ua,
  input                                ijrke0oayz6k,
  input                                in937eccpoct,
  input                                kc2beprm1o1chr7jv,
  input                                zhfmvvqqyhe6l74,



  input                               scadliwzjp0l78srd9p    ,

  input [64-1:0] e28x1bh5rb6,

  input                                o0gxucmy66th1ly2om5p,
  output wzqcq7ug3_gv3tuf0o,

  input                                hr0gt1i5t2qzoifxdtx3, 
  input                                tnr82i_e_q5p_n4o9w2cp5,

  input  n3zlo14nquu5l7zf3,
  output a_1o1o8345o28hui,
  output t8p1kh0tvb2ej56s,




  output y86fvwjf6k22ahfluzpt9, 
  input  q4gz66g470k0a1u_kk, 

  output hraqlcavq96j53yrbyif,
  output bf5ypgqi4grkg506x  ,

  output flv4ybjx_fxnt8ahli, 
  output mp50sb0x32pr82qg, 
  output r1mbz1476mmd6eb_2gb,
  output omlfl4p9_5zoeeas3, 
  output    p0e6oiwfprzmn8yx9hsoby9,
  output [64-1:0] ue5tzeds4j8o5wx5zkx,
  output i3fga9mifalr9g_siehz7127f4, 
  output sd8rqg0mey7v6mthfjratzooccvk9,
  output e0srj1jifo6i8ocnkw8xqhp  , 
  output ckrr5bi6ad3t5_60gouyjr9vvpfr,


  input [20-1:0]  u6f8hwzstewuo7nl0iywamw,
  input                            c9k79dqw2z4f63_8lcp4w,
  input                            o_4mw1alrjmdzl,
  input                            nkjxsm02z2_q5_0_,





  output                       o21b8ypt1xiu5ml63d,

  output                       badsf4ksbp3k6p_p5hnj2i, 
  input                        ed4kcy8s9nrisftgx_q, 


  output [32-1:0] bdqo1tgw2_bpi2e8alini, 
  output                       jp5nha2l14e7kx2jzpke,   
  output [64-1:0]      a4a48egkdkec8d9b_9, 
  output [8-1:0]   xwfmltfzahuj4qfn4qf2, 
  output [1:0]                 ggxoqcj7ytp1a4pjf7ee,
  output [4-1:0]oq9b5zfhza9yvdoj,
  output                       l3c127qdc9a2mfc13,
  output                       zdpamqgv7ddf1n3x5t2q,
  output                       wpsukhyqhl92dzoam7cm,
  output                       v3oo69y614hgiemyyld,
  output                       vy1zc0f0lrbzkonj3v,
  output                       uxlldm0w_h7kicit8gvhqv2,
  output                       yvu98r_7ji4o250r_u,
  output [4:0]                 szrgf24or2mbt7w_yleh_vt,   
  output                           an6zohwqn5kwj_tsi4_pczkvu,
  output                           bvvlopjoczq9r7vemdrzz3xd,
  output [64-1:0]          yuloizdmigr7b94rp,


  output  l_giy79jkzkxy7j  ,
  output  cw9xa748nw    ,
  output  x1huhi29x9mco   ,
  output  fpo04urqz74     ,
  output  a2i6e7_7    ,
  output  cque110xwd150_ ,
  output  m705cbtazx7y  ,
  output  etp831o_vh94  ,
  output  w3p1po3pu   ,
  output  nxy2oljfg0lssc  ,
  output  n2s7mr_zvl9k  ,
  output  mzwwsw0h6m1  ,
  output  lydg_n0cr655 ,
  output  tb62wswspbytv ,
  output  [64-1:0]      jttn_e63nm4n4lm9, 
  

  output  yixt0a_xmh    , 
  output  ej7frm_ut9j6y, 
  output  izjeme5aukvcc, 
  output  x5nbgu5ggtet3   , 

  input  [64-1:0] ttgsydregi0kgoj_z,

  input  dw0ku_p4sgs3627wdlt6,
  input  ygvgcd3cyi2ipiz53hbsp,






  input  gf33atgy,
  input  ru_wi
  );


  wire hgt2urny9_9; 
  wire nrxcyc791r8gksao; 

  wire qh14lwju0lrg29;
  wire rla2xv8ay27qlm  ;
  wire es_ankzl9_umwimii; 
  wire jq4n1p1ur; 
  wire egpatz0zaci0;
  wire h2oz0el3g2gltc1lq; 
  wire z_hzjzsz08cfoeut;
  wire [64-1:0] aj4uetnjind0y44r;
  wire djq1y534mfpar9a3_1t; 
  wire h7gvmmsamt7ctj9fg45jb;
  wire o0k24pennw4pm8buv2h6  ; 
  wire h0rjx9lkvgvgzd5q0znib2u;



  wire eqirqpxd2aybmhe839d4725ecig;
  wire [48-1:0] ybrrs0__m1aa00 = gyb1vfnsiaxnp;
  wire fj0lzkw_e2tjj = fl5uzx8oymfa;
  wire pkwcaygsgot_59n1  =  ijrke0oayz6k  ;
  wire vy1aysleh0imu4  =  in937eccpoct  ;
  wire pbjk7minp0n89j  =  kc2beprm1o1chr7jv  ;
  wire b4uk5z2pu_0s =  zhfmvvqqyhe6l74 ;
  wire [64-1:0]bi9zhg2zyeg = ibc9r3db5iet7;
  wire izavxptwkids56szaouo9_zj;
  wire k4zu6hd9_l91sgx;
  wire gp8w0vslru_r_rm7;
  wire o4u5pott58g;




  wire       w12tykr0sjk3cb    = ybrrs0__m1aa00 [5:5   ];
  wire       grfzm3doiudavltu   = ybrrs0__m1aa00 [6:6  ];
  wire       v2mydpki2mkh     = ybrrs0__m1aa00 [11:11    ];
  wire [1:0] i2x6qt_wyuanj  = ybrrs0__m1aa00 [28:27];

  wire [1:0] bwnqxkmv3793tn5    = ybrrs0__m1aa00 [8:7   ];
  wire       a02fqysr32bpia6b   = ybrrs0__m1aa00 [9:9  ];
  wire       m2q3ghpncvh    = ybrrs0__m1aa00 [10:10   ];
  wire       uadexzk_kh0g49nb = ybrrs0__m1aa00 [12:12];
  wire       r8x3j28xrzm0eq  = ybrrs0__m1aa00 [13:13 ];
  wire       m5ljd54icrby7u  = ybrrs0__m1aa00 [14:14 ];
  wire       ola68283_q7l   = ybrrs0__m1aa00 [15:15  ];
  wire       icz9kk4dx5uzjcoz  = ybrrs0__m1aa00 [16:16 ];
  wire       qpjjk_tptwhr4qvkz  = ybrrs0__m1aa00 [17:17 ];
  wire       mhi7m13i4tdp  = ybrrs0__m1aa00 [18:18 ];
  wire       qsexm8gncgpsd0 = ybrrs0__m1aa00 [19:19];
  wire       xsjat4ppp7fq3wj = ybrrs0__m1aa00 [20:20];
  wire       db5c7uyis59qjegezc = ybrrs0__m1aa00 [24:24];
  wire       o12r1q7fso07g4lk = ybrrs0__m1aa00 [22:22];
  wire       z5atnp0pqvut7tu3 = ybrrs0__m1aa00 [23:23];
  wire       my6482rcbzjsl0k = ybrrs0__m1aa00 [25:25];
  wire       foo1r_kdsxld_y28ot5 = ybrrs0__m1aa00 [26:26];

    wire       m7pgd062044v      = 1'b0 
                  ; 
    wire       bcz6wdcu6f4c      = 1'b0 
                  ; 
  wire       d8gxc7jp52uv      = w12tykr0sjk3cb  & (i2x6qt_wyuanj == 2'b10); 
  wire       vmlg53ng6oe      = grfzm3doiudavltu & (i2x6qt_wyuanj == 2'b10); 
  wire       av18nzhvobpoka      = w12tykr0sjk3cb  & (i2x6qt_wyuanj == 2'b11); 
  wire       p08f2oxj96slt      = grfzm3doiudavltu & (i2x6qt_wyuanj == 2'b11); 
  wire       jgah5jfw = m7pgd062044v | bcz6wdcu6f4c | d8gxc7jp52uv | vmlg53ng6oe | av18nzhvobpoka | p08f2oxj96slt;
  wire       bp9qt1h52k23 =  av18nzhvobpoka | p08f2oxj96slt;
  wire       t6ehcvrshdj =  m7pgd062044v | bcz6wdcu6f4c | d8gxc7jp52uv | vmlg53ng6oe;

  wire mus3nlhgqg8z3  = (bwnqxkmv3793tn5 == 2'b00);
  wire wlr32w09idkvg08 = (bwnqxkmv3793tn5 == 2'b01);
  wire csc54ee05lea_  = (bwnqxkmv3793tn5 == 2'b10);
  wire kwx1csxie28n7o  = (bwnqxkmv3793tn5 == 2'b11);

  wire cmxgyc59qlsu3szbo3pn2a = 
            (wlr32w09idkvg08 &  bdqo1tgw2_bpi2e8alini[0])
          | (csc54ee05lea_ &(|bdqo1tgw2_bpi2e8alini[1:0])) 
          | (kwx1csxie28n7o &(|bdqo1tgw2_bpi2e8alini[2:0]))
            ;


  wire jwgi6m_mhsmw95cqy5m1 = cmxgyc59qlsu3szbo3pn2a;

  wire cbalvtbhjuduth_a;

  wire gi5sx4wh1y = (w12tykr0sjk3cb | grfzm3doiudavltu);

  wire joddu4hrozwigoqc8ud = (~jwgi6m_mhsmw95cqy5m1) & gi5sx4wh1y;

  wire bwusl97ottvedusnq = jwgi6m_mhsmw95cqy5m1 & gi5sx4wh1y;

  wire l9_keysot8ddi96l = (jwgi6m_mhsmw95cqy5m1 & v2mydpki2mkh);

  wire ip9a_yuu2kn5f  = v2mydpki2mkh | ((w12tykr0sjk3cb | grfzm3doiudavltu) & m2q3ghpncvh); 
















  assign gp8w0vslru_r_rm7 = a2i6e7_7 | fpo04urqz74 | (l_giy79jkzkxy7j & exltui35irvvmodu205vw);

  assign izavxptwkids56szaouo9_zj = 
                       (
                             (gp8w0vslru_r_rm7  ? (~h7pglrrhtu6x34l5a21ern) : 1'b1)
                           & (gp8w0vslru_r_rm7  ? (~dw0ku_p4sgs3627wdlt6  ) : 1'b1) 
                       );


  assign k4zu6hd9_l91sgx = (uxlldm0w_h7kicit8gvhqv2 ? (~dw0ku_p4sgs3627wdlt6) : 1'b1);


  wire bzelinwijmbrd8ridm =    izavxptwkids56szaouo9_zj  
                         &  k4zu6hd9_l91sgx

                         & (o0gxucmy66th1ly2om5p | c9k79dqw2z4f63_8lcp4w)
                         ;

  wire vjgef0jjjb2bjablf3;
  wire ittjqpuh0jwnzsx9zt;
  wire y5lmpe1pw528nprhwfhjcw198;
  wire kdaater3onb4g112yxh4_1qxd1y;
  wire nnuy7nv12zz86zzsk3v3nlhb2jy;
  wire ztmxn3ljr221cia70thz28_n;
  wire r7bp_0qk912v3lonw6m9pdpilks;
  wire c8p765orxzwimt368eaghlkei;

  assign ypn14jlxvbvoxkesp     = bzelinwijmbrd8ridm & vjgef0jjjb2bjablf3;
  assign ittjqpuh0jwnzsx9zt = bzelinwijmbrd8ridm & fl5uzx8oymfa;

  assign o21b8ypt1xiu5ml63d  = ittjqpuh0jwnzsx9zt;



  assign vjgef0jjjb2bjablf3 = y5lmpe1pw528nprhwfhjcw198 & nrxcyc791r8gksao; 

  assign hgt2urny9_9            = y5lmpe1pw528nprhwfhjcw198 & ittjqpuh0jwnzsx9zt; 
  assign kdaater3onb4g112yxh4_1qxd1y = nrxcyc791r8gksao            & ittjqpuh0jwnzsx9zt;



  assign y5lmpe1pw528nprhwfhjcw198 = o4u5pott58g ? 1'b1 : nnuy7nv12zz86zzsk3v3nlhb2jy;
  assign ztmxn3ljr221cia70thz28_n = o4u5pott58g ? 1'b0 : kdaater3onb4g112yxh4_1qxd1y;





  assign nnuy7nv12zz86zzsk3v3nlhb2jy = gp8w0vslru_r_rm7 ? ygvgcd3cyi2ipiz53hbsp : r7bp_0qk912v3lonw6m9pdpilks;
  assign c8p765orxzwimt368eaghlkei = ztmxn3ljr221cia70thz28_n;

  assign badsf4ksbp3k6p_p5hnj2i = c8p765orxzwimt368eaghlkei;
  assign r7bp_0qk912v3lonw6m9pdpilks = ed4kcy8s9nrisftgx_q;





  wire e8zdez8sbero_ki, oj6_b0zewh20s7p4u;
  zu3cpta_6amki_tj3nyfxw7 do6b96j7qg1pmnqlnbfhoskvn0b(
    
    

    .j2f1_e0en     (pbjk7minp0n89j ),
    .aw82i964do     (pkwcaygsgot_59n1 ),
    .y8_gkxsfle     (vy1aysleh0imu4 ),
    .x6eruzvd5     (yuloizdmigr7b94rp      ),
    .kw2010ymt1iz5   (w12tykr0sjk3cb  ),
    .yeo38qe8mley55  (grfzm3doiudavltu ),
    .rvfxw53dft5    (v2mydpki2mkh   ),
    .r6dop3ru22     (1'b0   ),
    .n6a0r_0zddzrme8 (n6a0r_0zddzrme8),
    .azll7rq5fab5ou (azll7rq5fab5ou),

    .coeuovgdaw1  (e8zdez8sbero_ki  ),
    .o_gen1so7__xgr3pw2(oj6_b0zewh20s7p4u),
    .gf33atgy(gf33atgy),
    .ru_wi(ru_wi)
  );


  assign djq1y534mfpar9a3_1t   = e8zdez8sbero_ki  ;
  assign h7gvmmsamt7ctj9fg45jb = oj6_b0zewh20s7p4u;
  assign cbalvtbhjuduth_a = (h7gvmmsamt7ctj9fg45jb | djq1y534mfpar9a3_1t);

  assign aj4uetnjind0y44r = yuloizdmigr7b94rp;







  assign wzqcq7ug3_gv3tuf0o = v2mydpki2mkh | grfzm3doiudavltu;

  wire ebfq97xvdduyndg280qv;

  wire cler8gtj8253s3ld = v2mydpki2mkh | w12tykr0sjk3cb;
  wire zm5_ofuijsle46r = v2mydpki2mkh | grfzm3doiudavltu;

  
  
  
  wire qszb2sk2j_j82swem1 = 
                          vs6ryzcr0bwqs5so  ?  pi2nokcm8qf7och7l4g  :
                          
                          oa95jvzldxkjxnka5 ?  dl59edtk0_9k5jd65gxp :
                          cler8gtj8253s3ld;

  wire p_abbxlz8g37sezzdiz = 
                          vs6ryzcr0bwqs5so  ?  c0i0hs5tz64_ce5f0z  :
                          
                          oa95jvzldxkjxnka5 ?  unzbnfwje52jxr_9yt38_bmn :
                          zm5_ofuijsle46r;

  wire xztklfbn7v2ii3v_uevlo3r  = 
                          vs6ryzcr0bwqs5so  ?  dmzdczrqcueolg3dzufj_by5rmf  :
                          
                          oa95jvzldxkjxnka5 ?  qtcuhd18j5hjtx41o9tjmv0cm434 :
                          rvr30vvllni;

  wire xd167z8s0v_0qz__0jw86       = 
                          vs6ryzcr0bwqs5so  ?  a1sqko6fok9qzpbtyuw0  :
                          
                          oa95jvzldxkjxnka5 ?  srphqbnx3w67orxkuwvoz :
                          pkwcaygsgot_59n1;

  wire i05xjlghmnn2qbrl28vz       = 
                          vs6ryzcr0bwqs5so  ?  bquohubxiv2rsayn62v  :
                          
                          oa95jvzldxkjxnka5 ?  jbju6a9hecf_f8kg2bsz4 :
                          v3oo69y614hgiemyyld;

  wire [32-1:0] f1oe4mvkdfixfa21sr  = 
                          vs6ryzcr0bwqs5so  ?  j25ub196dc_agl8oovaex4  :
                          
                          oa95jvzldxkjxnka5 ?  hjbzyjew4g2fmth4l66ng8 :
                          bdqo1tgw2_bpi2e8alini;
  
  wire bmo63m4ok3ua6te7alj1bvii;

  d7stl61zflp21cls1tg tm9w0cgdh85kersg7vk9 (
      .sxvvsxtbhyvt    (sxvvsxtbhyvt),
      .pcr4upio7_tx37     (pcr4upio7_tx37   ), 
      .uzklqlncpqqm1rav  (uzklqlncpqqm1rav),
      .ortueunvnkx_l5m_j  (ortueunvnkx_l5m_j),
      .hwuhtb7ucto_utk56  (hwuhtb7ucto_utk56),
      .i1env2kmns7qvvuuc  (i1env2kmns7qvvuuc),
      .g3s3vpafvy3i  (g3s3vpafvy3i),

      .rm1dxjejhq7dh3q5m  (rm1dxjejhq7dh3q5m ),
      .xatytj_r0fv14q  (xztklfbn7v2ii3v_uevlo3r),

      .oily7    (qszb2sk2j_j82swem1),
      .ly3dor8    (p_abbxlz8g37sezzdiz),
      .p1m    (1'b0),

      .u2k4dyp52s_m(xd167z8s0v_0qz__0jw86 ),
      .bktu0z1mk56(i05xjlghmnn2qbrl28vz ),
      .e98zc_xde8d (f1oe4mvkdfixfa21sr  ),
      .foj6m18  (bmo63m4ok3ua6te7alj1bvii)
  );

  
  
  assign ebfq97xvdduyndg280qv = bmo63m4ok3ua6te7alj1bvii
                             & ~oa95jvzldxkjxnka5
                               ;

  assign  w66c528fqa9qnfz1btjnm = bmo63m4ok3ua6te7alj1bvii;

  assign  kqyojh1maxy0x834htg  = bmo63m4ok3ua6te7alj1bvii;
  









  assign es_ankzl9_umwimii = (1'b0
                       | l9_keysot8ddi96l 
                       | (bwusl97ottvedusnq & m2q3ghpncvh) 



              
                       | (exltui35irvvmodu205vw ? 1'b0 : bwusl97ottvedusnq)
                       )
                       ;

  wire gofn7tjm6he2;   
  assign eqirqpxd2aybmhe839d4725ecig = (o_4mw1alrjmdzl || nkjxsm02z2_q5_0_ 
                                   ) && c9k79dqw2z4f63_8lcp4w && !an6zohwqn5kwj_tsi4_pczkvu;
  assign z_hzjzsz08cfoeut =  (   
                                 o_4mw1alrjmdzl && !an6zohwqn5kwj_tsi4_pczkvu
                               )
                              & (~cbalvtbhjuduth_a)
                              
                              & (~es_ankzl9_umwimii)
                              ;

  assign h2oz0el3g2gltc1lq =  (    
                                  (   ebfq97xvdduyndg280qv  
                                  )
                               && !eqirqpxd2aybmhe839d4725ecig
                             || (nkjxsm02z2_q5_0_ && !an6zohwqn5kwj_tsi4_pczkvu)
                             )
                           & (~cbalvtbhjuduth_a)
                           
                           & (~es_ankzl9_umwimii)
                           & ~(z_hzjzsz08cfoeut)
                           ;



  assign o4u5pott58g = 1'b0
                     | cbalvtbhjuduth_a 
                     
                     | es_ankzl9_umwimii
                     | h2oz0el3g2gltc1lq
                     | z_hzjzsz08cfoeut



                     ;



  assign qh14lwju0lrg29 = 1'b0    

                        | (o4u5pott58g)

                        | (gp8w0vslru_r_rm7)
                        ;

  assign rla2xv8ay27qlm = 1'b0

                      | (gi5sx4wh1y & (~o4u5pott58g))

                      | (o4u5pott58g)

                      ;




  assign jq4n1p1ur      = w12tykr0sjk3cb;
  assign egpatz0zaci0   = grfzm3doiudavltu | v2mydpki2mkh;







  wire jr7bt1u761z2ss2hqtdtx9t9 = bwusl97ottvedusnq | v2mydpki2mkh | o4u5pott58g | m2q3ghpncvh;
  wire q78o6nh9n7wmaov7db8 = (~grfzm3doiudavltu) & (~jr7bt1u761z2ss2hqtdtx9t9);


































  
  assign bvvlopjoczq9r7vemdrzz3xd = !o0gxucmy66th1ly2om5p && 
                                  (   wlr32w09idkvg08 && (&bdqo1tgw2_bpi2e8alini[11:1] && |bdqo1tgw2_bpi2e8alini[0:0])
                                   || csc54ee05lea_  && (&bdqo1tgw2_bpi2e8alini[11:2] && |bdqo1tgw2_bpi2e8alini[1:0])
                                   || kwx1csxie28n7o  && (&bdqo1tgw2_bpi2e8alini[11:3] && |bdqo1tgw2_bpi2e8alini[2:0])
                                  );
  assign yuloizdmigr7b94rp   = ttgsydregi0kgoj_z[64-1:0];
  assign bdqo1tgw2_bpi2e8alini = o0gxucmy66th1ly2om5p ? yuloizdmigr7b94rp[32-1:0] : {u6f8hwzstewuo7nl0iywamw, yuloizdmigr7b94rp[11:0]};
  assign an6zohwqn5kwj_tsi4_pczkvu = o0gxucmy66th1ly2om5p;

  assign jp5nha2l14e7kx2jzpke = w12tykr0sjk3cb; 



  wire [64-1:0] n7ku2x7js0auxoew_ = 
            ({64{mus3nlhgqg8z3 }} & {8{bi9zhg2zyeg[ 7:0]}})
          | ({64{wlr32w09idkvg08}} & {4{bi9zhg2zyeg[15:0]}})
          | ({64{csc54ee05lea_ }} & {2{bi9zhg2zyeg[31:0]}})
          | ({64{kwx1csxie28n7o}}  & ( 
                                   db5c7uyis59qjegezc ? vyxop00ua6vr :  
                                   z5atnp0pqvut7tu3 ? p6rw9no76a3m :  
                                   foo1r_kdsxld_y28ot5 ? tvh1llq2i3_y :  
                                   o12r1q7fso07g4lk ?  zowrmckfhx7k5 :
                                   my6482rcbzjsl0k ?  hfsmpma3 :
                                              bi9zhg2zyeg[63:0]))
          ;


  wire [8-1:0] afztve62tee2r1 = 
            ({8{mus3nlhgqg8z3 }} & (8'b00000001 << bdqo1tgw2_bpi2e8alini[2:0]))
          | ({8{wlr32w09idkvg08}} & (8'b00000011 <<{bdqo1tgw2_bpi2e8alini[2:1],1'b0}))
          | ({8{csc54ee05lea_ }} & (8'b00001111 <<{bdqo1tgw2_bpi2e8alini[2  ],2'b0})) 
          | ({8{kwx1csxie28n7o }} & (8'b11111111));

  wire [64-1:0] rfzk0egtlh9={64{1'b0}}; 
  

  assign                szrgf24or2mbt7w_yleh_vt   = 5'b0;

  wire [64-1:0] vj7eqf1xjt6w49h6act = 
            (
               ({64{csc54ee05lea_ }} & {2{bi9zhg2zyeg[31:0]}}) 
             | ({64{kwx1csxie28n7o }} & bi9zhg2zyeg)
            );

  wire [8-1:0] o3g9z219e1_kgj7s0o4qt = 
            ({8{csc54ee05lea_ }} & (8'b0000_1111 << {bdqo1tgw2_bpi2e8alini[2],2'b0}))
          | ({8{kwx1csxie28n7o }} & (8'b1111_1111))
          ;

  assign a4a48egkdkec8d9b_9 =
                             jgah5jfw ? vj7eqf1xjt6w49h6act : 
                               n7ku2x7js0auxoew_
                           ;
  assign xwfmltfzahuj4qfn4qf2 = 
                             jgah5jfw ? o3g9z219e1_kgj7s0o4qt : 
                               afztve62tee2r1
                           ;


  assign oq9b5zfhza9yvdoj     = elf4ijc6zyn02ua;
  assign l3c127qdc9a2mfc13    = a02fqysr32bpia6b;
  assign ggxoqcj7ytp1a4pjf7ee     = bwnqxkmv3793tn5;
  assign v3oo69y614hgiemyyld     = pbjk7minp0n89j;
  assign vy1zc0f0lrbzkonj3v    = b4uk5z2pu_0s;


  wire fwmbk3wv_1qt = 
                (pbjk7minp0n89j ? sxvvsxtbhyvt : 1'b1) &
                 rm1dxjejhq7dh3q5m;

  wire y_yl6g1vnk = (fwmbk3wv_1qt) ? rvr30vvllni : (pkwcaygsgot_59n1 | pbjk7minp0n89j);

  assign zdpamqgv7ddf1n3x5t2q     = y_yl6g1vnk;

  
  wire kfjdozrxmb = (fwmbk3wv_1qt) ? z1cj655u31 : (vy1aysleh0imu4 & (~pbjk7minp0n89j));
  
  assign wpsukhyqhl92dzoam7cm     = kfjdozrxmb;

  assign  l_giy79jkzkxy7j  = jwgi6m_mhsmw95cqy5m1;
  assign  cw9xa748nw    = w12tykr0sjk3cb;
  assign  x1huhi29x9mco   = grfzm3doiudavltu;

  assign  fpo04urqz74     = v2mydpki2mkh     ;
  assign  a2i6e7_7    = m2q3ghpncvh    ;
  assign  cque110xwd150_ = uadexzk_kh0g49nb ;
  assign  m705cbtazx7y  = r8x3j28xrzm0eq  ;
  assign  etp831o_vh94  = m5ljd54icrby7u  ;
  assign  w3p1po3pu   = ola68283_q7l   ;
  assign  nxy2oljfg0lssc  = icz9kk4dx5uzjcoz  ;
  assign  n2s7mr_zvl9k  = qpjjk_tptwhr4qvkz  ;
  assign  mzwwsw0h6m1  = mhi7m13i4tdp  ;
  assign  lydg_n0cr655 = qsexm8gncgpsd0 ;
  assign  tb62wswspbytv = xsjat4ppp7fq3wj ;
  assign  jttn_e63nm4n4lm9 = bi9zhg2zyeg[64-1:0]; 

  assign yixt0a_xmh     = m7pgd062044v;
  assign ej7frm_ut9j6y = bp9qt1h52k23; 
  assign izjeme5aukvcc = t6ehcvrshdj; 
  assign x5nbgu5ggtet3    = jgah5jfw; 



  wc2lipjaiimwuy7fx9zp32mr  lbpbwc1x5lhcs71rg3inpdi1d2xu(
     .e98zc_xde8d   (bdqo1tgw2_bpi2e8alini),
     .lms849k     (yvu98r_7ji4o250r_u),  
     .dhzk00cwbk (uxlldm0w_h7kicit8gvhqv2)
  );





























  assign o0k24pennw4pm8buv2h6   = hr0gt1i5t2qzoifxdtx3  ;
  assign h0rjx9lkvgvgzd5q0znib2u = tnr82i_e_q5p_n4o9w2cp5;
  assign gofn7tjm6he2 = o0k24pennw4pm8buv2h6 | h0rjx9lkvgvgzd5q0znib2u;





  localparam ofr49_k0kstw57 = (
                        6
                       +1
                       +64
                       +4
                       );

  wire [ofr49_k0kstw57-1:0] vqvk5be0ew5;
  wire [ofr49_k0kstw57-1:0] uo1dbdf4eec96ry191bf;





  assign vqvk5be0ew5 = {
         qh14lwju0lrg29 
       , rla2xv8ay27qlm   
       , es_ankzl9_umwimii
       , jq4n1p1ur
       , egpatz0zaci0
       , h2oz0el3g2gltc1lq
       , z_hzjzsz08cfoeut
       , aj4uetnjind0y44r
       , djq1y534mfpar9a3_1t
       , h7gvmmsamt7ctj9fg45jb
       , o0k24pennw4pm8buv2h6  
       , h0rjx9lkvgvgzd5q0znib2u
       };

  assign {
         hraqlcavq96j53yrbyif 
       , bf5ypgqi4grkg506x   
       , flv4ybjx_fxnt8ahli
       , mp50sb0x32pr82qg
       , r1mbz1476mmd6eb_2gb
       , omlfl4p9_5zoeeas3
       , p0e6oiwfprzmn8yx9hsoby9
       , ue5tzeds4j8o5wx5zkx
       , i3fga9mifalr9g_siehz7127f4
       , sd8rqg0mey7v6mthfjratzooccvk9
       , e0srj1jifo6i8ocnkw8xqhp  
       , ckrr5bi6ad3t5_60gouyjr9vvpfr
       } = uo1dbdf4eec96ry191bf;


















































  assign uo1dbdf4eec96ry191bf = vqvk5be0ew5;
  assign y86fvwjf6k22ahfluzpt9 = hgt2urny9_9;
  assign nrxcyc791r8gksao      = q4gz66g470k0a1u_kk;

  assign a_1o1o8345o28hui   = y86fvwjf6k22ahfluzpt9 & q4gz66g470k0a1u_kk & q78o6nh9n7wmaov7db8;
  assign t8p1kh0tvb2ej56s = n3zlo14nquu5l7zf3;

endmodule                                      

























module iluwktw0594417cwb1su(





  input  fj5f6r_brv9, 
  output kdpypaw_l038t, 

  input  [64-1:0] tcdcik4o5zc,
  input  [64-1:0] d4lx9_3xlxjia1,
  input  [64-1:0] pa1go4rk4_,
  input  [64-1:0] nl8lrzq7,
  input  [34-1:0] h1ieg8rrdd,




  output c4znhmchls2i9, 
  input  fjclz58zhz4y4uf, 

  output [64-1:0] e0lrg61pa8jctwey_k,
  output [64-1:0] ldicihngwys9frt8r_q,
  input  [64-1:0] dytd_hd42_wbyvlhrmt9r7, 
  output ye3uidmavh9jbm9w4,
  output ulpu2wlvtk0b4i,

  output rb8jt7db79k4r076h,
  output g4gfgb2tm_ujg9dhex,
  output vyp0v8hghszoph ,
  output uzn0rxbzurqxprl ,
  output rz9jowsqb1lne29t6, 
  output uo8rfftroteg2gy267f,
  output h8j00pdvikgalx01_,
  output fxpfb14s16dp6ihm,
  output njgro75dfrjo_60y,
  output djpeelru7ruovogpcwr,
  output f8c0swke1b88ml,
  output hmbu9tiu4cl764c,

  output  v3e6l1k7eo9k3 ,
  output  hxrmt706n071lic0f7,







  output [64-1:0] bm6cerfr_1bou52muqp,
  output [64-1:0] tz3kfmltx71a5i0tmaln,
  output b9asx2rffq8fclg3_q ,
  output m1dubsueroj_o4i9hhxf ,
  output vupdzhdsf5tcdbcy3br3 ,
  output rzgzqvqbgh3abztkqck ,
  output n9_mxfs9poavrerrqf3ps,
  output a8ql4znkrbh_gj7cnnwc2j,
  output tz95dh49670qhxle1,

  input  ehhimwdiwsd20nyinnomx,
  input  [64-1:0] todxu2rm67fxk1x8y_tl4,

  input  gf33atgy,
  input  ru_wi
  );


  wire ux9e0dc   = h1ieg8rrdd [17:17 ]; 
  wire i6wn18or   = h1ieg8rrdd [18:18 ]; 
  wire b2nbojhb0   = h1ieg8rrdd [19:19 ]; 
  wire l64obb69 = h1ieg8rrdd [21:21 ]; 
  wire iqfzb2 = h1ieg8rrdd [22:22 ]; 
  wire k8p    = h1ieg8rrdd [16:16 ]; 
  wire fa2_s    = h1ieg8rrdd [5:5]; 
  wire u_vskhg4r   = h1ieg8rrdd [6:6]; 
  wire r0drxtm    = h1ieg8rrdd [8:8];
  wire d1v_   = h1ieg8rrdd [7:7];
  wire vlfahv69   = h1ieg8rrdd [4:4]; 

  wire zdfkhxahx = fa2_s | u_vskhg4r;

  wire fik76hef_4pi = h1ieg8rrdd [9:9 ];

  assign bm6cerfr_1bou52muqp = zdfkhxahx ? nl8lrzq7 : d4lx9_3xlxjia1;
  assign tz3kfmltx71a5i0tmaln = zdfkhxahx ? (vlfahv69 ? 64'd4 : 64'd2)
                                : pa1go4rk4_;

  wire [64-1:0] j5u33aiz66p_mnwyynoh = (k8p | fa2_s) ? nl8lrzq7 : d4lx9_3xlxjia1[64-1:0]; 
  wire [64-1:0] rbtx5k_3xjihbod8o =  tcdcik4o5zc[64-1:0]; 
  wire [64-1:0] k5gbfi75ml5lke9sjzauk5 = j5u33aiz66p_mnwyynoh + rbtx5k_3xjihbod8o;

  wire  crqdad2xg75t5dzsc;

  as9e9kibsg2lccbbj9#(64) ig0hk2uvk971tvgecb
  (   .ta7wib(j5u33aiz66p_mnwyynoh), 
      .g35wi_(rbtx5k_3xjihbod8o), 
      .h_kg5l(dytd_hd42_wbyvlhrmt9r7), 
      .ig1wj(crqdad2xg75t5dzsc), 
      .gf33atgy(gf33atgy), 
      .ru_wi(ru_wi)
  );

  assign ye3uidmavh9jbm9w4 = ~crqdad2xg75t5dzsc;

  assign rb8jt7db79k4r076h = k8p | zdfkhxahx;
  assign g4gfgb2tm_ujg9dhex = u_vskhg4r;
  assign vyp0v8hghszoph  = fa2_s ;
  assign uzn0rxbzurqxprl  = r0drxtm;
  assign rz9jowsqb1lne29t6 = d1v_;
  assign uo8rfftroteg2gy267f = ux9e0dc;
  assign h8j00pdvikgalx01_ = i6wn18or;
  assign fxpfb14s16dp6ihm = b2nbojhb0;
  assign njgro75dfrjo_60y = l64obb69;
  assign djpeelru7ruovogpcwr = iqfzb2;

  assign b9asx2rffq8fclg3_q  = h1ieg8rrdd [10:10  ]  
                             ;
  assign m1dubsueroj_o4i9hhxf  = h1ieg8rrdd [11:11  ]  
                             ;
  assign vupdzhdsf5tcdbcy3br3  = h1ieg8rrdd [12:12  ]; 
  assign rzgzqvqbgh3abztkqck  = h1ieg8rrdd [13:13  ]; 
  assign n9_mxfs9poavrerrqf3ps = h1ieg8rrdd [14:14 ]; 
  assign a8ql4znkrbh_gj7cnnwc2j = h1ieg8rrdd [15:15 ]; 




  assign tz95dh49670qhxle1  = zdfkhxahx;

  assign c4znhmchls2i9     = fj5f6r_brv9;
  assign kdpypaw_l038t     = fjclz58zhz4y4uf;
  assign f8c0swke1b88ml  = fik76hef_4pi;
  assign hmbu9tiu4cl764c  = 
                           zdfkhxahx ? 1'b1 : ehhimwdiwsd20nyinnomx;

  assign e0lrg61pa8jctwey_k  = todxu2rm67fxk1x8y_tl4;
  assign ldicihngwys9frt8r_q = k5gbfi75ml5lke9sjzauk5[64-1:0];
  assign ulpu2wlvtk0b4i   = 1'b0;

  assign v3e6l1k7eo9k3   = c4znhmchls2i9 & fjclz58zhz4y4uf & k8p;
  assign hxrmt706n071lic0f7  = ehhimwdiwsd20nyinnomx & k8p;














endmodule


















module xnt41w1r9gyu7e7lcjxkg92u(
  input  tywculgjyor8ndw,
  input  w2h8uh3l463qbgqmv,

  input  aw82i964do,
  input  y8_gkxsfle,
  input  pydatzxqqi,





  input  v7t8ipf7s3pkl, 
  output r30egqbrycq6277u, 

  input  [64-1:0] uhp5bzs36,
  input  [27-1:0] nybrz2cz78r,
  input  gr47f0gunxy4e1c,   

  output rb050tnl,
  output a94vd35etec4,
  output el7_p8jit09,
  output [12-1:0] e1go3iu,

  input  r0s7d8cr68i2qs1z,
  input  [64-1:0] l9erxxpnphqd26vg9,
  input  [64-1:0] hig2gwwbeuhnt65xrp,
  output [64-1:0] guuvp01vkcryglsu1p3,
  output [64-1:0] vf5xcr67bqhzlo43_,
  input  [64-1:0] zmfo8cca_77pc,
  output [64-1:0] bj7h5jqg66r51jxki6emra,

  output [64-1:0] vmx1fh4kmh4c,








  output wykc_imin5w, 
  input  xnta372agn8z7, 

  output [64-1:0] b6nv94op09myrtj3wy,
  output vp2vijaywqexo22ty08,   


  input  gf33atgy,
  input  ru_wi
  );






  assign wykc_imin5w      = v7t8ipf7s3pkl
                          ;


  assign r30egqbrycq6277u      = 
                             xnta372agn8z7
                           ; 

  assign vp2vijaywqexo22ty08   = r0s7d8cr68i2qs1z;
  assign b6nv94op09myrtj3wy  = 
                          l9erxxpnphqd26vg9
                          ;



  wire        wgp51487  = nybrz2cz78r[5:5 ];
  wire        puf_lwtj  = nybrz2cz78r[6:6 ];
  wire        klxytl1  = nybrz2cz78r[7:7 ];
  wire        dimd95ll = nybrz2cz78r[8:8];
  wire        m5zuks2mif = nybrz2cz78r[14:14];
  wire [4:0]  gjzlds   = nybrz2cz78r[13:9 ];
  wire [11:0] ve4o616ogbq = nybrz2cz78r[26:15];

  assign vmx1fh4kmh4c = dimd95ll ? {27'b0,gjzlds} : uhp5bzs36;

  assign el7_p8jit09 = v7t8ipf7s3pkl & 
    (
      (wgp51487 ? gr47f0gunxy4e1c : 1'b0) 
      | puf_lwtj | klxytl1 
     );
  assign a94vd35etec4 = v7t8ipf7s3pkl & (
                wgp51487 
               | ((puf_lwtj | klxytl1) & (~m5zuks2mif)) 
            );                                                                           

  assign e1go3iu = ve4o616ogbq;
  assign rb050tnl = wykc_imin5w & xnta372agn8z7 
                    & (~tywculgjyor8ndw);

  assign vf5xcr67bqhzlo43_ = 
              ({64{wgp51487}} & vmx1fh4kmh4c)
            | ({64{puf_lwtj}} & (  vmx1fh4kmh4c  | l9erxxpnphqd26vg9))
            | ({64{klxytl1}} & ((~vmx1fh4kmh4c) & l9erxxpnphqd26vg9));

  assign guuvp01vkcryglsu1p3 = 
              ({64{wgp51487}} & vmx1fh4kmh4c)
            | ({64{puf_lwtj}} & (  vmx1fh4kmh4c  | hig2gwwbeuhnt65xrp))
            | ({64{klxytl1}} & ((~vmx1fh4kmh4c) & hig2gwwbeuhnt65xrp));

  assign bj7h5jqg66r51jxki6emra = 
              ({64{wgp51487}} & vmx1fh4kmh4c)
            | ({64{puf_lwtj}} & (  vmx1fh4kmh4c  | zmfo8cca_77pc))
            | ({64{klxytl1}} & ((~vmx1fh4kmh4c) & zmfo8cca_77pc));

endmodule



















module wn2t_67c13cwq1_8a6(



  input  ktu3yhilgxp,

  input  odfbwv2n0hmkh9n2v ,
  input  vqqbidi8kkzgxc0qls ,
  input  ujg_tx8c5t9t0ddsmq ,
  input  xxf9gqnuyu__15_t1u ,
  input  f4uqn8qf5ljfnqy ,
  input  k0kxgs4dhk1hf26ky3 ,
  input  ngw96h2ls51cor4  ,
  input  cj5vhekber5gw1509m86 ,
  input  zouaj0qk3vke9quhfiqz ,
  input  u3s5vk_sv9c1gjjto,
  input  pm7lg8nzlruwwz9t29i ,
  input  [64-1:0] so01tnkdju7vnwezjvi,
  input  [64-1:0] hxad9091n05p_gjjo4,
  input tffp7jbfj_acgbf_htp  ,
  input mbmpk0lgl7bqaq0m7j  ,
  input fkbmt37lnc1cbn6h7f5q  ,
  input uhs5rs3m1apmo4oj3c7  ,
  input hkzo9ego93d08t8igz2  ,
  
  
  
  


  output [64-1:0] uk0gax2bf5vv97rrbosr,



  input  fv0c5k6cjre,

  input  [64-1:0] bm6cerfr_1bou52muqp,
  input  [64-1:0] tz3kfmltx71a5i0tmaln,
  input  b9asx2rffq8fclg3_q ,
  input  m1dubsueroj_o4i9hhxf ,
  input  vupdzhdsf5tcdbcy3br3 ,
  input  rzgzqvqbgh3abztkqck ,
  input  n9_mxfs9poavrerrqf3ps,
  input  a8ql4znkrbh_gj7cnnwc2j,
  input  tz95dh49670qhxle1,

  output ehhimwdiwsd20nyinnomx,
  output [64-1:0] todxu2rm67fxk1x8y_tl4,



  input  yvw7xod98x7,

  input  [64-1:0] tp6hfcjxcyp899mpksjl,
  input  [64-1:0] f4ds8dbk9kk_ic_,
  input  oso3fj0gx6pnvjni,
  input  xl9r7gr7wciuv2d00b ,
  input  htcsb0affil7c6q ,
  input  vrqdq7uwxf99gj_7  ,
  input  jqgtsdtxss_uios07 ,
  input  hn2h_gkqinydwsdg_i3 ,
  input  re8hncw6m47hrh6 ,
  input  tshku7fgpiu2j7ugwjj9,
  input  arc8ztjel_qlz3xfw0ya,
  input  dukom1hk2mc9i6m4,
  output [64-1:0] ttgsydregi0kgoj_z,

  input  e__67e1k5hdb4ctnr,
  input  [64-1:0] jay_5c6ndpwhj0vqzv,
  output [64-1:0] kn6tx97_rw9w0v,

  input  nc_3q2q5fz4e2,
  input  [64-1:0] a5y809wbv8w1d0,
  output [64-1:0] l0vxn4vg6wd,


  
  
  input  hgdur8q6gk2ak91b,
  input  r_aei1gc7v37oo9dghv,
  input  d1_eg4gq3uyxdyycybx,
  input  [64-1:0] od3rbv8xxz65lrcy,
  input  [64-1:0] du4qneuo7c4380bw33j,
  output [64-1:0] m2s376x2ngd1fz27iofg3yf1,
  output [64-1:0] f2mrhq1ax6cmfmtx_l5,

  input  gf33atgy,
  input  ru_wi
  );









       

  wire [64-1:0] az6qlcqsx_0;
  wire [64-1:0] cqqzeukmh;

  wire [64-1:0] yxz3vex1f = az6qlcqsx_0[64-1:0];
  wire [64-1:0] afthitl2 = cqqzeukmh[64-1:0];


  wire [64-1:0] svtp9g_orl2 = 
          hgdur8q6gk2ak91b ? od3rbv8xxz65lrcy : 
          so01tnkdju7vnwezjvi[64-1:0];
  wire [64-1:0] ovco_g1rr8cl = 
          hgdur8q6gk2ak91b ? du4qneuo7c4380bw33j : 
          hxad9091n05p_gjjo4[64-1:0];

  wire b1vnk2xf9;  
  wire nsc05do ; 
  wire cod1y7dl_;
  wire e7pwgmzzw54;

  wire mf5fcnu2azr;
  wire m0mq6jm4ys;
  wire uv65k1vtj = mf5fcnu2azr | m0mq6jm4ys; 

  wire zjk3uzc5cf;
  wire obmd5e6;
  wire qi__zhsq1zl9o_w = zjk3uzc5cf | obmd5e6; 

  wire nynmmk;
  wire oss8f_hhqe8;
  wire tqvnzdez;

  wire onsk4u1y9_e;
  wire tdz9d9;
  wire jxe3dht;

  wire b9bqr_g01;
  wire t1f2vol;
  wire w23f72vq40;

  wire fy1ybps5;
  wire q0brgn6;

  wire x1_dx841;


  wire g8dm1b58pm6xt ;
  wire bqmj8280_l ;
  wire egmgssvj3 ;
  wire nssum1cfr ;
  wire rn573wyhxlx2330;
  wire fm3pgkuczco;

  wire ufa33rbvjwk;

  wire t6d11eqb1s3;
  wire [64+1-1:0] yoibsjp7ouplcq;
  wire [64+1-1:0] tawrhvnsab;

  wire em10uopmr98x;
  wire [64+1-1:0] iajwu4x_2;
  wire [64+1-1:0] o7xczhh6fe;






  wire [64-1:0] eaks5rrtzx4;
  wire [6-1:0] qkr7a25rdze;
  wire [64-1:0] cvnvrq3lozc;

  wire [64-1:0]  rckctyqlnspj0, osmygk9ar45_; 
  genvar i;
  generate
    for (i=0;i<64;i=i+1) begin:ctx1tim9yd_vkndxkpsf8_9u
      if (i<32) begin :xqrf9su1zd
      assign rckctyqlnspj0[i] = (t1f2vol|w23f72vq40)? 1'b0 : svtp9g_orl2[64-1-i]; 
      end
      else begin :t3v_vnx8apzi6d
      assign rckctyqlnspj0[i] = svtp9g_orl2[64-1-i]; 
      end
      assign osmygk9ar45_[i] = cvnvrq3lozc[64-1-i]; 
    end
  endgenerate



  wire j4qv5sod = jxe3dht | onsk4u1y9_e | tdz9d9
                     | b9bqr_g01 | t1f2vol | w23f72vq40 
                  ; 
  wire bj8rlymm54x = 1'b0
                       | b9bqr_g01 | t1f2vol | w23f72vq40 
                     ; 



















  assign eaks5rrtzx4 = {64{j4qv5sod}} &
           ((jxe3dht | tdz9d9 | t1f2vol | w23f72vq40) ? rckctyqlnspj0 : svtp9g_orl2);
  assign qkr7a25rdze[6-1  ] =                    (!bj8rlymm54x) & ovco_g1rr8cl[6-1  ];
  assign qkr7a25rdze[6-2:0] = {6-1{j4qv5sod}} & ovco_g1rr8cl[6-2:0];

  assign cvnvrq3lozc = (eaks5rrtzx4 << qkr7a25rdze);

  wire [64-1:0] sr5i7o3ueuv3 = cvnvrq3lozc;
  wire [64-1:0] d8vbgw_alz_l =  osmygk9ar45_;












  wire [64-1:0] hvo606li = {64{1'b1}} >> qkr7a25rdze;
  wire [64-1:0] quqgtuvktbl  =
               (d8vbgw_alz_l & hvo606li) | ({64{svtp9g_orl2[64-1]}} & (~hvo606li));
  wire [31:0] c7w_3utqww = {32{1'b1}} >> qkr7a25rdze;
  wire [31:0] sm06jjtkd6dk8  = (d8vbgw_alz_l[31:0] & c7w_3utqww) | ({32{svtp9g_orl2[31]}} & (~c7w_3utqww));











  wire wxe9so32rgdol = q0brgn6 | rn573wyhxlx2330 | fm3pgkuczco | cod1y7dl_ | e7pwgmzzw54;
  wire [64-1:0] mw6r609jhxx60pytpgc = {{dukom1hk2mc9i6m4 ? yxz3vex1f[64-1:32] : {64-32{~wxe9so32rgdol && yxz3vex1f[31]}}}, yxz3vex1f[31:0]};
  wire [64-1:0] fmcbw4e6ixltp_33vlniu = {{dukom1hk2mc9i6m4 ? afthitl2[64-1:32] : {64-32{~wxe9so32rgdol && afthitl2[31]}}}, afthitl2[31:0]};
  wire [65-1:0] g0aqd08ou7rfnv3ndp =
      {{65-64{(~wxe9so32rgdol) & mw6r609jhxx60pytpgc[64-1]}},mw6r609jhxx60pytpgc[64-1:0]};
  wire [65-1:0] ccbzdmuytukdpcsy26d =
      {{65-64{(~wxe9so32rgdol) & fmcbw4e6ixltp_33vlniu[64-1]}},fmcbw4e6ixltp_33vlniu[64-1:0]};


  wire [65-1:0] ti2vpd9jde = 
      g0aqd08ou7rfnv3ndp;
  wire [65-1:0] xfvd9b_1bqsugi = 
      ccbzdmuytukdpcsy26d;

  wire knqibikmye3;
  wire [65-1:0] atsytx8oasf;
  wire [65-1:0] d_h0rtp1mu2fy;
  wire [65-1:0] wrcjvt7pl1j_;

  wire qqjhj5cz1ue;
  wire gn6aq7h3cy;

  assign qqjhj5cz1ue =
      mf5fcnu2azr | zjk3uzc5cf; 
  assign gn6aq7h3cy =
               (

               (m0mq6jm4ys | obmd5e6) 

             | (egmgssvj3 | nssum1cfr | 
                rn573wyhxlx2330 | fm3pgkuczco |
                b1vnk2xf9 | cod1y7dl_ |
                nsc05do | e7pwgmzzw54 |
                fy1ybps5 | q0brgn6 
               ));

  wire nuhvvo7aaoun4df0 = qqjhj5cz1ue | gn6aq7h3cy; 



  assign atsytx8oasf = {65{nuhvvo7aaoun4df0}} & (ti2vpd9jde);
  assign d_h0rtp1mu2fy = {65{nuhvvo7aaoun4df0}} & (gn6aq7h3cy ? (~xfvd9b_1bqsugi) : xfvd9b_1bqsugi);
  assign knqibikmye3 = nuhvvo7aaoun4df0 & gn6aq7h3cy;

  assign wrcjvt7pl1j_ = atsytx8oasf + d_h0rtp1mu2fy + { {65-1{1'b0}}, knqibikmye3 };








  wire [64-1:0] iept0vlz6lx;
  wire [64-1:0] orrbobw3ayx;

  wire fdy0cez8l = 
               oss8f_hhqe8

             | (g8dm1b58pm6xt | bqmj8280_l); 


  assign iept0vlz6lx = {64{fdy0cez8l}} & yxz3vex1f;
  assign orrbobw3ayx = {64{fdy0cez8l}} & afthitl2;

  wire [64-1:0] zk_1rdw8taxr5 = iept0vlz6lx ^ orrbobw3ayx;

  wire [64-1:0] s63w7cosk_nn  = yxz3vex1f | afthitl2; 
  wire [64-1:0] i3fuqkt9f0 = yxz3vex1f & afthitl2; 





  wire nvna3795  = (|zk_1rdw8taxr5); 
  wire mwi29p2u52  = (bqmj8280_l  & nvna3795);

  wire ucz1nud4yab  = g8dm1b58pm6xt  & (~nvna3795);

  wire tjuogza0f5v  = egmgssvj3  & wrcjvt7pl1j_[64];
  wire xi17iivz6ct = rn573wyhxlx2330 & wrcjvt7pl1j_[64];

  wire wj8lm_uex7d69  = (~wrcjvt7pl1j_[64]);
  wire i8lqt3tmbi2q_2  = nssum1cfr  & wj8lm_uex7d69;
  wire jp5cn3k6s_nnwub = fm3pgkuczco & wj8lm_uex7d69;

  assign ufa33rbvjwk = ucz1nud4yab 
                 | mwi29p2u52 
                 | tjuogza0f5v 
                 | i8lqt3tmbi2q_2  
                 | xi17iivz6ct 
                 | jp5cn3k6s_nnwub; 





  wire [64-1:0] pai2o8ss6k6 = {{(64-32){afthitl2[31]}}, afthitl2[31:0]};
  wire [64-1:0] spnkcpp24vpcjr = pm7lg8nzlruwwz9t29i? pai2o8ss6k6 : afthitl2;





  wire m3lbds76y = (fy1ybps5 | q0brgn6);


  wire hcd2t4f_9lkiz9_lw = m3lbds76y & wrcjvt7pl1j_[64];
  wire [64-1:0] b2110r1fhss = 
               hcd2t4f_9lkiz9_lw ?
               64'b1 : 64'b0;



  wire jkt85o2_yqxb87ehr_y =  ((b1vnk2xf9 | cod1y7dl_) &   wj8lm_uex7d69) 
                      |  ((nsc05do | e7pwgmzzw54) & (~wj8lm_uex7d69));


  wire [64-1:0] qxzve6id9_hb8olf = az6qlcqsx_0[64-1:0];
  wire [64-1:0] sr13svb5rwk75f0 = dukom1hk2mc9i6m4 ? cqqzeukmh[64-1:0] : {{64-32{cqqzeukmh[31]}},cqqzeukmh[31:0]};
  wire [64-1:0] ivcpoenlvs_zrk8  = jkt85o2_yqxb87ehr_y ? qxzve6id9_hb8olf : sr13svb5rwk75f0;  



  wire [64-1:0] gxt8kdblxpj6h_q7 = 
        ({64{nynmmk       }} & s63w7cosk_nn )
      | ({64{tqvnzdez      }} & i3fuqkt9f0)
      | ({64{oss8f_hhqe8      }} & zk_1rdw8taxr5)
      | ({64{uv65k1vtj   }} & wrcjvt7pl1j_[64-1:0])
      | ({64{qi__zhsq1zl9o_w  }} & {{64-32{wrcjvt7pl1j_[31]}},wrcjvt7pl1j_[31:0]})
      | ({64{tdz9d9      }} & d8vbgw_alz_l)
      | ({64{onsk4u1y9_e      }} & sr5i7o3ueuv3)
      | ({64{jxe3dht      }} & quqgtuvktbl)
      | ({64{t1f2vol     }} & {{64-32{d8vbgw_alz_l[31]}},d8vbgw_alz_l[31:0]})
      | ({64{b9bqr_g01     }} & {{64-32{sr5i7o3ueuv3[31]}},sr5i7o3ueuv3[31:0]})
      | ({64{w23f72vq40     }} & {{64-32{sm06jjtkd6dk8[31]}},sm06jjtkd6dk8[31:0]})
      | ({64{x1_dx841    }} & spnkcpp24vpcjr)
      | ({64{m3lbds76y    }} & b2110r1fhss)
      | ({64{b1vnk2xf9 | cod1y7dl_ | nsc05do | e7pwgmzzw54}} & ivcpoenlvs_zrk8)
        ;



  ux607_gnrl_dffl #(64+1) zjut_2sqlm7t_n (t6d11eqb1s3, yoibsjp7ouplcq, tawrhvnsab, gf33atgy, ru_wi);
  ux607_gnrl_dffl #(64+1) cvcju2l8uvyvs2g (em10uopmr98x, iajwu4x_2, o7xczhh6fe, gf33atgy, ru_wi);






  localparam wxbg7z6hn_1rfi1anz2 = ((64*2)+26);

  assign  {
     az6qlcqsx_0
    ,cqqzeukmh
    ,b1vnk2xf9  
    ,nsc05do  
    ,cod1y7dl_ 
    ,e7pwgmzzw54 
    ,mf5fcnu2azr
    ,m0mq6jm4ys
    ,zjk3uzc5cf
    ,obmd5e6
    ,nynmmk
    ,oss8f_hhqe8
    ,tqvnzdez
    ,onsk4u1y9_e
    ,tdz9d9
    ,jxe3dht
    ,b9bqr_g01
    ,t1f2vol
    ,w23f72vq40
    ,fy1ybps5
    ,q0brgn6
    ,x1_dx841
    ,g8dm1b58pm6xt 
    ,bqmj8280_l 
    ,egmgssvj3 
    ,nssum1cfr 
    ,rn573wyhxlx2330
    ,fm3pgkuczco
    }
    = 
        ({wxbg7z6hn_1rfi1anz2{ktu3yhilgxp}} & {
             so01tnkdju7vnwezjvi            
            ,hxad9091n05p_gjjo4            
            ,1'b0                       
            ,1'b0                       
            ,1'b0                       
            ,1'b0                       
            ,odfbwv2n0hmkh9n2v            
            ,vqqbidi8kkzgxc0qls            
            ,tffp7jbfj_acgbf_htp           
            ,mbmpk0lgl7bqaq0m7j           
            ,ngw96h2ls51cor4             
            ,ujg_tx8c5t9t0ddsmq            
            ,cj5vhekber5gw1509m86            
            ,xxf9gqnuyu__15_t1u            
            ,f4uqn8qf5ljfnqy            
            ,k0kxgs4dhk1hf26ky3            
            ,fkbmt37lnc1cbn6h7f5q           
            ,uhs5rs3m1apmo4oj3c7           
            ,hkzo9ego93d08t8igz2           
            ,zouaj0qk3vke9quhfiqz            
            ,u3s5vk_sv9c1gjjto           
            ,pm7lg8nzlruwwz9t29i            
            ,1'b0                       
            ,1'b0                       
            ,1'b0                       
            ,1'b0                       
            ,1'b0                       
            ,1'b0                       
        })
      | ({wxbg7z6hn_1rfi1anz2{fv0c5k6cjre}} & {
             bm6cerfr_1bou52muqp            
            ,tz3kfmltx71a5i0tmaln            
            ,1'b0                       
            ,1'b0                       
            ,1'b0                       
            ,1'b0                       
            ,tz95dh49670qhxle1            
            ,1'b0                       
            ,1'b0                       
            ,1'b0                       
            ,1'b0                       
            ,1'b0                       
            ,1'b0                       
            ,1'b0                       
            ,1'b0                       
            ,1'b0                       
            ,1'b0                       
            ,1'b0                       
            ,1'b0                       
            ,1'b0                       
            ,1'b0                       
            ,1'b0                       
            ,b9asx2rffq8fclg3_q         
            ,m1dubsueroj_o4i9hhxf         
            ,vupdzhdsf5tcdbcy3br3         
            ,rzgzqvqbgh3abztkqck         
            ,n9_mxfs9poavrerrqf3ps        
            ,a8ql4znkrbh_gj7cnnwc2j        
        })
      | ({wxbg7z6hn_1rfi1anz2{yvw7xod98x7}} & {
             tp6hfcjxcyp899mpksjl            
            ,f4ds8dbk9kk_ic_            
            ,hn2h_gkqinydwsdg_i3            
            ,re8hncw6m47hrh6            
            ,tshku7fgpiu2j7ugwjj9           
            ,arc8ztjel_qlz3xfw0ya           
            ,xl9r7gr7wciuv2d00b            
            ,1'b0                       
            ,1'b0                       
            ,1'b0                       
            ,vrqdq7uwxf99gj_7             
            ,jqgtsdtxss_uios07            
            ,htcsb0affil7c6q            
            ,1'b0                       
            ,1'b0                       
            ,1'b0                       
            ,1'b0                       
            ,1'b0                       
            ,1'b0                       
            ,1'b0                       
            ,1'b0                       
            ,oso3fj0gx6pnvjni           
            ,1'b0                       
            ,1'b0                       
            ,1'b0                       
            ,1'b0                       
            ,1'b0                       
            ,1'b0                       
        })
      | ({wxbg7z6hn_1rfi1anz2{hgdur8q6gk2ak91b}} & {
             32'b0                      
            ,32'b0                      
            ,1'b0                       
            ,1'b0                       
            ,1'b0                       
            ,1'b0                       
            ,1'b0                       
            ,1'b0                       
            ,1'b0                       
            ,1'b0                       
            ,1'b0                       
            ,1'b0                       
            ,1'b0                       
            ,r_aei1gc7v37oo9dghv            
            ,1'b0                       
            ,d1_eg4gq3uyxdyycybx            
            ,1'b0                       
            ,1'b0                       
            ,1'b0                       
            ,1'b0                       
            ,1'b0                       
            ,1'b0                       
            ,1'b0                       
            ,1'b0                       
            ,1'b0                       
            ,1'b0                       
            ,1'b0                       
            ,1'b0                       
        })                               
        ;                                

  assign m2s376x2ngd1fz27iofg3yf1 = sr5i7o3ueuv3[64-1:0];
  assign f2mrhq1ax6cmfmtx_l5 = quqgtuvktbl[64-1:0];
  assign uk0gax2bf5vv97rrbosr     = gxt8kdblxpj6h_q7[64-1:0];
  assign ttgsydregi0kgoj_z     = gxt8kdblxpj6h_q7[64-1:0];
  assign todxu2rm67fxk1x8y_tl4 = gxt8kdblxpj6h_q7[64-1:0];
  assign ehhimwdiwsd20nyinnomx = ufa33rbvjwk;

  assign t6d11eqb1s3 = 
                 e__67e1k5hdb4ctnr;
  assign em10uopmr98x = 
                 nc_3q2q5fz4e2;

  assign yoibsjp7ouplcq = 
                 {1'b0,jay_5c6ndpwhj0vqzv};
  assign iajwu4x_2 = 
                 {1'b0,a5y809wbv8w1d0};

  assign kn6tx97_rw9w0v = tawrhvnsab[64-1:0];
  assign l0vxn4vg6wd = o7xczhh6fe[64-1:0];


endmodule                                      

























module n9fwcab7kdqyokfwizktfw(
























































  output  [64-1:0] yqs98coa39vu7,
  output  [64-1:0] cd0szp_7s1jnw,




  input  fj0lzkw_e2tjj, 
  output im2j_m47n4mhs, 

  input  [64-1:0] c5lrjuy9t_f,
  input  [64-1:0] bi9zhg2zyeg,
  input  [64-1:0] iet1_xpdj,
  input  [64-1:0] utdfnsgxzrzt14u,
  input  [48-1:0] ybrrs0__m1aa00,
  input  [4-1:0]        jythgzdjfospqb,
  input                                pkwcaygsgot_59n1,
  input                                vy1aysleh0imu4,
  input                                pbjk7minp0n89j,
  input                                b4uk5z2pu_0s,








  output hgt2urny9_9, 
  input  nrxcyc791r8gksao, 














































































  
  
  
  
  
  
     
  output xl9r7gr7wciuv2d00b,
  output [64-1:0] tp6hfcjxcyp899mpksjl,
  output [64-1:0] f4ds8dbk9kk_ic_,
  input  [64-1:0] ttgsydregi0kgoj_z,


  input  gf33atgy,
  input  ru_wi
  );






  wire       w12tykr0sjk3cb    = ybrrs0__m1aa00 [5:5   ];
  wire       grfzm3doiudavltu   = ybrrs0__m1aa00 [6:6  ];
  wire       v2mydpki2mkh     = ybrrs0__m1aa00 [11:11    ];
  wire [1:0] i2x6qt_wyuanj  = ybrrs0__m1aa00 [28:27];

  wire [1:0] bwnqxkmv3793tn5    = ybrrs0__m1aa00 [8:7   ];
  wire       a02fqysr32bpia6b   = ybrrs0__m1aa00 [9:9  ];
  wire       m2q3ghpncvh    = ybrrs0__m1aa00 [10:10   ];
  wire       uadexzk_kh0g49nb = ybrrs0__m1aa00 [12:12];
  wire       r8x3j28xrzm0eq  = ybrrs0__m1aa00 [13:13 ];
  wire       m5ljd54icrby7u  = ybrrs0__m1aa00 [14:14 ];
  wire       ola68283_q7l   = ybrrs0__m1aa00 [15:15  ];
  wire       icz9kk4dx5uzjcoz  = ybrrs0__m1aa00 [16:16 ];
  wire       qpjjk_tptwhr4qvkz  = ybrrs0__m1aa00 [17:17 ];
  wire       mhi7m13i4tdp  = ybrrs0__m1aa00 [18:18 ];
  wire       qsexm8gncgpsd0 = ybrrs0__m1aa00 [19:19];
  wire       xsjat4ppp7fq3wj = ybrrs0__m1aa00 [20:20];
  wire       db5c7uyis59qjegezc = ybrrs0__m1aa00 [24:24];
  wire       o12r1q7fso07g4lk = ybrrs0__m1aa00 [22:22];
  wire       z5atnp0pqvut7tu3 = ybrrs0__m1aa00 [23:23];
  wire       my6482rcbzjsl0k = ybrrs0__m1aa00 [25:25];
  wire       foo1r_kdsxld_y28ot5 = ybrrs0__m1aa00 [26:26];

    wire       m7pgd062044v      = 1'b0 
                  ; 
    wire       bcz6wdcu6f4c      = 1'b0 
                  ; 
  wire       d8gxc7jp52uv      = w12tykr0sjk3cb  & (i2x6qt_wyuanj == 2'b10); 
  wire       vmlg53ng6oe      = grfzm3doiudavltu & (i2x6qt_wyuanj == 2'b10); 
  wire       av18nzhvobpoka      = w12tykr0sjk3cb  & (i2x6qt_wyuanj == 2'b11); 
  wire       p08f2oxj96slt      = grfzm3doiudavltu & (i2x6qt_wyuanj == 2'b11); 
  wire       jgah5jfw = m7pgd062044v | bcz6wdcu6f4c | d8gxc7jp52uv | vmlg53ng6oe | av18nzhvobpoka | p08f2oxj96slt;
  wire       bp9qt1h52k23 =  av18nzhvobpoka | p08f2oxj96slt;
  wire       t6ehcvrshdj =  m7pgd062044v | bcz6wdcu6f4c | d8gxc7jp52uv | vmlg53ng6oe;
































  wire ip9a_yuu2kn5f  = v2mydpki2mkh | ((w12tykr0sjk3cb | grfzm3doiudavltu) & m2q3ghpncvh); 









  wire [64-1:0] zynejvtsl0wzmfbs8tvbi = 
           jgah5jfw ? utdfnsgxzrzt14u :
          ip9a_yuu2kn5f ? 64'b0 : 
          (db5c7uyis59qjegezc || z5atnp0pqvut7tu3 || o12r1q7fso07g4lk) ? {iet1_xpdj[64-2:0],1'b0} :
          (foo1r_kdsxld_y28ot5 || my6482rcbzjsl0k) ? {iet1_xpdj[64-2:0],1'b0} :
          iet1_xpdj;

  assign xl9r7gr7wciuv2d00b = 1'b1;
  assign tp6hfcjxcyp899mpksjl = 
            (pbjk7minp0n89j & b4uk5z2pu_0s) ? 32'h00000000 :
                         c5lrjuy9t_f; 
  assign f4ds8dbk9kk_ic_ = zynejvtsl0wzmfbs8tvbi ;

  assign yqs98coa39vu7 = tp6hfcjxcyp899mpksjl;
  assign cd0szp_7s1jnw = f4ds8dbk9kk_ic_;









  assign im2j_m47n4mhs =



      nrxcyc791r8gksao  



      ;
















  assign hgt2urny9_9 = 

         fj0lzkw_e2tjj 




          ;
























































































































































































































































































































































































































































endmodule                                      
























module uflzl0cx7tik0xzqybt(
  

  
  
  
  
  input  kg5ogiwmi4x2jcasma, 
  output rbjqmkcrkr7uyq4dauq, 

  input  [64-1:0] w56hh_dniqksvhf,
  input  [64-1:0] q6e0lb86_tx2afeh,
  input  [64-1:0] i5vvhea8kczaa,
  input  [19-1:0] umfak1vbx2r1b,
  input  [4-1:0] i1gdm9hju_gidl,

  output l3kh5v32kt2mkcqz6t,

  input  dnmtm28bd2t,

  
  
  
  output qqrzyv7p9gfzn99, 
  input  ori3109ceulwf9p, 
  output [64-1:0] p3nl1p59c7tkqhr5l8rl,
  output sw6cd2q81orxwjah_hdqq9,   
  

  
  
  
  
     
  output [67-1:0] alse1t6spxo4msbspebwy3y,
  output [67-1:0] x0er7wym12k2zbbkwic3tk,
  output                                g35fohnhd6cn9np610_ ,
  output                                nn3y8_8tdpg0r00cfh22 ,
  input  [67-1:0] tvohxqv2vynsps11_n8jcm1,

     
  output          b9_gjh0acfnkvdnxisky4,
  output [64:0] kjts4h4q5dfneeyrrdrxw,
  input  [64:0] sco_wqinvslwrh,

  output          sj_mdw9rcnoy3tw08nw,
  output [64:0] bx56_yppcspoez2oo86i,
  input  [64:0] tjsikyyrigiuo_,

  input  gf33atgy,
  input  ru_wi
  );

  wire fngy_43kvde0i7yr84 = kg5ogiwmi4x2jcasma & rbjqmkcrkr7uyq4dauq;
  wire db1wnjxow71e6n = qqrzyv7p9gfzn99 & ori3109ceulwf9p;

  
  
  
  
  
  
  assign b9_gjh0acfnkvdnxisky4 = 1'b0;
  assign kjts4h4q5dfneeyrrdrxw = {(64+1){1'b0}};

  assign sj_mdw9rcnoy3tw08nw = 1'b0;
  assign bx56_yppcspoez2oo86i = {(64+1){1'b0}};

  wire fm5qvc    = umfak1vbx2r1b[9:9   ];
  wire ms_4ed   = umfak1vbx2r1b[10:10  ];
  wire i7sstsvqw    = umfak1vbx2r1b[11:11   ];
  wire p4ggl84x_   = umfak1vbx2r1b[12:12  ];

  wire vmw3ij0a96    = umfak1vbx2r1b[15:15    ];
  wire zt4egkm   = umfak1vbx2r1b[16:16   ];
  wire wslud0u    = umfak1vbx2r1b[17:17    ];
  wire ujsqugs   = umfak1vbx2r1b[18:18   ];
      
  
  
  wire cgsm38lhmu = 1'b0;

  wire luu15_fyftf_60kh = cgsm38lhmu;


  
  wire j8b98unuymzt50 = vmw3ij0a96 | zt4egkm | wslud0u  | ujsqugs;
  
  wire qgrzkmut1_u9xo = fm5qvc | ms_4ed | i7sstsvqw  | p4ggl84x_;
  wire knuud64iei = kg5ogiwmi4x2jcasma;
  
  
  wire do24aunj403 = fm5qvc | ms_4ed | vmw3ij0a96 | zt4egkm;
  
  wire a7y71nasc = i7sstsvqw | p4ggl84x_ | wslud0u | ujsqugs;
  
  
  localparam rvvscbdtnunwl5maq8dwovl = 3;

  wire [rvvscbdtnunwl5maq8dwovl-1:0] cwhmtt4bjkyoq2_y;
  wire [rvvscbdtnunwl5maq8dwovl-1:0] xu9sew5enzxvf9nd;
  wire j34mx2nxumsr8qih7e;

  
  localparam pxkzjnxua20t78mk = 3'd0;
  
  localparam cwsvs_tblgh_ip_yu7hw74xe = 3'd1;
  
  localparam vis5wo38luh8olawd3yfg = 3'd2;
  
  localparam dzjqnfvvynffsk4yf6s45w11dxn = 3'd3;
  
  localparam ox_3fqrgcckzzp549az65wysdk = 3'd4;
  
  localparam cvali5t66a_ecwrukwqd4m6xr8 = 3'd5;
  
  localparam rjx0c_5hu03xaw7i_old4c2vq0 = 3'd6;
  
  localparam kcrgmvlnv0aew5yzl_juvo3c = 3'd7;

  wire [rvvscbdtnunwl5maq8dwovl-1:0] fuyfhz6vib9mmow_;
  wire [rvvscbdtnunwl5maq8dwovl-1:0] a2dvifs7ouklsdypatj16;
  wire [rvvscbdtnunwl5maq8dwovl-1:0] nfaffkiutfil4ozf__b;
  wire [rvvscbdtnunwl5maq8dwovl-1:0] hfxd7uehbu5gxfnp4kf;
  wire [rvvscbdtnunwl5maq8dwovl-1:0] yc_p6zm9chckcdpvelu7;
  wire [rvvscbdtnunwl5maq8dwovl-1:0] xuezb11hk022u644tt5d;
  wire [rvvscbdtnunwl5maq8dwovl-1:0] umozcax8c__jn9217ev_kr6;
  wire [rvvscbdtnunwl5maq8dwovl-1:0] w6czcbj6628j7_dt9;

  wire emzbemdseyus6f56bkir7;
  wire vayxkylokyi6tov7_8vpi0jl47_y4kf;
  wire sufue9iopakxbuyxa_u;
  wire mgv19caed0r5x4i1r8tvm6j1;
  wire clm755bo643p6w08dbql_ean;
  wire t221bf_qpb_zxne6bm4s59bidk7;
  wire ul1h3698licmbmnzglsrzaogq4qa;
  wire yak839qok7m09acgj84zgsuz6zb;

  wire zlw2z06rh9jw8sq;
  wire nic33i142fgdyocr6vrotyt = kg5ogiwmi4x2jcasma & (~luu15_fyftf_60kh) & (~zlw2z06rh9jw8sq);

  
  wire   tctggwwx9ewc2bnbum7rgp          = (xu9sew5enzxvf9nd == pxkzjnxua20t78mk        );
  wire   at44jvmwzm87ug8_qz3intfeb055kf  = (xu9sew5enzxvf9nd == cwsvs_tblgh_ip_yu7hw74xe);
  wire   ol1caffg7ftaluj4jy0b         = (xu9sew5enzxvf9nd == vis5wo38luh8olawd3yfg       );
  wire   mtfz_0a_x9uvv8pxxcgu5o7hszz    = (xu9sew5enzxvf9nd == dzjqnfvvynffsk4yf6s45w11dxn  );
  wire   z_1u5zn8t754l0hxm5qcqea_d1jd    = (xu9sew5enzxvf9nd == ox_3fqrgcckzzp549az65wysdk  );
  wire   yf1hpaj7zyyyzd1dicudtlr0oar    = (xu9sew5enzxvf9nd == cvali5t66a_ecwrukwqd4m6xr8  );
  wire   u_90mukpto0u7au4dgn0xciq0xg77   = (xu9sew5enzxvf9nd == rjx0c_5hu03xaw7i_old4c2vq0 );
  wire   s91yobxezoiswejay4ga8v63y      = (xu9sew5enzxvf9nd == kcrgmvlnv0aew5yzl_juvo3c    );
  
    
  
          
  assign emzbemdseyus6f56bkir7 = tctggwwx9ewc2bnbum7rgp & nic33i142fgdyocr6vrotyt & (~dnmtm28bd2t);
  assign fuyfhz6vib9mmow_      = cwsvs_tblgh_ip_yu7hw74xe;

      
          
  assign vayxkylokyi6tov7_8vpi0jl47_y4kf = (at44jvmwzm87ug8_qz3intfeb055kf & (dnmtm28bd2t | 1'b1));
  assign a2dvifs7ouklsdypatj16      = dnmtm28bd2t ? pxkzjnxua20t78mk : vis5wo38luh8olawd3yfg;

      
  wire tvmuha1_tqa;
  wire aejagosb1fvtgozqa7l7rgsi; 
  assign sufue9iopakxbuyxa_u =  ol1caffg7ftaluj4jy0b & ((
          
                           aejagosb1fvtgozqa7l7rgsi 
              
                         & (knuud64iei ? 1'b1
              
                                            : db1wnjxow71e6n))
            | dnmtm28bd2t);
  assign nfaffkiutfil4ozf__b      = 
                (
                         dnmtm28bd2t ? pxkzjnxua20t78mk :
              
                                       dzjqnfvvynffsk4yf6s45w11dxn
                );

      
          
          
  wire y07pr2allup91cvwe9o; 
  wire nnex5qu4d62mmyuuef; 
  wire ljbp87zj73pp;
  
  assign mgv19caed0r5x4i1r8tvm6j1 = (mtfz_0a_x9uvv8pxxcgu5o7hszz & ( dnmtm28bd2t | 1'b1)); 
  assign hfxd7uehbu5gxfnp4kf      = dnmtm28bd2t                                     ? pxkzjnxua20t78mk :
              
                                    (do24aunj403 & nnex5qu4d62mmyuuef)                 ? ox_3fqrgcckzzp549az65wysdk :
              
                                    (do24aunj403 & ~nnex5qu4d62mmyuuef & ljbp87zj73pp)   ? kcrgmvlnv0aew5yzl_juvo3c :
              
                                    (a7y71nasc & y07pr2allup91cvwe9o)                  ? cvali5t66a_ecwrukwqd4m6xr8 :
              
                                    (a7y71nasc & ~y07pr2allup91cvwe9o)                 ? rjx0c_5hu03xaw7i_old4c2vq0 :
              
                                                                                      pxkzjnxua20t78mk;

      
          
  assign clm755bo643p6w08dbql_ean = (z_1u5zn8t754l0hxm5qcqea_d1jd & (dnmtm28bd2t | 1'b1));
  assign yc_p6zm9chckcdpvelu7      = dnmtm28bd2t ? pxkzjnxua20t78mk :
                                    ljbp87zj73pp  ? kcrgmvlnv0aew5yzl_juvo3c :
                                                  pxkzjnxua20t78mk;

                
      
              
  assign t221bf_qpb_zxne6bm4s59bidk7 = (yf1hpaj7zyyyzd1dicudtlr0oar & (dnmtm28bd2t | 1'b1));
  assign xuezb11hk022u644tt5d      = dnmtm28bd2t ?   pxkzjnxua20t78mk : 
                                                    rjx0c_5hu03xaw7i_old4c2vq0;
  
      
         
  assign ul1h3698licmbmnzglsrzaogq4qa = (u_90mukpto0u7au4dgn0xciq0xg77 & (dnmtm28bd2t | 1'b1));
  assign umozcax8c__jn9217ev_kr6 = dnmtm28bd2t         ? pxkzjnxua20t78mk :
                                tvmuha1_tqa          ? kcrgmvlnv0aew5yzl_juvo3c :
                                                      pxkzjnxua20t78mk;

      
          
  assign yak839qok7m09acgj84zgsuz6zb = (s91yobxezoiswejay4ga8v63y & (dnmtm28bd2t | 1'b1));
  assign w6czcbj6628j7_dt9      = pxkzjnxua20t78mk;


  
  assign j34mx2nxumsr8qih7e = emzbemdseyus6f56bkir7 
                          | vayxkylokyi6tov7_8vpi0jl47_y4kf  
                          | sufue9iopakxbuyxa_u  
                          | mgv19caed0r5x4i1r8tvm6j1  
                          | clm755bo643p6w08dbql_ean  
                          | t221bf_qpb_zxne6bm4s59bidk7  
                          | ul1h3698licmbmnzglsrzaogq4qa
                          | yak839qok7m09acgj84zgsuz6zb  
                          ;

  
  assign cwhmtt4bjkyoq2_y = 
              ({rvvscbdtnunwl5maq8dwovl{emzbemdseyus6f56bkir7        }} & fuyfhz6vib9mmow_        )
            | ({rvvscbdtnunwl5maq8dwovl{vayxkylokyi6tov7_8vpi0jl47_y4kf}} & a2dvifs7ouklsdypatj16)            
            | ({rvvscbdtnunwl5maq8dwovl{sufue9iopakxbuyxa_u       }} & nfaffkiutfil4ozf__b       )
            | ({rvvscbdtnunwl5maq8dwovl{mgv19caed0r5x4i1r8tvm6j1  }} & hfxd7uehbu5gxfnp4kf  )
            | ({rvvscbdtnunwl5maq8dwovl{clm755bo643p6w08dbql_ean  }} & yc_p6zm9chckcdpvelu7  )
            | ({rvvscbdtnunwl5maq8dwovl{t221bf_qpb_zxne6bm4s59bidk7  }} & xuezb11hk022u644tt5d  )
            | ({rvvscbdtnunwl5maq8dwovl{ul1h3698licmbmnzglsrzaogq4qa }} & umozcax8c__jn9217ev_kr6 )            
            | ({rvvscbdtnunwl5maq8dwovl{yak839qok7m09acgj84zgsuz6zb    }} & w6czcbj6628j7_dt9    )            
              ;

  ux607_gnrl_dfflr #(rvvscbdtnunwl5maq8dwovl) ummoxvcagl4gsz63jh (j34mx2nxumsr8qih7e, cwhmtt4bjkyoq2_y, xu9sew5enzxvf9nd, gf33atgy, ru_wi);
  
  wire rm11i0fhvrvpa2j4j8fhanxxybj6 = j34mx2nxumsr8qih7e & (cwhmtt4bjkyoq2_y == cwsvs_tblgh_ip_yu7hw74xe);
  wire gilndp855iiulx68zkl50 = j34mx2nxumsr8qih7e & (cwhmtt4bjkyoq2_y == vis5wo38luh8olawd3yfg);
  localparam jt3ho7cizyka  = 7;
  localparam mjj76ct8o1p  = 7'd0 ;
  localparam cj0jb1qkpn  = 7'd1 ;
  localparam hwwdbfi52t4tum = 7'd32;
  localparam pm42q8y0fkk5_sq = 7'd64;
  localparam m6d1zd37y4qv2qt_e5 = 7'd16;  
  localparam p0u0coqmf6fkp75 = 7'd32;  
  localparam tj72am0aq9mmw_seuh = 7'd64;  
  localparam xqgqwa5rixv = 7;
  localparam uic4wt9w_k = 6;
  localparam nz92trl63p09bhd = 7'd18;
  localparam dzttnj6s8jqu7a = 7'd34;


  wire[jt3ho7cizyka-1:0] l2m2s106w95k;
  wire on52gxi2i1_8p5_ = rm11i0fhvrvpa2j4j8fhanxxybj6; 
  wire mdp_a_1uzeiv = gilndp855iiulx68zkl50;
  wire z3q0v1s1_muk73 = ol1caffg7ftaluj4jy0b & (~aejagosb1fvtgozqa7l7rgsi); 
  wire g59yhxfbkwd12 = z3q0v1s1_muk73 | mdp_a_1uzeiv | on52gxi2i1_8p5_; 
    
  wire[jt3ho7cizyka-1:0] ecpjvly4p6z78t = on52gxi2i1_8p5_ ? mjj76ct8o1p : 
                                      mdp_a_1uzeiv ? cj0jb1qkpn : 
                                                     (l2m2s106w95k + {{jt3ho7cizyka-1{1'b0}},1'b1});
  ux607_gnrl_dfflr #(jt3ho7cizyka) mbui732ruwohkr (g59yhxfbkwd12, ecpjvly4p6z78t, l2m2s106w95k, gf33atgy, ru_wi);
  

  wire imnkcvuxli11  = l2m2s106w95k == mjj76ct8o1p;
  
  
  wire uxstct0v10h4tde = (l2m2s106w95k == m6d1zd37y4qv2qt_e5);
  
  wire mg126ouq2dqjk = (l2m2s106w95k == dzttnj6s8jqu7a);

  wire[xqgqwa5rixv-1:0] toomwmpbxsmlbhqtx0oi8y4pw;
  assign aejagosb1fvtgozqa7l7rgsi = knuud64iei & (l2m2s106w95k == toomwmpbxsmlbhqtx0oi8y4pw );








 
  wire g88mwavu3olf = (ms_4ed | p4ggl84x_ | zt4egkm | ujsqugs) ? 1'b0 : 
                      (vmw3ij0a96 | wslud0u)                     ? w56hh_dniqksvhf[31]  :
                                                              w56hh_dniqksvhf[64-1];
  wire ybtjcyiwk275d = (ms_4ed | p4ggl84x_ | zt4egkm | ujsqugs) ? 1'b0 : 
                      (vmw3ij0a96 | wslud0u)                     ? q6e0lb86_tx2afeh[31]  :
                                                              q6e0lb86_tx2afeh[64-1];
  
  
  
  wire hwh65zabyknriqont = g88mwavu3olf & (i7sstsvqw | wslud0u);
  wire uhsepkgpelpn0p = at44jvmwzm87ug8_qz3intfeb055kf;
  ux607_gnrl_dfflr #(1) v56i02t7d4czdn (uhsepkgpelpn0p, hwh65zabyknriqont, tvmuha1_tqa, gf33atgy, ru_wi);


  wire g8fx0qh5o49qm6d6 = (g88mwavu3olf ^ ybtjcyiwk275d) & (fm5qvc | vmw3ij0a96);
  wire aza6vs1oui8scst8 = at44jvmwzm87ug8_qz3intfeb055kf;
  ux607_gnrl_dfflr #(1) rodyya_ynntagpf2 (aza6vs1oui8scst8, g8fx0qh5o49qm6d6, ljbp87zj73pp, gf33atgy, ru_wi);



  
  wire [67-1:0] q70hd825o9qzbjbjck_nkdbjw;

  wire pu0twvle6ws8u7d = ( (vmw3ij0a96 | wslud0u) & w56hh_dniqksvhf[31] ) | ( (fm5qvc | i7sstsvqw) & w56hh_dniqksvhf[64-1] );
  wire o1iwv1o5h4362hx7ih4wwt = ~pu0twvle6ws8u7d;
  
  wire [64-1:0] prooawqnpajt1laptu = pu0twvle6ws8u7d? ~w56hh_dniqksvhf : w56hh_dniqksvhf;
  
  wire b95_l8ftvsr7lpu6b2d = ( (vmw3ij0a96 | wslud0u) & q6e0lb86_tx2afeh[31] ) | ( (fm5qvc | i7sstsvqw) & q6e0lb86_tx2afeh[64-1] );
  
  wire [64-1:0] aypc6it61ljlyo7fl8 = q70hd825o9qzbjbjck_nkdbjw[64-1:0];
  wire [64-1:0] hz0h3cdzl_s9ramg8_z = b95_l8ftvsr7lpu6b2d? aypc6it61ljlyo7fl8 :  q6e0lb86_tx2afeh;

  wire [64-1:0] purxqwoq9lnp7ectr = (vmw3ij0a96 | zt4egkm | wslud0u | ujsqugs) ? {prooawqnpajt1laptu[31:0], 32'b0} : prooawqnpajt1laptu;
  wire [64-1:0] tplwh7047vgl7fiatx5  = (vmw3ij0a96 | zt4egkm | wslud0u | ujsqugs) ? {hz0h3cdzl_s9ramg8_z[31:0], 32'b0} : hz0h3cdzl_s9ramg8_z;
  
  wire [64-1:0] oxmqqogsjqsx78fh;
  wire yim0q0jmj06649ub = tctggwwx9ewc2bnbum7rgp & knuud64iei;
  ux607_gnrl_dfflr #(64) yfy12oxq2liksuz9y_t (yim0q0jmj06649ub, tplwh7047vgl7fiatx5, oxmqqogsjqsx78fh, gf33atgy, ru_wi);

  
  wire [uic4wt9w_k-1:0] pun0eqbgync25oxt8;
  wire [uic4wt9w_k-1:0] lk6k6mq63szqj9buqf;
  wire asdj74mldfl30j_5j37wb9br = at44jvmwzm87ug8_qz3intfeb055kf & knuud64iei;
  ux607_gnrl_dfflr #(uic4wt9w_k) t90qhin2_cspdzrs87desq0 (asdj74mldfl30j_5j37wb9br, pun0eqbgync25oxt8, lk6k6mq63szqj9buqf, gf33atgy, ru_wi);

  crj9jaav6wgkqbu1 #(.onr7l(64),.hw3qvr(6)) b6xrt0rr88sbo0  (.bjh(oxmqqogsjqsx78fh), .ht70(pun0eqbgync25oxt8));

  assign toomwmpbxsmlbhqtx0oi8y4pw = lk6k6mq63szqj9buqf[uic4wt9w_k-1:1]+1'b1;

  wire [64-1:0] qimb_d7m_730jbt5j48_k_; 
  wire [64-1:0] kfw9_6qenp0if86lrw1vdq4v0ow = oxmqqogsjqsx78fh << pun0eqbgync25oxt8;
  wire s6b5h8rrun5fg2aurot43nd3f = at44jvmwzm87ug8_qz3intfeb055kf;
  ux607_gnrl_dfflr #(64) eluy9pwcfd6awd4g0g3v59nb (s6b5h8rrun5fg2aurot43nd3f, kfw9_6qenp0if86lrw1vdq4v0ow, qimb_d7m_730jbt5j48_k_, gf33atgy, ru_wi);

  wire [68-1:0] mjx3_lt0fd_ = {4'b0,purxqwoq9lnp7ectr};
  wire [68-1:0] uw_hf_3q  = {3'b0,qimb_d7m_730jbt5j48_k_,1'b0};

  wire [68-1:0] jgc8ze0wjsbov451fa88rr =  uw_hf_3q;
  wire [68-1:0] mv7gmrm_p6q993kpqk = ~uw_hf_3q;

  wire [68-1:0] rkcxlhptlv8k8zsuxv4;
  wire [68-1:0] bk4ft_fijbgsyx_;
  wire [68-1:0] n77tq9d9umlm_q0v6yb;
  wire [68-1:0] s2cksdp0bmh__nk3;
  wire [68-1:0] xxdi9_qz2jew54h;

  
  wire l_sb2nwq4d1xsvxf38q = mdp_a_1uzeiv & knuud64iei;
  wire rdku4m3qpoja9iicn6wh = z3q0v1s1_muk73 & knuud64iei; 

  wire vhogvq2t73k0zvs6i = l_sb2nwq4d1xsvxf38q | rdku4m3qpoja9iicn6wh | sufue9iopakxbuyxa_u | t221bf_qpb_zxne6bm4s59bidk7;
  

  wire [67-1:0] u_g9a1qe8dho70ggv3ae624yp;
  wire [67-1:0] hil28bjka808mauzn50b7l1xq; 
  wire [67-1:0] topbsq9vgz4_chsttkg7n; 
  wire [64-1:0] rdf2np3w;
  wire [64-1:0] vttcbkxuic7ybtrh;

  wire [68-1:0] jior3mbjv6sgdl;
  wire [68-1:0] dvooronxj88s4wy =  ({68{imnkcvuxli11               }} & mjx3_lt0fd_                     )                      
                                            | ({68{ol1caffg7ftaluj4jy0b      }} & rkcxlhptlv8k8zsuxv4               )
                                            | ({68{mtfz_0a_x9uvv8pxxcgu5o7hszz }} & {1'b0, hil28bjka808mauzn50b7l1xq})
                                            | ({68{yf1hpaj7zyyyzd1dicudtlr0oar }} & {1'b0, topbsq9vgz4_chsttkg7n})
                                            | ({68{u_90mukpto0u7au4dgn0xciq0xg77}} & {4'b0, vttcbkxuic7ybtrh         })
                                            ;
                                                                                                        
  wire qeiwllctq_d1db73j = vhogvq2t73k0zvs6i | mtfz_0a_x9uvv8pxxcgu5o7hszz | u_90mukpto0u7au4dgn0xciq0xg77;
  ux607_gnrl_dffl #(68) goy993rzja07b20io_fp(qeiwllctq_d1db73j, dvooronxj88s4wy, jior3mbjv6sgdl, gf33atgy, ru_wi);

  wire [68-1:0] l8elw6lkpkwm2lgm5s = o1iwv1o5h4362hx7ih4wwt ? {68{1'b0}} : 
                                             j8b98unuymzt50           ? {35'b0,1'b1,32'b0}    :
                                                                   {{(68-1){1'b0}}, 1'b1};

  wire [68-1:0] har15kbia_8670;
  wire [68-1:0] gkrmlupuwwhley9gs = mtfz_0a_x9uvv8pxxcgu5o7hszz ?  {68{1'b0}}:
                                             imnkcvuxli11 ?                l8elw6lkpkwm2lgm5s : 
                                                                        bk4ft_fijbgsyx_;

  wire o1o6ho80flf8qk1v73n = vhogvq2t73k0zvs6i | mtfz_0a_x9uvv8pxxcgu5o7hszz;
  ux607_gnrl_dffl #(68) trm6lzh224boye01116eb(o1o6ho80flf8qk1v73n, gkrmlupuwwhley9gs, har15kbia_8670, gf33atgy, ru_wi);

  wire [68-1:0] rrdj9beol47k9qwcte;
  wire [68-1:0] nvfyzrhxggm8d4x57 = imnkcvuxli11 ? {68{1'b0}} : n77tq9d9umlm_q0v6yb; 
  ux607_gnrl_dffl #(68) nnfpkouay1l48khdt1qx(vhogvq2t73k0zvs6i, nvfyzrhxggm8d4x57, rrdj9beol47k9qwcte, gf33atgy, ru_wi);

  wire [68-1:0] l70r12wporrm20;
  wire [64-1:0] y94wq56bk3vnomt_ = l70r12wporrm20[64+2:3] >> (64-1-lk6k6mq63szqj9buqf);
  wire uyxgfxu16eskur3nt = vhogvq2t73k0zvs6i | mtfz_0a_x9uvv8pxxcgu5o7hszz | z_1u5zn8t754l0hxm5qcqea_d1jd ;
  wire [68-1:0] lkf0ta9fwl1rthw0nla0 =  ({68{imnkcvuxli11              }} & {68{1'b0}        })
                                            | ({68{ol1caffg7ftaluj4jy0b     }} & {s2cksdp0bmh__nk3             })
                                            | ({68{mtfz_0a_x9uvv8pxxcgu5o7hszz}} & {4'b0, y94wq56bk3vnomt_         })
                                            | ({68{z_1u5zn8t754l0hxm5qcqea_d1jd}} & {1'b0, u_g9a1qe8dho70ggv3ae624yp})
                                            ;

  ux607_gnrl_dffl #(68) svvmfr0z3pehqsxi(uyxgfxu16eskur3nt, lkf0ta9fwl1rthw0nla0, l70r12wporrm20, gf33atgy, ru_wi);


  wire [68-1:0] hxn0kheaar53byy;
  wire [68-1:0] va6kvorr04ff34tab = imnkcvuxli11 ? {68{1'b0}} : xxdi9_qz2jew54h;
  ux607_gnrl_dffl #(68) l1wsyj6f4anwfmwz6(vhogvq2t73k0zvs6i, va6kvorr04ff34tab, hxn0kheaar53byy, gf33atgy, ru_wi);

  wire k2xz1iocfj4qk7btop = ~lk6k6mq63szqj9buqf[0] & aejagosb1fvtgozqa7l7rgsi;


  jvwuov7by1m8upbjlyy6 egutfe1kb9mrcsmlryeiun(
    .rydw                (jior3mbjv6sgdl),
    .d4y                (har15kbia_8670),
    .iev4j_o4            (jgc8ze0wjsbov451fa88rr),
    .hfl_1crp            (mv7gmrm_p6q993kpqk),
    .h891r               (rrdj9beol47k9qwcte),
    .m48h                (l70r12wporrm20),
    .r04h               (hxn0kheaar53byy),
    .k2xz1iocfj4qk7btop    (k2xz1iocfj4qk7btop),

    .kktrbu07             (rkcxlhptlv8k8zsuxv4),
    .kf9hl8c_             (bk4ft_fijbgsyx_),
    .spfqyly64           (n77tq9d9umlm_q0v6yb),
    .dqm4y5o             (s2cksdp0bmh__nk3),
    .tzwq6o86            (xxdi9_qz2jew54h)
    );


       
       
       
           

  wire [64-1:0] qhjeo561rub87 = mtfz_0a_x9uvv8pxxcgu5o7hszz ? y94wq56bk3vnomt_ : tvohxqv2vynsps11_n8jcm1[64-1:0];


  wire [67-1:0] b13rowm96j8tw7ylhiu1u = 
                                            (vmw3ij0a96 | wslud0u) ? {{67-64{1'b0}},32'b0, ~q6e0lb86_tx2afeh[31:0]} :
                                            {{67-64{1'b0}}, ~q6e0lb86_tx2afeh};

  wire [67-1:0] hxgjhh23aui05xqtg5f9bxz7h = {{(67-1){1'b0}},1'b1};

  wire dec916j3r2kt10vqxhap5u = 1'b1;
  wire vv0_j637dpg5b6n4ckkem = 1'b0;
 
  assign q70hd825o9qzbjbjck_nkdbjw = tvohxqv2vynsps11_n8jcm1; 

  
  assign hil28bjka808mauzn50b7l1xq = tvohxqv2vynsps11_n8jcm1;
  wire [67-1:0] jhkcorqz91nr_rgl65lrkk = jior3mbjv6sgdl[67-1:0];
  wire [67-1:0] mfpizpziwuw6sxkonddalx = har15kbia_8670[67-1:0];
  wire p0cthoh7mrvh6ea4hqf3j = 1'b1; 
  wire bng35hngtrw10ln9w4fek5rrdh = 1'b0; 
  
  assign y07pr2allup91cvwe9o = hil28bjka808mauzn50b7l1xq[67-1] & a7y71nasc;
  assign nnex5qu4d62mmyuuef = hil28bjka808mauzn50b7l1xq[67-1] & do24aunj403;
  

  assign u_g9a1qe8dho70ggv3ae624yp = tvohxqv2vynsps11_n8jcm1;
  wire [67-1:0] w33jdq7vfismzww2ajvuy6n = {{67-64{1'b0}}, l70r12wporrm20[64-1:0]};
  wire [67-1:0] xchyn0dpmgd_hjajz528eg = {{(67-1){1'b0}}, 1'b1};
  wire n598ep7r9jm04bk34zmlc2dyua = 1'b0;
  wire jchfur14o10iq8hk53nzt = 1'b1;

  assign topbsq9vgz4_chsttkg7n = tvohxqv2vynsps11_n8jcm1;
  wire [67-1:0] xw6vae9ktdr7ai1f1x06r610u4 = jior3mbjv6sgdl[67-1:0];
  wire [67-1:0] dhg2fu358rxsvd8az8ydnz5 = uw_hf_3q[67-1:0];
  wire te1ug32hvsiuidvsmeb0cxuy = 1'b1;
  wire noko_faipjic3du4_u6pwlz = 1'b0;


  wire [64-1:0] cpqevr1sbluf2vtuagep_u8 = tvohxqv2vynsps11_n8jcm1[64-1:0];
  wire [67-1:0] e8ornbgozwvrhsc484js77xw = ljbp87zj73pp ?  {{67-64{1'b1}},~l70r12wporrm20[64-1:0]} : {{67-64{1'b1}}, ~jior3mbjv6sgdl[64-1:0]};
  wire [67-1:0] j6v8x95y_q4ghbmmin5397f = {{(67-1){1'b0}},1'b1};
  wire dr0ydrozi_owdg77zer = 1'b1;
  wire izorepwjzxcb317s53sjme1 = 1'b0;
 


  wire [64-1:0] k6b39gmh_vqvzhin = (wslud0u | ujsqugs) ? {{(64/2){1'b0}}, jior3mbjv6sgdl[64:64/2+1]} :  jior3mbjv6sgdl[64:1];
  assign vttcbkxuic7ybtrh = k6b39gmh_vqvzhin >> lk6k6mq63szqj9buqf;

  wire [64-1:0] pjse89toq0f7cyuut = cpqevr1sbluf2vtuagep_u8;


  assign rdf2np3w = s91yobxezoiswejay4ga8v63y    ? pjse89toq0f7cyuut : 
                    u_90mukpto0u7au4dgn0xciq0xg77 ? vttcbkxuic7ybtrh :
                                               topbsq9vgz4_chsttkg7n[64-1:0];

  wire[64-1:0] bcpc42f7 = (fm5qvc | ms_4ed | vmw3ij0a96 | zt4egkm ) ? qhjeo561rub87[64-1:0] : rdf2np3w[64-1:0];
  

  



  wire pbnf388q25tg_q8 = ~(|q6e0lb86_tx2afeh);
  wire v17qh3l8zn8sg_ = j8b98unuymzt50 & (~(|q6e0lb86_tx2afeh[31:0]));
  wire bq1jtw_wg7ht = pbnf388q25tg_q8 | v17qh3l8zn8sg_;

  wire hu_ub8tznh7e47cd6 = (fm5qvc | i7sstsvqw ) & (&q6e0lb86_tx2afeh)  
                        
                     & w56hh_dniqksvhf[64-1] & (~(|w56hh_dniqksvhf[64-2:0]));
  wire c_vwhek_9xyf = (vmw3ij0a96 | wslud0u) & (&q6e0lb86_tx2afeh[31:0]) & w56hh_dniqksvhf[31] & (~(|w56hh_dniqksvhf[30:0]));
  wire vtoxra6 = hu_ub8tznh7e47cd6 | c_vwhek_9xyf;

  wire rz1_ifrea7y8b_a6f6 = vmw3ij0a96 & (w56hh_dniqksvhf == 64'd9) & (q6e0lb86_tx2afeh == 64'd7); 

  wire[64-1:0] tsfrfbnur6pyx7wmb = ~64'b0;
  
  wire[64-1:0] s4n7oocjmwj88wbbkr = (wslud0u | ujsqugs) ? {{64/2{w56hh_dniqksvhf[64/2-1]}}, w56hh_dniqksvhf[64/2-1:0]} :  w56hh_dniqksvhf[64-1:0];
  
  wire[64-1:0] nb80y93tuo2ieimbw = (fm5qvc | ms_4ed | vmw3ij0a96 | zt4egkm) ? tsfrfbnur6pyx7wmb : s4n7oocjmwj88wbbkr;

  wire[64-1:0] hi9r1vhsx607_tnzh  = (vmw3ij0a96) ? {{64/2+1{1'b1}},{64/2-1{1'b0}}} : {1'b1,{64-1{1'b0}}};
  wire[64-1:0] ntimmdhpytkts505  = 64'b0;
  
  wire[64-1:0] hh7lzf537ly6ek3 = (fm5qvc | vmw3ij0a96) ? hi9r1vhsx607_tnzh : ntimmdhpytkts505;
  wire[64-1:0] vt3rj774l75g34d41de0djyf = {{(64-1){1'b0}},1'b1};


  wire nl6zemz9mxoe59gusvnn = knuud64iei & (bq1jtw_wg7ht | vtoxra6 | rz1_ifrea7y8b_a6f6);
  
  wire[64-1:0] lbeu_v4zoishx6w = bq1jtw_wg7ht ? nb80y93tuo2ieimbw 
                                       : vtoxra6  ? hh7lzf537ly6ek3
                                       :            vt3rj774l75g34d41de0djyf
                                       ;







  assign zlw2z06rh9jw8sq = nl6zemz9mxoe59gusvnn;
  wire[64-1:0] jh7_lyxa4z44z_sv = lbeu_v4zoishx6w;

  
  

    
    
    
    
  wire mtvxxowxa9 = (luu15_fyftf_60kh | zlw2z06rh9jw8sq) ? 1'b1 : 
                       (
                           (ol1caffg7ftaluj4jy0b & aejagosb1fvtgozqa7l7rgsi & (~knuud64iei))
                         | (mtfz_0a_x9uvv8pxxcgu5o7hszz & (do24aunj403) & (~nnex5qu4d62mmyuuef) & (~ljbp87zj73pp) )
                         | (z_1u5zn8t754l0hxm5qcqea_d1jd & (~ljbp87zj73pp))
                         | (u_90mukpto0u7au4dgn0xciq0xg77 & (~tvmuha1_tqa))
                         | (s91yobxezoiswejay4ga8v63y)
                       );
                       
  assign qqrzyv7p9gfzn99 = mtvxxowxa9 & kg5ogiwmi4x2jcasma;
  assign rbjqmkcrkr7uyq4dauq = mtvxxowxa9 & ori3109ceulwf9p;
  wire gsdm0k7q0pb_f = zlw2z06rh9jw8sq;
  wire xpzybyn4n22  = (~luu15_fyftf_60kh) & (~zlw2z06rh9jw8sq) & qgrzkmut1_u9xo;
  wire i5qwugguk8muyt7 = (~luu15_fyftf_60kh) & (~zlw2z06rh9jw8sq) & j8b98unuymzt50;
  assign p3nl1p59c7tkqhr5l8rl = 
               ({64{gsdm0k7q0pb_f}} & jh7_lyxa4z44z_sv)
             | ({64{xpzybyn4n22}} & bcpc42f7)
             | ({64{i5qwugguk8muyt7}} & {{32{bcpc42f7[31]}},bcpc42f7[31:0]})
             ;

  
  assign sw6cd2q81orxwjah_hdqq9 = 1'b0;

     
  wire ckphz278a4bkhg = knuud64iei & tctggwwx9ewc2bnbum7rgp;
  wire sw736m_p2mupr1mfk = knuud64iei & mtfz_0a_x9uvv8pxxcgu5o7hszz;
  wire m10asfr9f1sq = knuud64iei & z_1u5zn8t754l0hxm5qcqea_d1jd;
  wire rsp_p6j830ce7p_8 = knuud64iei & yf1hpaj7zyyyzd1dicudtlr0oar;
  wire yxzdrswl5m2n1c = knuud64iei & s91yobxezoiswejay4ga8v63y  ;

  assign alse1t6spxo4msbspebwy3y = 
             ({67{ckphz278a4bkhg}} & b13rowm96j8tw7ylhiu1u)
           | ({67{sw736m_p2mupr1mfk}} & jhkcorqz91nr_rgl65lrkk)
           | ({67{m10asfr9f1sq}} & w33jdq7vfismzww2ajvuy6n)
           | ({67{rsp_p6j830ce7p_8}} & xw6vae9ktdr7ai1f1x06r610u4)
           | ({67{yxzdrswl5m2n1c}} & e8ornbgozwvrhsc484js77xw  );

  assign x0er7wym12k2zbbkwic3tk =
             ({67{ckphz278a4bkhg}} & hxgjhh23aui05xqtg5f9bxz7h)
           | ({67{sw736m_p2mupr1mfk}} & mfpizpziwuw6sxkonddalx)
           | ({67{m10asfr9f1sq}} & xchyn0dpmgd_hjajz528eg)
           | ({67{rsp_p6j830ce7p_8}} & dhg2fu358rxsvd8az8ydnz5) 
           | ({67{yxzdrswl5m2n1c}} & j6v8x95y_q4ghbmmin5397f  );

  assign g35fohnhd6cn9np610_  = 
             (ckphz278a4bkhg & dec916j3r2kt10vqxhap5u)
           | (sw736m_p2mupr1mfk & p0cthoh7mrvh6ea4hqf3j)
           | (m10asfr9f1sq & n598ep7r9jm04bk34zmlc2dyua)
           | (rsp_p6j830ce7p_8 & te1ug32hvsiuidvsmeb0cxuy) 
           | (yxzdrswl5m2n1c & dr0ydrozi_owdg77zer  );

  assign nn3y8_8tdpg0r00cfh22  = 
             (ckphz278a4bkhg & vv0_j637dpg5b6n4ckkem)
           | (sw736m_p2mupr1mfk & bng35hngtrw10ln9w4fek5rrdh)
           | (m10asfr9f1sq & jchfur14o10iq8hk53nzt)
           | (rsp_p6j830ce7p_8 & noko_faipjic3du4_u6pwlz) 
           | (yxzdrswl5m2n1c & izorepwjzxcb317s53sjme1  );


  
  assign l3kh5v32kt2mkcqz6t = 1'b0;





endmodule                                      























module q8buuqlskug7714mfcon71(





  input  c6cxk8927p4f, 
  output m2_8aknpfse, 

  input  [64-1:0] dn0217a1asgpu,
  input  [64-1:0] jzpnr2l6ruhz,
  input  [64-1:0] nlpn_dhtplj1_,
  input  [64-1:0] biu3jln6jgq,
  input  [47-1:0] zojgfxfr_e4,




  output r9hdxtws4mibgldl, 
  input  olti9ndjvk_sohpa, 

  output [64-1:0] n67h_nt2we0os531a,
  output nblksiin2hjdghpd,   
  output cqss2zfmm9gkyqrwf,   
  output yamns_fbsulfpji691,   
  output hyram4bhtm3b2uv_2,   







  output odfbwv2n0hmkh9n2v ,
  output vqqbidi8kkzgxc0qls ,
  output ujg_tx8c5t9t0ddsmq ,
  output xxf9gqnuyu__15_t1u ,
  output f4uqn8qf5ljfnqy ,
  output k0kxgs4dhk1hf26ky3 ,
  output ngw96h2ls51cor4  ,
  output cj5vhekber5gw1509m86 ,
  output zouaj0qk3vke9quhfiqz ,
  output u3s5vk_sv9c1gjjto,
  output pm7lg8nzlruwwz9t29i ,
  output tffp7jbfj_acgbf_htp  ,
  output mbmpk0lgl7bqaq0m7j  ,
  output fkbmt37lnc1cbn6h7f5q  ,
  output uhs5rs3m1apmo4oj3c7  ,
  output hkzo9ego93d08t8igz2  ,
  
  
  
  
  output [64-1:0] so01tnkdju7vnwezjvi,
  output [64-1:0] hxad9091n05p_gjjo4,


  input  [64-1:0] uk0gax2bf5vv97rrbosr,

  input  gf33atgy,
  input  ru_wi
  );


  wire yc1860sc  = zojgfxfr_e4 [16:16 ];
  wire lu4q7um   = zojgfxfr_e4 [17:17  ];

  assign so01tnkdju7vnwezjvi  = lu4q7um  ? biu3jln6jgq  : dn0217a1asgpu;
  assign hxad9091n05p_gjjo4  = 
                            yc1860sc ? nlpn_dhtplj1_ : jzpnr2l6ruhz;

  wire opp2c8    = zojgfxfr_e4 [18:18 ] ;
  wire wao52c9  = zojgfxfr_e4 [19:19 ];
  wire djo84wp_5uy = zojgfxfr_e4 [20:20 ];
  wire cvok75_q    = zojgfxfr_e4 [21:21 ];


  assign odfbwv2n0hmkh9n2v  = zojgfxfr_e4 [5:5 ] & (~opp2c8) 
                            ;
  assign vqqbidi8kkzgxc0qls  = zojgfxfr_e4 [6:6 ];
  assign ujg_tx8c5t9t0ddsmq  = 
                            zojgfxfr_e4 [7:7 ];
  assign xxf9gqnuyu__15_t1u  = 
                            zojgfxfr_e4 [8:8 ];
  assign f4uqn8qf5ljfnqy  = 
                            zojgfxfr_e4 [9:9 ];
  assign k0kxgs4dhk1hf26ky3  = zojgfxfr_e4 [10:10 ];
  assign ngw96h2ls51cor4   = zojgfxfr_e4 [11:11  ];
  assign cj5vhekber5gw1509m86  = zojgfxfr_e4 [12:12 ];
  assign zouaj0qk3vke9quhfiqz  = zojgfxfr_e4 [13:13 ];
  assign u3s5vk_sv9c1gjjto = zojgfxfr_e4 [14:14];
  assign pm7lg8nzlruwwz9t29i  = zojgfxfr_e4 [15:15 ];

  assign tffp7jbfj_acgbf_htp  = zojgfxfr_e4 [42:42  ];
  assign mbmpk0lgl7bqaq0m7j  = zojgfxfr_e4 [43:43  ];
  assign fkbmt37lnc1cbn6h7f5q  = zojgfxfr_e4 [44:44  ];
  assign uhs5rs3m1apmo4oj3c7  = zojgfxfr_e4 [45:45  ];
  assign hkzo9ego93d08t8igz2  = zojgfxfr_e4 [46:46  ];
  
  
  
  

  assign r9hdxtws4mibgldl = c6cxk8927p4f;
  assign m2_8aknpfse = olti9ndjvk_sohpa;
  assign n67h_nt2we0os531a = 
                           uk0gax2bf5vv97rrbosr;

  assign cqss2zfmm9gkyqrwf  = wao52c9;   
  assign yamns_fbsulfpji691 = djo84wp_5uy;   
  assign hyram4bhtm3b2uv_2 = cvok75_q;   


  assign nblksiin2hjdghpd = cqss2zfmm9gkyqrwf | yamns_fbsulfpji691 | hyram4bhtm3b2uv_2
                        ;

endmodule






















module m0m7t4t8fpmv #(
 parameter hcl69mdlw0ykna4ue4_t1 = 1 
)(
  input t9b41sw5vpr,
  input bfo1il0du_,
  input gnb98c7tbqat,
  input w4kjodkdva03q,
  input zawjtr32pktig,
  input [48-1:0]  hy14_6z7grvldvw, 
  input scadliwzjp0l78srd9p,
  input w2h8uh3l463qbgqmv,

  input nrebzehsuam,
  input [64-1:0] bvzc7t76o17,

  input i7vhyhns, 
  input veibgbyke,
  input lu44s70ub62,
  input [64-1:0] yocn4o2zav, 


  input   tywculgjyor8ndw,



  input  rvr30vvllni,
  input  z1cj655u31,
  input  lhu2z948o3n,

  input  pw3qcykea5ib_ieka,
  input  g6xvfy8tj0zmajl ,



  input  jjzotrbn, 
  output hw1_k1jmu, 


  input  ryc6z1c7rmzrnlno, 


  input  [4-1:0] qbpmsk2,

  input  [64-1:0] tc88s6cm5b,
  input  [64-1:0] c3sszdooylrw,
  input  [3-1:0] vc529nuu,
  input  xh52jycxcjs,
  input  rnx27onf2lbe,
  output ya8t4ev_aidf0t0x4or,
  input  [64-1:0] l6s_gf8go82fwn,
  input  [64-1:0] afifdv1w9,
  input  [64-1:0] u2bhabgcppcy,
  input  [64-1:0] aziir_r1p,          

  input                           cj2osby26qlape,

  input  [64-1:0] b_sdf8,
  input  [31:0] n1rp2mggtiknd88,
  input  [64-1:0] begxws3d6mwhnm,
  input  [64-1:0] z1nw2lilgog_,
  input  [64-1:0] x6ywulzbb7jp,
  input b9mfhl8am_whqquz,
  input [19-1:0] bqen_oh1ujvq9lj4,
  input [105-1:0] e19iv2rqeu5,
  input [50-1:0] m4y6v4ncsg,
  input le3dqob2,
  input  [5-1:0] cpt0qfwiz,
  input [64-1:0]qpyjufa5h7y   ,
  input [64-1:0]hvv94pmafz   ,
  input j_rvclhfbeig5cqeb3_,
  input [64-1:0]sjunepbdn  ,
  input  [64-1:0] bwjyqadn,
  input  [64-1:0] binjv97px9r7dt04h0,
  input  o_d157fc5_l,
  input  ajl4tppx98ihuirj_mxih,
  input  [32-1:0] k0xug5g,
  input  ipht6ss_sh6h,
  input  [5-1:0] fhhe7189lmum,
  input  ojbpo5z6urt,
  input  q8977k41y4,
  input  ciiwo7qhifea,
  input  al4xeg8mukgfg,
  input  rhufxsnopy0n,
  input  wbhvg_1r9435,
  input  s1woka0byzgo,
  input  piwiqvrjoq,
  input  b7ilo27jne5k,
  input  u2k4dyp52s_m,
  input  djvj1e_,
  input  bktu0z1mk56,
  input  l6z1pzhjg5az,

  input  v35y3qnk7mx3l1695,

  output [27-1:0]      phofig8d5zd_8v9g8,     
  output [26-1:0]    js0ml55dtie8qenb4eoj2,
  output [64-1:0]                  p343qo1j,
  output [64-1:0]                  h8m3g7a,
  output                                   r9ix0zzks6zej,
  output                                   l8xeqkc,






  output                     gqe6zqljzhgt5wz98      ,
  output                     tisftwun8guh8lnibary2gz ,
  output                     wdgj6jexv3_u8sb4gnsv5 ,
  output                     c_qlgbc7oqwu9as946yqls ,
  output [64-1:0] nc5hf3a4mwl257q       ,
  output                     cqq719hbl6kax00mwmrhj   ,
  output                     a_x852mvzp7z5occs1   ,




  output  v3e6l1k7eo9k3 ,
  output  hxrmt706n071lic0f7,
  output lrhkvgg4x13sq245, 
  output [64-1:0] y45254ns5fjfjnwjiwr1_quk,
  output sshjsyphxbyaqk3kr,
  output mf10lk374lxu341vp3kpfl6,
  output isvwkofue95j9ud7p3nrgntc,
  output nkemiexuw_o6b34go,
  output bnnsit7f_1yqs20xcxk3l,
  output [64-1:0] c2vqeph9snojapvdushbj,

  output zu8yygom_ioh, 
  input  od8eje0yjk8, 
  output l_km9bow2ubqs5dtd,  
  output [64-1:0] cv8rkirz,  
  output [32-1:0] mbnh9clp6pd3t,  
  output [64-1:0]    z091v3i7q4_rty4,
  output w8wwz5822d7298zis7,
  output tsml_wqqwnty,      

  output pdz01l48nt,
  output l5zrepfg8it,
  output aq4b6s94dp0f,
  output dmg1a5xdc9 ,
  output v1j50zesdgxioc ,
  output tkhm63y407b,
  output nh1gz4628x89,
  output l4anyablbw3gt,
  output qhkm8drwygkskh_,
  output vn5b662w76_a3npe,
  output wigtf10_bybfdpp_x,
  output w2gbqib7zable3o,
  output zp24wdce6ufxkpbs,
  output xxee65tc1tureck,
  output wr1tfb0_sg9,
  output enhpakthwj3e65vldt,
  output mz47ksy6nekv1cbaq75,
  output egplp36i1ttcggdv2b0xo2e,
  output rbsutocgtudusq3v,
  output sgy1x259o9ltvsfe,
  output tr2dgjt2yqfzjaos9o,
  output [64-1:0] o8m475rdcb4y71zte3fbd30,
  output nzm80hh72kwblbx4fcg, 
  output l9wonwtwviy4i8w6s, 
  output wuw4k4dyuslqkjap, 
  output s4o6xx8w0dylrebxlqmia79t5, 

  output br6lhce3u3l01blvxzrqphj5svlum,
  output zq261z2pygzc0_h44fo,
  output g_w5s5kg5qk2w1gyo7odo2nubrxo0 ,
  output b1iduhkyfb7xynn3btxh6lhgev7_ ,
  output ndtc71v47ribx6u_eqsx8tdk0 ,
  output efp001u9ffq4ypu8uk4l8tbblt8 ,
  output fce921hmrlbrv4qdu4cb0pee ,
  output twjiv2hewisn6o,
  output l4i6kd5vs494chi,












  output [31:0] d7kpxfpyhil_2nt,








  output jugi02ecegnos3, 
  input  rxjuugktc38un, 
  output [64-1:0] h8wu7unf_ixmxfeh,
  output [5-1:0] b84l246u4jmnu,
  output uh251o1pav, 
  output [4-1:0] kdpgigzs75vcc1d  ,
  output vjkz8n6i44pc7o,     
  output cwmxezrc3jv6hzxcfc,
  input  uig3ujuyq0_61kqb,
  output xc2becmsn4fcniw6ks,
  output [64-1:0] nb3w1rq_ny95rvrt,
  output [4-1:0] p_yx415so7q1vohijb,

  output suxmggt9hea4ao3r,
  output kwn45x5pjj_5mi,
  output lp9c9xlhbpjow4k,
  output ts1jnweqrdhomp,
  output ze26d9sog9r3thx,






  
  
  output                        isz7jw04u7k3s7b398, 
  input                         q4_7fnx90rztwn6_8dybi, 
  output [64-1:0]       zq2e9j_emlri_qjtg,
  output                        qv749hsiom75nyn49v,
  output [4-1:0] gw6s_h2ymbn1ds50q8,
  
  
  output vo_fj58ip6ok0srq7t5, 
  input  qq819v1yyh8derngk15k1, 
  output [64-1:0] o_q0qt9vjpibgshm714a,
  output melkey3fxhhc3e649p,
  output [4-1:0] iqx3cqyh7_mpvu_9om,



  output rb050tnl,
  output a94vd35etec4,
  output el7_p8jit09,
  output [12-1:0] e1go3iu,

  input  af5qc04tmn51e4u2h1z,
  input  qwcb6hcmvfqmf032z,
  input  r0s7d8cr68i2qs1z,
  input  kakelc68be0x7tdm9b9o,
  input  j3j1czgoam48vhs8auo,
  input  gm1r5itc44uxw_y0_msk,
  input  [64-1:0] l9erxxpnphqd26vg9,
  input  [64-1:0] hig2gwwbeuhnt65xrp,
  output [64-1:0] guuvp01vkcryglsu1p3,
  output [64-1:0] vf5xcr67bqhzlo43_,

  output [64-1:0] vmx1fh4kmh4c,

  input  [64-1:0] zmfo8cca_77pc,
  output [64-1:0] bj7h5jqg66r51jxki6emra,























































  
  
  
  
  output v657dksgaz1cki9,
  output qzz1jhwf_vd0r8g, 
  input  dwn42a1uvd9x3myec, 
  output [4 -1:0] uiojikf9vcnz,
  output [64 -1:0] x1_k6oouttg7m3f,
  output [64 -1:0] fcvvhg9v3mx,
  output [64 -1:0] l_v5xmhbzqc,
  output [3-1:0] i7iq7ecm_d9pi6uw6,
  input  p5fn_ooo9rctbxkgm_jui,
  input  a5z_23_ryr_m29hhia_p ,



  input  gf33atgy,
  input  ru_wi
  );





  wire [64-1:0] yqs98coa39vu7;
  wire [64-1:0] cd0szp_7s1jnw;





  wire hnf_wyxvz1jn9wt8 = b7ilo27jne5k;  











  wire [48-1:0]  qsngsdmvoowsh = {48{t9b41sw5vpr}} & hy14_6z7grvldvw;
  wire [48-1:0]  f02j1_1eastxoh = {48{bfo1il0du_}} & hy14_6z7grvldvw;
  wire [48-1:0]  x8dt7e21kqfww7n = {48{gnb98c7tbqat}} & hy14_6z7grvldvw;
  wire [48-1:0]  tk5ngec81k = {48{w4kjodkdva03q}} & hy14_6z7grvldvw;


  wire j1we4o_jq6 = t9b41sw5vpr;
  wire bx89ng51ifc5n = bfo1il0du_;
  wire yas5k1_0cqxw9t = gnb98c7tbqat;
  wire n66q34nf3o1 = w4kjodkdva03q;

  wire cgn5_8ym11 = zawjtr32pktig;
  wire tgh4hil0u4nn0mih = cj2osby26qlape;
  wire gml_tzlxi8mv = cgn5_8ym11 | tgh4hil0u4nn0mih;

  wire qherdpqlgbhx1 = (~hnf_wyxvz1jn9wt8) & j1we4o_jq6 ;
  wire ei82smlw45m = qherdpqlgbhx1 & i7vhyhns;
  wire esr71bul94s1v = (~hnf_wyxvz1jn9wt8) & bx89ng51ifc5n;
  wire n3w1kpphj = esr71bul94s1v;
  wire bycddb3mhn1ga = (~hnf_wyxvz1jn9wt8) & yas5k1_0cqxw9t;
  wire khaw8p = bycddb3mhn1ga & lu44s70ub62;
  wire j61lgkdibp_nr8n = (~hnf_wyxvz1jn9wt8) & n66q34nf3o1;
  wire a7bzgrh = j61lgkdibp_nr8n;
  wire xt6eqjulr16w = le3dqob2;

  wire mxn4wdlge = (~hnf_wyxvz1jn9wt8) & xt6eqjulr16w;

  wire s66_nzq5i23lbo;
  wire v51v27wp_7tuha;
  wire isrgf76t7pxi;
  wire b7nkstim3k = (~hnf_wyxvz1jn9wt8) & cgn5_8ym11;
  wire cdlm5zrwv = (~hnf_wyxvz1jn9wt8) & tgh4hil0u4nn0mih;
  wire w86hm036xqu9hguo = b7nkstim3k | cdlm5zrwv;

  wire w93iw99udtpi6y = b9mfhl8am_whqquz;
  wire ft7ipo4vuxj = (~hnf_wyxvz1jn9wt8) & b9mfhl8am_whqquz;
  wire hvf_5lrj = ft7ipo4vuxj;
  wire opddptxe1    = bqen_oh1ujvq9lj4[5:5   ];
  wire rm85kx   = bqen_oh1ujvq9lj4[6:6  ];
  wire xt2jzmuzqs = bqen_oh1ujvq9lj4[7:7];
  wire w_wyjws0ma  = bqen_oh1ujvq9lj4[8:8 ];
  wire fm5qvc    = bqen_oh1ujvq9lj4[9:9   ];
  wire ms_4ed   = bqen_oh1ujvq9lj4[10:10  ];
  wire i7sstsvqw    = bqen_oh1ujvq9lj4[11:11   ];
  wire p4ggl84x_   = bqen_oh1ujvq9lj4[12:12  ];
  wire bu2stjoruwb  = bqen_oh1ujvq9lj4[14:14  ];
  wire vmw3ij0a96  = bqen_oh1ujvq9lj4[15:15  ];
  wire zt4egkm = bqen_oh1ujvq9lj4[16:16 ];
  wire wslud0u  = bqen_oh1ujvq9lj4[17:17  ];
  wire ujsqugs = bqen_oh1ujvq9lj4[18:18 ];
  wire wvr9_ddra61 = opddptxe1 | rm85kx | xt2jzmuzqs | w_wyjws0ma | bu2stjoruwb;
  wire yi3gmyct = fm5qvc | ms_4ed | i7sstsvqw    | p4ggl84x_ | vmw3ij0a96 | zt4egkm | wslud0u | ujsqugs;

  wire gifgw_z2iuu5s = w93iw99udtpi6y & wvr9_ddra61;
  wire e0tqa5udo7q_4 = w93iw99udtpi6y & yi3gmyct;
  wire zwzzi2nr = hvf_5lrj & wvr9_ddra61;
  wire ncphj0b = hvf_5lrj & yi3gmyct;
  wire xgpp07s3jj0vxd;
  generate
    if (hcl69mdlw0ykna4ue4_t1) begin: hp_2oabslchbydhgtobyfv4_
      assign xgpp07s3jj0vxd = (t9b41sw5vpr  & (~i7vhyhns)) 
                        | (gnb98c7tbqat & (~lu44s70ub62))
                        | w4kjodkdva03q 
                        | b9mfhl8am_whqquz
                        | zawjtr32pktig
                        | cj2osby26qlape
                        | le3dqob2
                        ;

    end else begin: yib8enrc4ileycrljs45
      assign xgpp07s3jj0vxd = (t9b41sw5vpr  & (~i7vhyhns)) 
                    | (gnb98c7tbqat & (~lu44s70ub62))


                    ;
    end
  endgenerate

  wire pz2bb_5njek = (~hnf_wyxvz1jn9wt8) & xgpp07s3jj0vxd;









  wire bwvpn4pm5q2m2 = jjzotrbn & zwzzi2nr;
  wire z4za08k83of9q = jjzotrbn & ncphj0b;
  wire ictx5fosbsup6y = jjzotrbn & mxn4wdlge;
  wire mt0f3958vekbx9 = jjzotrbn & w86hm036xqu9hguo;
  wire fj0lzkw_e2tjj = jjzotrbn & n3w1kpphj;
  wire c6cxk8927p4f = jjzotrbn & ei82smlw45m;
  wire fj5f6r_brv9 = jjzotrbn & khaw8p;
  wire v7t8ipf7s3pkl = jjzotrbn & a7bzgrh;
  wire fi816rwfszigkucl7ys = jjzotrbn & hnf_wyxvz1jn9wt8;
  wire dq_qnrmwcl6dcke = jjzotrbn & pz2bb_5njek;

  wire p7t1k5doyho;
  wire e79c5kbq9c5f;
  wire d9f119ap_n00k;
  wire x9a3z87q3adhgofd;
  wire im2j_m47n4mhs;
  wire m2_8aknpfse;
  wire kdpypaw_l038t;
  wire r30egqbrycq6277u;
  wire ycy6z9hc84ajgm9k;

  wire j6osee8dtbl;



  assign hw1_k1jmu =   ((im2j_m47n4mhs & n3w1kpphj)
                   | (e79c5kbq9c5f & zwzzi2nr)
                   | (d9f119ap_n00k & ncphj0b)
                   | (x9a3z87q3adhgofd & w86hm036xqu9hguo)
                   | (m2_8aknpfse & ei82smlw45m)
                   | (ycy6z9hc84ajgm9k & hnf_wyxvz1jn9wt8)
                   | (kdpypaw_l038t & khaw8p)
                   | (r30egqbrycq6277u & a7bzgrh)


                   | (p7t1k5doyho & pz2bb_5njek)
                   | (s66_nzq5i23lbo & mxn4wdlge)
                   )
                     ;


  wire ah6dvj4hwj480v;
  wire ogtxqxlymgsff9qr;
  wire i1517rq45m7oy8;






  wire sq6asp7q1ph0o1;   

  wire gm39_778;

  assign  {sq6asp7q1ph0o1, gm39_778} = 

                      ({1'b1,1'b0} & {2{ei82smlw45m}}) 

                    | ({1'b1,1'b0} & {2{a7bzgrh}}) 

                    | ({1'b1,1'b0} & {2{khaw8p}}) 

                    | ({1'b1,1'b0} & {2{pz2bb_5njek}}) 

                    | ({1'b1,1'b1} & {2{hnf_wyxvz1jn9wt8}}) 

                    | ({pw3qcykea5ib_ieka,g6xvfy8tj0zmajl} & {2{n3w1kpphj}}) 

                       
                    | ({2{ogtxqxlymgsff9qr}} & {2{ncphj0b}}) 
                    | ({2{ah6dvj4hwj480v}} & {2{zwzzi2nr}}) 
                    | ({~i1517rq45m7oy8, 1'b0} & {2{w86hm036xqu9hguo}}) 
                    | ({1'b0,1'b0} & {2{mxn4wdlge}})
                   ;







  wire                  lbd_qikbfejcglzz;
  wire                  g6j_bkwxdy36w;
  wire [64-1:0] vr1msvsauqfuz4s;

  assign lbd_qikbfejcglzz = dq_qnrmwcl6dcke;
  assign p7t1k5doyho = g6j_bkwxdy36w;
  assign vr1msvsauqfuz4s = ({64{~i7vhyhns}} & yocn4o2zav);








  wire wykc_imin5w;
  wire xnta372agn8z7;
  wire [64-1:0] b6nv94op09myrtj3wy;
  wire vp2vijaywqexo22ty08;



  wire  [64-1:0]           uhp5bzs36   = {64         {n66q34nf3o1}} & tc88s6cm5b;
  wire  [64-1:0]           b6rgihnhymh   = {64         {n66q34nf3o1}} & c3sszdooylrw;
  wire  [64-1:0]           gk0itvt5u   = {64         {n66q34nf3o1}} & b_sdf8;
  wire  [48-1:0]  nybrz2cz78r  = {48{n66q34nf3o1}} & tk5ngec81k;  
  wire                             gr47f0gunxy4e1c =                      n66q34nf3o1   & ojbpo5z6urt;  


  generate 
  if (hcl69mdlw0ykna4ue4_t1) begin: rlvc4ycafb809udjxpi5e

  xnt41w1r9gyu7e7lcjxkg92u wz81_gm5tcxyen17x0vxwk5hlmd7s(
    .tywculgjyor8ndw    (1'b0   ),                
    .w2h8uh3l463qbgqmv(1'b0),

    .aw82i964do(1'b0),
    .y8_gkxsfle(1'b0),
    .pydatzxqqi(1'b0),


    .v7t8ipf7s3pkl      (v7t8ipf7s3pkl),
    .r30egqbrycq6277u      (r30egqbrycq6277u),

    .uhp5bzs36        (64'h0),
    .nybrz2cz78r       (nybrz2cz78r[27-1:0]),
    .gr47f0gunxy4e1c      (1'b0),

    .rb050tnl          (rb050tnl           ),
    .e1go3iu          (e1go3iu           ),
    .el7_p8jit09        (el7_p8jit09         ),
    .a94vd35etec4        (a94vd35etec4         ),
    .l9erxxpnphqd26vg9     (64'h0                 ),
    .vf5xcr67bqhzlo43_     (vf5xcr67bqhzlo43_      ),
    .hig2gwwbeuhnt65xrp    (64'h0                 ),
    .guuvp01vkcryglsu1p3( guuvp01vkcryglsu1p3),
    .r0s7d8cr68i2qs1z  (1'b0),

    .vmx1fh4kmh4c          ( vmx1fh4kmh4c          ),

    .zmfo8cca_77pc    (64'h0    ), 
    .bj7h5jqg66r51jxki6emra(bj7h5jqg66r51jxki6emra),
    .wykc_imin5w      (wykc_imin5w      ),   
    .xnta372agn8z7      (xnta372agn8z7      ),   
    .b6nv94op09myrtj3wy  (b6nv94op09myrtj3wy  ),
    .vp2vijaywqexo22ty08   (vp2vijaywqexo22ty08   ),

    .gf33atgy             (gf33atgy),
    .ru_wi           (ru_wi)
  );
  end else begin: e2mwxe3ab9zc_1nlgpc463c

  xnt41w1r9gyu7e7lcjxkg92u z8n554ymjobf_kogxbvg448w76cu3i(
    .tywculgjyor8ndw    (tywculgjyor8ndw   ),
    .w2h8uh3l463qbgqmv(w2h8uh3l463qbgqmv),

    .aw82i964do(u2k4dyp52s_m),
    .y8_gkxsfle(djvj1e_),
    .pydatzxqqi(bktu0z1mk56),


    .v7t8ipf7s3pkl      (v7t8ipf7s3pkl),
    .r30egqbrycq6277u      (r30egqbrycq6277u),

    .uhp5bzs36        (uhp5bzs36  ),
    .nybrz2cz78r       (nybrz2cz78r[27-1:0]),
    .gr47f0gunxy4e1c      (gr47f0gunxy4e1c),

    .rb050tnl          (rb050tnl),
    .e1go3iu          (e1go3iu),
    .el7_p8jit09        (el7_p8jit09),
    .a94vd35etec4        (a94vd35etec4),
    .l9erxxpnphqd26vg9     (l9erxxpnphqd26vg9),
    .vf5xcr67bqhzlo43_     (vf5xcr67bqhzlo43_),
    .hig2gwwbeuhnt65xrp    (hig2gwwbeuhnt65xrp),
    .guuvp01vkcryglsu1p3(guuvp01vkcryglsu1p3),
    .r0s7d8cr68i2qs1z  (r0s7d8cr68i2qs1z),

    .vmx1fh4kmh4c          (vmx1fh4kmh4c),

    .zmfo8cca_77pc    (zmfo8cca_77pc),
    .bj7h5jqg66r51jxki6emra     (bj7h5jqg66r51jxki6emra),
    .wykc_imin5w      (wykc_imin5w      ),   
    .xnta372agn8z7      (xnta372agn8z7      ),   
    .b6nv94op09myrtj3wy  (b6nv94op09myrtj3wy  ),
    .vp2vijaywqexo22ty08   (vp2vijaywqexo22ty08   ),

    .gf33atgy             (gf33atgy),
    .ru_wi           (ru_wi)
  );
  end
  endgenerate





  wire c4znhmchls2i9; 
  wire fjclz58zhz4y4uf; 
  wire [64-1:0] e0lrg61pa8jctwey_k;
  wire [64-1:0] ldicihngwys9frt8r_q;
  wire ye3uidmavh9jbm9w4;
  wire ulpu2wlvtk0b4i;
  wire rb8jt7db79k4r076h;
  wire g4gfgb2tm_ujg9dhex;
  wire vyp0v8hghszoph ;
  wire uzn0rxbzurqxprl ;
  wire rz9jowsqb1lne29t6 ;
  wire uo8rfftroteg2gy267f;
  wire h8j00pdvikgalx01_;
  wire fxpfb14s16dp6ihm;
  wire njgro75dfrjo_60y;
  wire djpeelru7ruovogpcwr;
  wire f8c0swke1b88ml;
  wire hmbu9tiu4cl764c;

  wire [64-1:0] bm6cerfr_1bou52muqp;
  wire [64-1:0] tz3kfmltx71a5i0tmaln;
  wire b9asx2rffq8fclg3_q ;
  wire m1dubsueroj_o4i9hhxf ;
  wire vupdzhdsf5tcdbcy3br3 ;
  wire rzgzqvqbgh3abztkqck ;
  wire n9_mxfs9poavrerrqf3ps;
  wire a8ql4znkrbh_gj7cnnwc2j;
  wire tz95dh49670qhxle1;
  wire ehhimwdiwsd20nyinnomx;
  wire [64-1:0] todxu2rm67fxk1x8y_tl4;

  wire  [64-1:0]           d4lx9_3xlxjia1  = {64         {yas5k1_0cqxw9t}} & tc88s6cm5b;
  wire  [64-1:0]           pa1go4rk4_  = {64         {yas5k1_0cqxw9t}} & c3sszdooylrw;
  wire  [64-1:0]           tcdcik4o5zc  = {64         {yas5k1_0cqxw9t}} & bvzc7t76o17;
  wire  [48-1:0]  h1ieg8rrdd = {48{yas5k1_0cqxw9t}} & x8dt7e21kqfww7n;  
  wire  [64-1:0]        nl8lrzq7   = {64      {yas5k1_0cqxw9t}} & bwjyqadn;  




  generate 
  if (hcl69mdlw0ykna4ue4_t1) begin: j_jfy_pajdxuzfrcte18


     wire nu7hc86wz44pessqgvceajddmn3s;
     wire cj4f17jo0s_z9vmi5htht = nu7hc86wz44pessqgvceajddmn3s & (~qwcb6hcmvfqmf032z);
     wire a0itdy0a5fts62ldu_woafqynzc;
     wire zn5lc4nu61e0ms4p0u4v2siuxjz_6;
     wire r0nx0iuols_4pg0z96k6ifhert;
     wire [64-1:0] ztfuyixi1aw62ttyksukyd   ;
     wire d3vybluuijhl4u65a3wsn_n6i1;
     wire y0nferrzezge90_qml8ypux7i;

  iluwktw0594417cwb1su l9ut8gfoezyeajynt04fdqcy(
      .fj5f6r_brv9         (fj5f6r_brv9         ),
      .kdpypaw_l038t         (kdpypaw_l038t         ),
      .d4lx9_3xlxjia1           (d4lx9_3xlxjia1           ),
      .pa1go4rk4_           (pa1go4rk4_           ),
      .h1ieg8rrdd          (h1ieg8rrdd[34-1:0]),
      .tcdcik4o5zc           (tcdcik4o5zc           ),
      .nl8lrzq7            (nl8lrzq7            ),

      .c4znhmchls2i9         (c4znhmchls2i9  ),
      .fjclz58zhz4y4uf         (fjclz58zhz4y4uf  ),
      .e0lrg61pa8jctwey_k     (e0lrg61pa8jctwey_k  ),
      .ldicihngwys9frt8r_q    (ldicihngwys9frt8r_q ),
      .dytd_hd42_wbyvlhrmt9r7   (binjv97px9r7dt04h0    ),  
      .ye3uidmavh9jbm9w4        (ye3uidmavh9jbm9w4     ),
      .ulpu2wlvtk0b4i      (ulpu2wlvtk0b4i   ),

      .v3e6l1k7eo9k3        (v3e6l1k7eo9k3 ),
      .hxrmt706n071lic0f7       (hxrmt706n071lic0f7),
      .rb8jt7db79k4r076h       (rb8jt7db79k4r076h    ),
      .g4gfgb2tm_ujg9dhex      (g4gfgb2tm_ujg9dhex    ),
      .vyp0v8hghszoph       (vyp0v8hghszoph     ),
      .uzn0rxbzurqxprl       (uzn0rxbzurqxprl     ),
      .rz9jowsqb1lne29t6      (rz9jowsqb1lne29t6    ),
      .uo8rfftroteg2gy267f      (uo8rfftroteg2gy267f    ),
      .h8j00pdvikgalx01_      (h8j00pdvikgalx01_    ),
      .fxpfb14s16dp6ihm      (fxpfb14s16dp6ihm    ),
      .njgro75dfrjo_60y    (njgro75dfrjo_60y  ),
      .djpeelru7ruovogpcwr    (djpeelru7ruovogpcwr  ),
      .f8c0swke1b88ml      (f8c0swke1b88ml   ),
      .hmbu9tiu4cl764c      (hmbu9tiu4cl764c   ),

      .bm6cerfr_1bou52muqp     (bm6cerfr_1bou52muqp       ),
      .tz3kfmltx71a5i0tmaln     (tz3kfmltx71a5i0tmaln       ),
      .b9asx2rffq8fclg3_q  (b9asx2rffq8fclg3_q    ),
      .m1dubsueroj_o4i9hhxf  (m1dubsueroj_o4i9hhxf    ),
      .vupdzhdsf5tcdbcy3br3  (vupdzhdsf5tcdbcy3br3    ),
      .rzgzqvqbgh3abztkqck  (rzgzqvqbgh3abztkqck    ),
      .n9_mxfs9poavrerrqf3ps (n9_mxfs9poavrerrqf3ps   ),
      .a8ql4znkrbh_gj7cnnwc2j (a8ql4znkrbh_gj7cnnwc2j   ),
      .tz95dh49670qhxle1     (tz95dh49670qhxle1       ),
      .ehhimwdiwsd20nyinnomx (ehhimwdiwsd20nyinnomx   ),
      .todxu2rm67fxk1x8y_tl4 (todxu2rm67fxk1x8y_tl4   ),

      .gf33atgy                 (gf33atgy),
      .ru_wi               (ru_wi)
  );

  lqqd_zj04p6o3_g6h1le u_ux607_exu_branchslv(
    .r21i4by0bu3ks                   (2'b11),
    .ip4b_cj6h98z45oey8l           (1'b0),

    .w5rbttl5mj11z                 (), 
    .lu3guz5hxinmv_i4vg2k             (lrhkvgg4x13sq245    ),  
    .tbncz5fmqkrrvgqd9n8lz        (ldicihngwys9frt8r_q),
    .m5qoggt2in4ie_llz91            (ye3uidmavh9jbm9w4),

    .d2cosjdh8e6u1zldf6kf09           (o_d157fc5_l),
    .l9wonwtwviy4i8w6s            (l9wonwtwviy4i8w6s ), 
    .nwpj2xvetia76ai6nkrnv5k8cpxq   (br6lhce3u3l01blvxzrqphj5svlum),
    .xlzi1qrfl8ef8u0                  (pdz01l48nt    ),  
    .uiqmdx8tnsb                   (l5zrepfg8it     ),  
    .c9q9b8x3r05mpe5                  (aq4b6s94dp0f  ),  
    .ntedv1bjeakd                   (dmg1a5xdc9   ),  
    .i1a3ajcrp                   (v1j50zesdgxioc   ),  
    .wokc20mug9u1gn                  (tkhm63y407b  ),  
    .asl4zsbrnfn7                (1'b0),
    .psf3mvojppotcy                (1'b0),
    .yec_1lu2ooyq                  (1'b0  ),
    .hhimu5qv7me_z                  (1'b0  ),
    .bn3gk8oaq6g3ax                  (1'b0  ),
    .obqt4l21562rgtgxh              (1'b0  ),
    .otv3n61fdzkg6gt              (twjiv2hewisn6o),
    .bq_u11fb64d2bir3vxj              (l4i6kd5vs494chi),
    .sfs34sstg9pk                    (cv8rkirz      ),
    .c_fnucn4hvf3g               (z091v3i7q4_rty4),


    .l7r_xp04shn9v4n12        (al4xeg8mukgfg    ),
    .ouj04k7brubwkv_h9qhnkh    (ryc6z1c7rmzrnlno),
    .c00vdqa8yvwhd6r55g      (s1woka0byzgo   ),
    .lovkp0eqfnxtb7            (                        ),

    .rrujrlc85mhm            (                  ),
    .s_m3pbf5m2tr6v            (                  ),



    .jw4fsjecr0u919fr7            (                   ),
    .gfod0nmy6eta29jeeg6mr2      (s4o6xx8w0dylrebxlqmia79t5),
    .n4soswat5yihd74b         (wuw4k4dyuslqkjap),
    .y8wz7aud_fd6dfiakjtx2i0g   (mf10lk374lxu341vp3kpfl6),
    .a3xib90kwk4_hm1         (nkemiexuw_o6b34go),
    .nfzexr8q9g893gi          (bnnsit7f_1yqs20xcxk3l),
    .opkkwp3eg8g3448t         (c2vqeph9snojapvdushbj),
    .tv3_4qrynvnaoy4riz           (w8wwz5822d7298zis7),
    .pldoasxyzlvx2              ( 64'h0    ),


    .bde41te346q515l              ( 64'h0    ),
    .hn85hkp2yav               (  64'h0   ),

    .pydatzxqqi                (bktu0z1mk56),
    .aw82i964do                  (u2k4dyp52s_m),
    .rvr30vvllni              (rvr30vvllni),
    .y8_gkxsfle                  (djvj1e_),
    .z1cj655u31              (z1cj655u31),
    .lhu2z948o3n              (lhu2z948o3n),

    .glime27x19feqrvvsa2nmeh5f(1'b0),
    .llyh4o81vzcbw0zjekct       (1'b1    ),
    .mnqkmoietusiwyf95g       (nu7hc86wz44pessqgvceajddmn3s ), 
    .bq75f6k903dwxcstjv1wpw2cg09  (a0itdy0a5fts62ldu_woafqynzc),  
    .m1yqe0cmaq2_frcfgf_1c1qtgm7  (zn5lc4nu61e0ms4p0u4v2siuxjz_6),  
    .t2uejj01ae4b5d7shv4q2x  (r0nx0iuols_4pg0z96k6ifhert),  
    .sdsekm12iz4x32pwrh        (ztfuyixi1aw62ttyksukyd    ),  
    .tskef3o28v1jcu97th07m_    (d3vybluuijhl4u65a3wsn_n6i1),
    .nd7mxlwd9xekhy2oqb88dre5    (y0nferrzezge90_qml8ypux7i),  

    .gf33atgy   (gf33atgy  ),
    .ru_wi (ru_wi)
  );



  assign gqe6zqljzhgt5wz98      = cj4f17jo0s_z9vmi5htht;
  assign tisftwun8guh8lnibary2gz = a0itdy0a5fts62ldu_woafqynzc;
  assign wdgj6jexv3_u8sb4gnsv5 = zn5lc4nu61e0ms4p0u4v2siuxjz_6;
  assign c_qlgbc7oqwu9as946yqls = r0nx0iuols_4pg0z96k6ifhert;
  assign nc5hf3a4mwl257q       = ztfuyixi1aw62ttyksukyd;
  assign cqq719hbl6kax00mwmrhj   = d3vybluuijhl4u65a3wsn_n6i1;
  assign a_x852mvzp7z5occs1   = y0nferrzezge90_qml8ypux7i;
  assign isvwkofue95j9ud7p3nrgntc = cj4f17jo0s_z9vmi5htht;

  end else begin: e_firlcc7jrw9z_h9
  iluwktw0594417cwb1su ahq2gjyu63kizw98qpp5qvr(
      .fj5f6r_brv9         (fj5f6r_brv9 ),
      .kdpypaw_l038t         (kdpypaw_l038t ),
      .d4lx9_3xlxjia1           (d4lx9_3xlxjia1           ),
      .pa1go4rk4_           (pa1go4rk4_           ),
      .h1ieg8rrdd          (h1ieg8rrdd[34-1:0]),
      .tcdcik4o5zc           (tcdcik4o5zc           ),
      .nl8lrzq7            (nl8lrzq7            ),

      .c4znhmchls2i9         (c4znhmchls2i9      ),
      .fjclz58zhz4y4uf         (fjclz58zhz4y4uf      ),
      .e0lrg61pa8jctwey_k     (e0lrg61pa8jctwey_k  ),
      .ldicihngwys9frt8r_q    (ldicihngwys9frt8r_q ),
      .dytd_hd42_wbyvlhrmt9r7   (binjv97px9r7dt04h0    ),  
      .ye3uidmavh9jbm9w4        (ye3uidmavh9jbm9w4     ),
      .ulpu2wlvtk0b4i      (ulpu2wlvtk0b4i   ),

      .v3e6l1k7eo9k3        (v3e6l1k7eo9k3 ),
      .hxrmt706n071lic0f7       (hxrmt706n071lic0f7),
      .rb8jt7db79k4r076h       (rb8jt7db79k4r076h    ),
      .g4gfgb2tm_ujg9dhex      (g4gfgb2tm_ujg9dhex    ),
      .vyp0v8hghszoph       (vyp0v8hghszoph     ),
      .uzn0rxbzurqxprl       (uzn0rxbzurqxprl     ),
      .rz9jowsqb1lne29t6      (rz9jowsqb1lne29t6    ),
      .uo8rfftroteg2gy267f      (uo8rfftroteg2gy267f    ),
      .fxpfb14s16dp6ihm      (fxpfb14s16dp6ihm    ),
      .h8j00pdvikgalx01_      (h8j00pdvikgalx01_    ),
      .njgro75dfrjo_60y    (njgro75dfrjo_60y  ),
      .djpeelru7ruovogpcwr    (djpeelru7ruovogpcwr  ),
      .f8c0swke1b88ml      (f8c0swke1b88ml   ),
      .hmbu9tiu4cl764c      (hmbu9tiu4cl764c   ),

      .bm6cerfr_1bou52muqp     (bm6cerfr_1bou52muqp       ),
      .tz3kfmltx71a5i0tmaln     (tz3kfmltx71a5i0tmaln       ),
      .b9asx2rffq8fclg3_q  (b9asx2rffq8fclg3_q    ),
      .m1dubsueroj_o4i9hhxf  (m1dubsueroj_o4i9hhxf    ),
      .vupdzhdsf5tcdbcy3br3  (vupdzhdsf5tcdbcy3br3    ),
      .rzgzqvqbgh3abztkqck  (rzgzqvqbgh3abztkqck    ),
      .n9_mxfs9poavrerrqf3ps (n9_mxfs9poavrerrqf3ps   ),
      .a8ql4znkrbh_gj7cnnwc2j (a8ql4znkrbh_gj7cnnwc2j   ),
      .tz95dh49670qhxle1     (tz95dh49670qhxle1       ),
      .ehhimwdiwsd20nyinnomx (ehhimwdiwsd20nyinnomx   ),
      .todxu2rm67fxk1x8y_tl4 (todxu2rm67fxk1x8y_tl4   ),

      .gf33atgy                 (gf33atgy),
      .ru_wi               (ru_wi)
  );


  assign gqe6zqljzhgt5wz98    = 1'b0;
  assign tisftwun8guh8lnibary2gz = 1'b0;
  assign wdgj6jexv3_u8sb4gnsv5 = 1'b0;
  assign c_qlgbc7oqwu9as946yqls = 1'b0;
  assign nc5hf3a4mwl257q       = 64'h0;
  assign cqq719hbl6kax00mwmrhj   = 1'b0;
  assign a_x852mvzp7z5occs1   = 1'b0;
  assign l9wonwtwviy4i8w6s = 1'b0; 
  assign wuw4k4dyuslqkjap = 1'b0; 
  assign mf10lk374lxu341vp3kpfl6 = 1'b0;
  assign s4o6xx8w0dylrebxlqmia79t5 = 1'b0; 
  assign isvwkofue95j9ud7p3nrgntc = 1'b0;
  assign nkemiexuw_o6b34go = 1'b0;
  assign bnnsit7f_1yqs20xcxk3l = 1'b0;
  assign c2vqeph9snojapvdushbj = 64'b0;
  assign w8wwz5822d7298zis7 = 1'b0;



  end
  endgenerate






  wire hgt2urny9_9; 
  wire nrxcyc791r8gksao; 
















    wire [64-1:0] tp6hfcjxcyp899mpksjl;
    wire [64-1:0] f4ds8dbk9kk_ic_;
    wire                  xl9r7gr7wciuv2d00b ;
    wire [64-1:0] ttgsydregi0kgoj_z;



  wire  [64-1:0]           c5lrjuy9t_f  = {64         {bx89ng51ifc5n}} & tc88s6cm5b;
  wire  [64-1:0]           bi9zhg2zyeg  = {64         {bx89ng51ifc5n}} & c3sszdooylrw;
  wire  [64-1:0]           iet1_xpdj  = {64         {bx89ng51ifc5n}} & b_sdf8;
  wire  [48-1:0]  ybrrs0__m1aa00 = {48{bx89ng51ifc5n}} & f02j1_1eastxoh;  
  wire  [4-1:0]     jythgzdjfospqb = {4   {bx89ng51ifc5n}} & qbpmsk2;  

  wire pkwcaygsgot_59n1  = bx89ng51ifc5n & u2k4dyp52s_m;
  wire vy1aysleh0imu4  = bx89ng51ifc5n & djvj1e_;
  wire pbjk7minp0n89j  = bx89ng51ifc5n & bktu0z1mk56;
  wire b4uk5z2pu_0s = bx89ng51ifc5n & l6z1pzhjg5az;

  wire  [64-1:0] q02_ci8ru207_lx;
  generate 
  if (hcl69mdlw0ykna4ue4_t1) begin: l_4ic6e8kjn4rc1ja2xb
  n9fwcab7kdqyokfwizktfw  gaw1808otgpaa6hnszair2fy(

      .fj0lzkw_e2tjj         (fj0lzkw_e2tjj     ),
      .im2j_m47n4mhs         (im2j_m47n4mhs     ),
      .c5lrjuy9t_f           (c5lrjuy9t_f       ),
      .bi9zhg2zyeg           (bi9zhg2zyeg       ),
      .yqs98coa39vu7           (yqs98coa39vu7       ),
      .cd0szp_7s1jnw           (cd0szp_7s1jnw       ),
      .iet1_xpdj           (iet1_xpdj       ),
      .utdfnsgxzrzt14u          (aziir_r1p),
      .ybrrs0__m1aa00          (ybrrs0__m1aa00),

      .jythgzdjfospqb          (jythgzdjfospqb      ),
      .pkwcaygsgot_59n1         (pkwcaygsgot_59n1     ),
      .vy1aysleh0imu4         (vy1aysleh0imu4     ),
      .pbjk7minp0n89j         (pbjk7minp0n89j     ),
      .b4uk5z2pu_0s        (b4uk5z2pu_0s    ),

      .hgt2urny9_9         (hgt2urny9_9         ),
      .nrxcyc791r8gksao         (nrxcyc791r8gksao         ),

      .tp6hfcjxcyp899mpksjl     (tp6hfcjxcyp899mpksjl     ),
      .f4ds8dbk9kk_ic_     (f4ds8dbk9kk_ic_     ),
      .xl9r7gr7wciuv2d00b     (xl9r7gr7wciuv2d00b     ),
      .ttgsydregi0kgoj_z     (ttgsydregi0kgoj_z     ),

      .gf33atgy                 (gf33atgy),
      .ru_wi               (ru_wi)
  );

  assign q02_ci8ru207_lx   = ttgsydregi0kgoj_z; 
















































end  else begin: aiq2_9u5umsbcmigx

  assign q02_ci8ru207_lx = 64'h0;

  assign hgt2urny9_9  = fj0lzkw_e2tjj; 
  assign im2j_m47n4mhs  = nrxcyc791r8gksao;




































  assign tp6hfcjxcyp899mpksjl = 64'h0;
  assign f4ds8dbk9kk_ic_ = 64'h0;
  assign xl9r7gr7wciuv2d00b = 1'b0;                




























  end
  endgenerate




  wire r9hdxtws4mibgldl; 
  wire olti9ndjvk_sohpa; 
  wire [64-1:0] n67h_nt2we0os531a;
  wire nblksiin2hjdghpd;   
  wire cqss2zfmm9gkyqrwf;
  wire yamns_fbsulfpji691;
  wire hyram4bhtm3b2uv_2;

  wire odfbwv2n0hmkh9n2v ;
  wire vqqbidi8kkzgxc0qls ;
  wire ujg_tx8c5t9t0ddsmq ;
  wire xxf9gqnuyu__15_t1u ;
  wire f4uqn8qf5ljfnqy ;
  wire k0kxgs4dhk1hf26ky3 ;
  wire ngw96h2ls51cor4  ;
  wire cj5vhekber5gw1509m86 ;
  wire zouaj0qk3vke9quhfiqz ;
  wire u3s5vk_sv9c1gjjto;
  wire pm7lg8nzlruwwz9t29i ;
  wire tffp7jbfj_acgbf_htp  ;
  wire mbmpk0lgl7bqaq0m7j  ;
  wire fkbmt37lnc1cbn6h7f5q  ;
  wire uhs5rs3m1apmo4oj3c7  ;
  wire hkzo9ego93d08t8igz2  ;
  wire [64-1:0] so01tnkdju7vnwezjvi;
  wire [64-1:0] hxad9091n05p_gjjo4;

  wire [64-1:0] uk0gax2bf5vv97rrbosr;

  wire  [64-1:0]           dn0217a1asgpu  =  {64         {j1we4o_jq6}} & tc88s6cm5b;
  wire  [64-1:0]           jzpnr2l6ruhz  =  {64         {j1we4o_jq6}} & c3sszdooylrw;
  wire  [64-1:0]           nlpn_dhtplj1_  =  {64         {j1we4o_jq6}} & b_sdf8;
  wire  [48-1:0]  zojgfxfr_e4 =  {48{j1we4o_jq6}} & qsngsdmvoowsh;  
  wire  [64-1:0]        biu3jln6jgq   =  {64      {j1we4o_jq6}} & bwjyqadn;  


  q8buuqlskug7714mfcon71 nvb1tn63mvz1n_hu659d(

      .c6cxk8927p4f         (c6cxk8927p4f     ),
      .m2_8aknpfse         (m2_8aknpfse     ),
      .dn0217a1asgpu           (dn0217a1asgpu           ),
      .jzpnr2l6ruhz           (jzpnr2l6ruhz           ),
      .zojgfxfr_e4          (zojgfxfr_e4[47-1:0]),
      .nlpn_dhtplj1_           (nlpn_dhtplj1_           ),
      .biu3jln6jgq            (biu3jln6jgq            ),

      .r9hdxtws4mibgldl         (r9hdxtws4mibgldl         ),
      .olti9ndjvk_sohpa         (olti9ndjvk_sohpa         ),
      .n67h_nt2we0os531a     (n67h_nt2we0os531a     ),
      .nblksiin2hjdghpd      (nblksiin2hjdghpd      ),
      .cqss2zfmm9gkyqrwf     (cqss2zfmm9gkyqrwf     ),
      .yamns_fbsulfpji691    (yamns_fbsulfpji691    ),
      .hyram4bhtm3b2uv_2       (hyram4bhtm3b2uv_2       ),

      .odfbwv2n0hmkh9n2v     (odfbwv2n0hmkh9n2v       ),
      .vqqbidi8kkzgxc0qls     (vqqbidi8kkzgxc0qls       ),
      .ujg_tx8c5t9t0ddsmq     (ujg_tx8c5t9t0ddsmq       ),
      .xxf9gqnuyu__15_t1u     (xxf9gqnuyu__15_t1u       ),
      .f4uqn8qf5ljfnqy     (f4uqn8qf5ljfnqy       ),
      .k0kxgs4dhk1hf26ky3     (k0kxgs4dhk1hf26ky3       ),
      .ngw96h2ls51cor4      (ngw96h2ls51cor4        ),
      .cj5vhekber5gw1509m86     (cj5vhekber5gw1509m86       ),
      .zouaj0qk3vke9quhfiqz     (zouaj0qk3vke9quhfiqz       ),
      .u3s5vk_sv9c1gjjto    (u3s5vk_sv9c1gjjto      ),
      .pm7lg8nzlruwwz9t29i     (pm7lg8nzlruwwz9t29i       ),
      .tffp7jbfj_acgbf_htp    (tffp7jbfj_acgbf_htp      ),
      .mbmpk0lgl7bqaq0m7j    (mbmpk0lgl7bqaq0m7j      ),
      .fkbmt37lnc1cbn6h7f5q    (fkbmt37lnc1cbn6h7f5q      ),
      .uhs5rs3m1apmo4oj3c7    (uhs5rs3m1apmo4oj3c7      ),
      .hkzo9ego93d08t8igz2    (hkzo9ego93d08t8igz2      ),
      .so01tnkdju7vnwezjvi     (so01tnkdju7vnwezjvi       ),
      .hxad9091n05p_gjjo4     (hxad9091n05p_gjjo4       ),
      .uk0gax2bf5vv97rrbosr     (uk0gax2bf5vv97rrbosr       ),

      .gf33atgy                 (gf33atgy           ),
      .ru_wi               (ru_wi         ) 
  );


  
  
  
  
  wire [64-1:0]           loc9a4t09i4  = begxws3d6mwhnm;
  wire [64-1:0]           k2jxyry72hc9nl  = z1nw2lilgog_;
  wire [64-1:0]           xtlt33xlczy37q  = x6ywulzbb7jp;
  wire [19-1:0]  uzxs4linfwcrjy = bqen_oh1ujvq9lj4;  
  wire  [4-1:0]    t86na4x45h4ficw = qbpmsk2;  

  wire i_swuedh0b3s; 
  wire qvhs4kakyng1sk; 



  
  
  
  

  generate
  if (hcl69mdlw0ykna4ue4_t1) begin: q_m7ocsob2lizblb6kenunv4ro
  vnidphqictr3gtptdwbgr os3lyxvkdsazef54hkw_3pb (

      .bwvpn4pm5q2m2            (1'b0), 
      .e79c5kbq9c5f            (e79c5kbq9c5f), 

      .loc9a4t09i4              (64'b0      ),
      .k2jxyry72hc9nl              (64'b0      ),
      .xtlt33xlczy37q              (xtlt33xlczy37q      ),
      .uzxs4linfwcrjy             (uzxs4linfwcrjy[19-1:0]),

      .ah6dvj4hwj480v         (ah6dvj4hwj480v ),
      .t86na4x45h4ficw             (t86na4x45h4ficw     ),

      .i_swuedh0b3s            (i_swuedh0b3s),
      .qvhs4kakyng1sk            (qvhs4kakyng1sk),

      .baeb5atyeipjmjtwdx66m       (vo_fj58ip6ok0srq7t5), 
      .zf3zgw37xlcc2o5eprc5k       (qq819v1yyh8derngk15k1), 
      .a9rvmf7a9nbie6nd923        (o_q0qt9vjpibgshm714a),
      .gzyfsm1lj5vk008         (melkey3fxhhc3e649p),   
      .w6xoq8do9qo8kitx8e        (iqx3cqyh7_mpvu_9om),


      .gf33atgy                    (gf33atgy            ),
      .ru_wi                  (ru_wi          ) 
  );
  end else begin: ivau4plyjjazjyn1z_ikvxibk
  vnidphqictr3gtptdwbgr os3lyxvkdsazef54hkw_3pb (

      .bwvpn4pm5q2m2            (bwvpn4pm5q2m2), 
      .e79c5kbq9c5f            (e79c5kbq9c5f), 

      .loc9a4t09i4              (loc9a4t09i4      ),
      .k2jxyry72hc9nl              (k2jxyry72hc9nl      ),
      .xtlt33xlczy37q              (xtlt33xlczy37q      ),
      .uzxs4linfwcrjy             (uzxs4linfwcrjy[19-1:0]),

      .ah6dvj4hwj480v         (ah6dvj4hwj480v ),
      .t86na4x45h4ficw             (t86na4x45h4ficw     ),

      .i_swuedh0b3s            (i_swuedh0b3s),
      .qvhs4kakyng1sk            (qvhs4kakyng1sk),

      .baeb5atyeipjmjtwdx66m       (vo_fj58ip6ok0srq7t5), 
      .zf3zgw37xlcc2o5eprc5k       (qq819v1yyh8derngk15k1), 
      .a9rvmf7a9nbie6nd923        (o_q0qt9vjpibgshm714a),
      .gzyfsm1lj5vk008         (melkey3fxhhc3e649p),   
      .w6xoq8do9qo8kitx8e        (iqx3cqyh7_mpvu_9om),


      .gf33atgy                    (gf33atgy            ),
      .ru_wi                  (ru_wi          ) 
  );
  end
  endgenerate

  
  
  
  wire [64-1:0]           dq0a9sotg74w  = {64         {e0tqa5udo7q_4}} & begxws3d6mwhnm;
  wire [64-1:0]           netnmrvccmf  = {64         {e0tqa5udo7q_4}} & z1nw2lilgog_;
  wire [64-1:0]           qaxmne8xc_  = {64         {e0tqa5udo7q_4}} & x6ywulzbb7jp;
  wire [19-1:0]  v48iyoy1fdeh = {19{e0tqa5udo7q_4}} & bqen_oh1ujvq9lj4;  
  wire  [4-1:0]    gcl2zxzh4brhr = {4   {e0tqa5udo7q_4}} & qbpmsk2;  

  wire jfgbmn4y_79lt81; 
  wire tsa8otson44it2;
  wire [64-1:0] du9nxa6qo7knx2et1gw6;
  wire h7szh92q4s7x6vx_;

  generate
  if (hcl69mdlw0ykna4ue4_t1) begin: re1y7nl_9ivvawq53vjo
  a3zxpqwwtl53hi anbbns1qjybpcxm6(
      .z4za08k83of9q      (1'b0    ),
      .d9f119ap_n00k      (d9f119ap_n00k    ),
       
      .dq0a9sotg74w        (64'h0 ),
      .netnmrvccmf        (64'h0 ),
      .qaxmne8xc_        (64'h0 ),
      .v48iyoy1fdeh       ({19{1'b0}}),
      .ogtxqxlymgsff9qr   (ogtxqxlymgsff9qr ),
      .gcl2zxzh4brhr       (4'h0),
                          
      .jfgbmn4y_79lt81      (jfgbmn4y_79lt81    ),
      .tsa8otson44it2      (tsa8otson44it2    ),
      .du9nxa6qo7knx2et1gw6  (du9nxa6qo7knx2et1gw6),
      .h7szh92q4s7x6vx_   (h7szh92q4s7x6vx_ ),

      .isz7jw04u7k3s7b398(isz7jw04u7k3s7b398),
      .q4_7fnx90rztwn6_8dybi(1'b0),
      .zq2e9j_emlri_qjtg (zq2e9j_emlri_qjtg),
      .qv749hsiom75nyn49v  (qv749hsiom75nyn49v ),
      .gw6s_h2ymbn1ds50q8 (gw6s_h2ymbn1ds50q8),

      .gf33atgy              (gf33atgy            ),
      .ru_wi            (ru_wi          ) 

  );
  end else begin: td2_e_jkendk04g9d
  a3zxpqwwtl53hi anbbns1qjybpcxm6(

      .z4za08k83of9q      (z4za08k83of9q    ),
      .d9f119ap_n00k      (d9f119ap_n00k    ),
       
      .dq0a9sotg74w        (dq0a9sotg74w      ),
      .netnmrvccmf        (netnmrvccmf      ),
      .qaxmne8xc_        (qaxmne8xc_      ),
      .v48iyoy1fdeh       (v48iyoy1fdeh[19-1:0]),
      .ogtxqxlymgsff9qr   (ogtxqxlymgsff9qr ),
      .gcl2zxzh4brhr       (gcl2zxzh4brhr     ),
                          
      .jfgbmn4y_79lt81      (jfgbmn4y_79lt81    ),
      .tsa8otson44it2      (tsa8otson44it2    ),
      .du9nxa6qo7knx2et1gw6  (du9nxa6qo7knx2et1gw6),
      .h7szh92q4s7x6vx_   (h7szh92q4s7x6vx_ ),

      .isz7jw04u7k3s7b398(isz7jw04u7k3s7b398),
      .q4_7fnx90rztwn6_8dybi(q4_7fnx90rztwn6_8dybi),
      .zq2e9j_emlri_qjtg (zq2e9j_emlri_qjtg),
      .qv749hsiom75nyn49v  (qv749hsiom75nyn49v ),
      .gw6s_h2ymbn1ds50q8 (gw6s_h2ymbn1ds50q8),

      .gf33atgy              (gf33atgy            ),
      .ru_wi            (ru_wi          ) 
  );
  end
  endgenerate



  wire c0z4i4kyokyx7sug; 
  wire w2kcsfod60d_68;
  wire [64-1:0] ntu21o6bz2w2777k4u;
  wire ffyib96xpww6adq;
  wire owq8xep05y1_39287n92;
  
generate
if (hcl69mdlw0ykna4ue4_t1) begin: fyk1k_6pctrhbnvw5f3pe
  assign c0z4i4kyokyx7sug = 1'b0; 
  assign x9a3z87q3adhgofd = w2kcsfod60d_68;
  assign ntu21o6bz2w2777k4u = {64{1'b0}};
  assign ffyib96xpww6adq = 1'b0;
  assign owq8xep05y1_39287n92 = 1'b0;
  
  assign v657dksgaz1cki9   = 1'b0;
  assign qzz1jhwf_vd0r8g = 1'b0;
  assign uiojikf9vcnz  = {4-1{1'b0}};
  assign x1_k6oouttg7m3f   = {64{1'b0}};
  assign fcvvhg9v3mx   = {64{1'b0}};
  assign l_v5xmhbzqc   = {64{1'b0}};
  assign i7iq7ecm_d9pi6uw6 = 3'b0;
  assign ya8t4ev_aidf0t0x4or = 1'b0;
  assign i1517rq45m7oy8 = 1'b0;


end else begin: qaj528xmf_nxaos6
  
  
  
  
  wire  [4-1:0]    lefkd05cxbpmfb = {4{gml_tzlxi8mv}} & qbpmsk2;  
  wire  [64-1:0]          wvg6yggd3_ngr  = l6s_gf8go82fwn;  
  wire  [64-1:0]          fvamtne5n7  = afifdv1w9;  
  wire  [64-1:0]          w6fv3puuz49wu  = u2bhabgcppcy;  
  wire  [3-1:0]                   ahi4ptho3r9  = {3{gml_tzlxi8mv}} & vc529nuu;
  wire                            tvy3ej4fztwicmyr  = gml_tzlxi8mv & xh52jycxcjs;

  wire esw3r2fugnssgn13j4;

  assign ya8t4ev_aidf0t0x4or = esw3r2fugnssgn13j4
                          | (j1we4o_jq6 & af5qc04tmn51e4u2h1z & xh52jycxcjs) 
                          ;



  ybdbqemjrr2kv71i ck_5yw2o4r7850yg(
      .rnx27onf2lbe       (rnx27onf2lbe),
      .ya8t4ev_aidf0t0x4or (esw3r2fugnssgn13j4),

      .af5qc04tmn51e4u2h1z (af5qc04tmn51e4u2h1z),

      .mt0f3958vekbx9      (mt0f3958vekbx9    ),
      .x9a3z87q3adhgofd      (x9a3z87q3adhgofd    ),
       
      .i1517rq45m7oy8   (i1517rq45m7oy8 ),
      .lefkd05cxbpmfb       (lefkd05cxbpmfb     ),
      .wvg6yggd3_ngr        (wvg6yggd3_ngr      ),
      .fvamtne5n7        (fvamtne5n7      ),
      .w6fv3puuz49wu        (w6fv3puuz49wu      ),
      .ahi4ptho3r9      (ahi4ptho3r9    ),
      .tvy3ej4fztwicmyr      (tvy3ej4fztwicmyr    ),
                          
      .c0z4i4kyokyx7sug      (c0z4i4kyokyx7sug    ),
      .w2kcsfod60d_68      (w2kcsfod60d_68    ),
      .ntu21o6bz2w2777k4u  (ntu21o6bz2w2777k4u),
      .ffyib96xpww6adq   (ffyib96xpww6adq ),
      .owq8xep05y1_39287n92(owq8xep05y1_39287n92),

      .v657dksgaz1cki9      (v657dksgaz1cki9   ),
      .qzz1jhwf_vd0r8g    (qzz1jhwf_vd0r8g ),
      .dwn42a1uvd9x3myec    (dwn42a1uvd9x3myec ),
      .uiojikf9vcnz     (uiojikf9vcnz  ),
      .x1_k6oouttg7m3f      (x1_k6oouttg7m3f   ),
      .fcvvhg9v3mx      (fcvvhg9v3mx   ),
      .l_v5xmhbzqc      (l_v5xmhbzqc   ),
      .i7iq7ecm_d9pi6uw6    (i7iq7ecm_d9pi6uw6   ),
      .p5fn_ooo9rctbxkgm_jui (p5fn_ooo9rctbxkgm_jui),
      .a5z_23_ryr_m29hhia_p(a5z_23_ryr_m29hhia_p),

      .gf33atgy              (gf33atgy            ),
      .ru_wi            (ru_wi          ) 
  );


  end
endgenerate






  
  wire r_aei1gc7v37oo9dghv; 
  wire d1_eg4gq3uyxdyycybx;
  wire [64-1:0] od3rbv8xxz65lrcy;
  wire [64-1:0] du4qneuo7c4380bw33j;
  wire [64-1:0] m2s376x2ngd1fz27iofg3yf1;
  wire [64-1:0] f2mrhq1ax6cmfmtx_l5;
  wire hgdur8q6gk2ak91b = (r_aei1gc7v37oo9dghv | d1_eg4gq3uyxdyycybx) & xt6eqjulr16w;

  
  
  
  
  wire  [4-1:0] ker4nfxz2b_p53w = {4{xt6eqjulr16w}} & qbpmsk2;  




generate
if (hcl69mdlw0ykna4ue4_t1) begin: v93e2vcumx2a1vun_e

  
  assign r_aei1gc7v37oo9dghv = 1'b0; 
  assign d1_eg4gq3uyxdyycybx = 1'b0;
  assign od3rbv8xxz65lrcy = {64{1'b0}};
  assign du4qneuo7c4380bw33j = {64{1'b0}};


  assign vjkz8n6i44pc7o           = 1'b0;     
  assign cwmxezrc3jv6hzxcfc  = 1'b0;
  assign xc2becmsn4fcniw6ks    = 1'b0;
  assign nb3w1rq_ny95rvrt   = {64{1'b0}}; 
  assign p_yx415so7q1vohijb = {4{1'b0}};



  assign v51v27wp_7tuha = 1'b0;
  assign s66_nzq5i23lbo = isrgf76t7pxi;


end else begin: vyxfknvdh1syinun2v

  rkhmkn86ap95zo99 ig2zt6006mogto63df9qge7 (
      .artnbioj                         ( qpyjufa5h7y                      ),
      .emfjxicm                         ( hvv94pmafz                      ),
      .ehzolf0                          ( sjunepbdn                   ),
      .fhhe7189lmum                       ( fhhe7189lmum                    ),
      .cpt0qfwiz                      ( cpt0qfwiz                   ), 
      .ker4nfxz2b_p53w                    ( ker4nfxz2b_p53w           ),
      .vjkz8n6i44pc7o                 ( vjkz8n6i44pc7o              ),  
      .cwmxezrc3jv6hzxcfc              ( cwmxezrc3jv6hzxcfc     ), 
      .uig3ujuyq0_61kqb              ( uig3ujuyq0_61kqb     ), 
      .nb3w1rq_ny95rvrt               ( nb3w1rq_ny95rvrt      ),
      .xc2becmsn4fcniw6ks                ( xc2becmsn4fcniw6ks       ),
      .p_yx415so7q1vohijb               ( p_yx415so7q1vohijb      ),
      .j_rvclhfbeig5cqeb3_             ( j_rvclhfbeig5cqeb3_          ),
      .e19iv2rqeu5                    ( e19iv2rqeu5                 ),
      .m4y6v4ncsg                    ( m4y6v4ncsg                 ),
      .wkzq9xwwp9c3wcf3616c             ( r_aei1gc7v37oo9dghv            ), 
      .juy4d3jn2_92c7jefm1i6             ( d1_eg4gq3uyxdyycybx            ), 
      .qebmlqd6ka70065zibcx             ( od3rbv8xxz65lrcy            ),
      .hftmbp4yfjjsgcltu             ( du4qneuo7c4380bw33j            ),
      .iont49tufvh5v7eetbw0m         ( m2s376x2ngd1fz27iofg3yf1        ),
      .u2yurbi1gylta0pv_xpnz8ppo         ( f2mrhq1ax6cmfmtx_l5        ),

      .ictx5fosbsup6y                   (ictx5fosbsup6y),
      .s66_nzq5i23lbo                   (s66_nzq5i23lbo),
                                                             
      .v51v27wp_7tuha                   (v51v27wp_7tuha),
      .isrgf76t7pxi                   (isrgf76t7pxi),
                                                       
      .gf33atgy                           (gf33atgy                        ), 
      .ru_wi                         (ru_wi                      )
    );
  end
endgenerate








  wire ktu3yhilgxp = j1we4o_jq6;
  wire fv0c5k6cjre = yas5k1_0cqxw9t;
  wire yvw7xod98x7 = bx89ng51ifc5n;

  wn2t_67c13cwq1_8a6 hnddk5wg7l5nzt535efo(
      .ktu3yhilgxp         (ktu3yhilgxp           ),    
      .odfbwv2n0hmkh9n2v     (odfbwv2n0hmkh9n2v       ),
      .vqqbidi8kkzgxc0qls     (vqqbidi8kkzgxc0qls       ),
      .ujg_tx8c5t9t0ddsmq     (ujg_tx8c5t9t0ddsmq       ),
      .xxf9gqnuyu__15_t1u     (xxf9gqnuyu__15_t1u       ),
      .f4uqn8qf5ljfnqy     (f4uqn8qf5ljfnqy       ),
      .k0kxgs4dhk1hf26ky3     (k0kxgs4dhk1hf26ky3       ),
      .ngw96h2ls51cor4      (ngw96h2ls51cor4        ),
      .cj5vhekber5gw1509m86     (cj5vhekber5gw1509m86       ),
      .zouaj0qk3vke9quhfiqz     (zouaj0qk3vke9quhfiqz       ),
      .u3s5vk_sv9c1gjjto    (u3s5vk_sv9c1gjjto      ),
      .pm7lg8nzlruwwz9t29i     (pm7lg8nzlruwwz9t29i       ),
      .tffp7jbfj_acgbf_htp    (tffp7jbfj_acgbf_htp     ),
      .mbmpk0lgl7bqaq0m7j    (mbmpk0lgl7bqaq0m7j     ),
      .fkbmt37lnc1cbn6h7f5q    (fkbmt37lnc1cbn6h7f5q     ),
      .uhs5rs3m1apmo4oj3c7    (uhs5rs3m1apmo4oj3c7     ),
      .hkzo9ego93d08t8igz2    (hkzo9ego93d08t8igz2     ),
      .so01tnkdju7vnwezjvi     (so01tnkdju7vnwezjvi       ),
      .hxad9091n05p_gjjo4     (hxad9091n05p_gjjo4       ),
      .uk0gax2bf5vv97rrbosr     (uk0gax2bf5vv97rrbosr       ),

      .fv0c5k6cjre         (fv0c5k6cjre           ),
      .bm6cerfr_1bou52muqp     (bm6cerfr_1bou52muqp       ),
      .tz3kfmltx71a5i0tmaln     (tz3kfmltx71a5i0tmaln       ),
      .b9asx2rffq8fclg3_q  (b9asx2rffq8fclg3_q    ),
      .m1dubsueroj_o4i9hhxf  (m1dubsueroj_o4i9hhxf    ),
      .vupdzhdsf5tcdbcy3br3  (vupdzhdsf5tcdbcy3br3    ),
      .rzgzqvqbgh3abztkqck  (rzgzqvqbgh3abztkqck    ),
      .n9_mxfs9poavrerrqf3ps (n9_mxfs9poavrerrqf3ps   ),
      .a8ql4znkrbh_gj7cnnwc2j (a8ql4znkrbh_gj7cnnwc2j   ),
      .tz95dh49670qhxle1     (tz95dh49670qhxle1       ),
      .ehhimwdiwsd20nyinnomx (ehhimwdiwsd20nyinnomx   ),
      .todxu2rm67fxk1x8y_tl4 (todxu2rm67fxk1x8y_tl4   ),

      .yvw7xod98x7         (yvw7xod98x7           ),
      .tp6hfcjxcyp899mpksjl     (tp6hfcjxcyp899mpksjl       ),
      .f4ds8dbk9kk_ic_     (f4ds8dbk9kk_ic_       ),
      .oso3fj0gx6pnvjni    (1'b0      ),
      .xl9r7gr7wciuv2d00b     (xl9r7gr7wciuv2d00b       ),
      .htcsb0affil7c6q     (1'b0      ),
      .vrqdq7uwxf99gj_7      (1'b0      ),
      .jqgtsdtxss_uios07     (1'b0      ),
      .hn2h_gkqinydwsdg_i3     (1'b0      ),
      .re8hncw6m47hrh6     (1'b0      ),
      .tshku7fgpiu2j7ugwjj9    (1'b0      ),
      .arc8ztjel_qlz3xfw0ya    (1'b0      ),
      .dukom1hk2mc9i6m4      (1'b1      ),
      .ttgsydregi0kgoj_z     (ttgsydregi0kgoj_z       ),
             
      .e__67e1k5hdb4ctnr       (1'b0         ),
      .jay_5c6ndpwhj0vqzv       (64'b0         ),
      .kn6tx97_rw9w0v         (),
            
      .nc_3q2q5fz4e2       (1'b0         ),
      .a5y809wbv8w1d0       (64'b0         ),
      .l0vxn4vg6wd         (),      


      .hgdur8q6gk2ak91b         (hgdur8q6gk2ak91b       ),    
      .r_aei1gc7v37oo9dghv     (r_aei1gc7v37oo9dghv   ),    
      .d1_eg4gq3uyxdyycybx     (d1_eg4gq3uyxdyycybx   ),    
      .od3rbv8xxz65lrcy     (od3rbv8xxz65lrcy   ),
      .du4qneuo7c4380bw33j     (du4qneuo7c4380bw33j   ),
      .m2s376x2ngd1fz27iofg3yf1 (m2s376x2ngd1fz27iofg3yf1   ),
      .f2mrhq1ax6cmfmtx_l5 (f2mrhq1ax6cmfmtx_l5   ),


      .gf33atgy                 (gf33atgy           ),
      .ru_wi               (ru_wi         ) 
    );


  wire bdmoj3mcktel1_qus3;
  wire lab1_4glh2j8sgkl6pofw;
  wire [64-1:0] alitplyh4w0svbs48nie1m;
  wire r0a9ex23qxn7tddwq0ip;

  assign ycy6z9hc84ajgm9k = lab1_4glh2j8sgkl6pofw;
  assign bdmoj3mcktel1_qus3 = fi816rwfszigkucl7ys;
  assign alitplyh4w0svbs48nie1m = 64'b0;
  assign r0a9ex23qxn7tddwq0ip  = 1'b1;




  wire l55er67nkdneeatw =   (khaw8p      & c4znhmchls2i9     );

  wire l7076zhst5 = (ei82smlw45m      & r9hdxtws4mibgldl     )
               | (khaw8p      & c4znhmchls2i9     )
               | (a7bzgrh      & wykc_imin5w     )
               | (n3w1kpphj      & hgt2urny9_9     )
               | (hnf_wyxvz1jn9wt8 & bdmoj3mcktel1_qus3)
                | (zwzzi2nr      & i_swuedh0b3s     )
                | (ncphj0b      & jfgbmn4y_79lt81     )
               | (mxn4wdlge & v51v27wp_7tuha)
               | (w86hm036xqu9hguo  & c0z4i4kyokyx7sug     )
               | (pz2bb_5njek      & lbd_qikbfejcglzz     )
               ;
























  assign lab1_4glh2j8sgkl6pofw = hnf_wyxvz1jn9wt8 & j6osee8dtbl;
  assign olti9ndjvk_sohpa      = ei82smlw45m & j6osee8dtbl;
  assign nrxcyc791r8gksao      = n3w1kpphj & j6osee8dtbl;
  assign qvhs4kakyng1sk      = zwzzi2nr & j6osee8dtbl;
  assign tsa8otson44it2      = ncphj0b & j6osee8dtbl;

  assign isrgf76t7pxi      = mxn4wdlge & j6osee8dtbl;

  assign g6j_bkwxdy36w      = pz2bb_5njek & j6osee8dtbl;

  assign w2kcsfod60d_68      = w86hm036xqu9hguo & j6osee8dtbl;
  assign fjclz58zhz4y4uf      = khaw8p & j6osee8dtbl;
  assign xnta372agn8z7      = a7bzgrh & j6osee8dtbl;


  wire [64-1:0] lojt0eer4uu4n07ak = 
                    ({64{ei82smlw45m}} & n67h_nt2we0os531a)
                  | ({64{khaw8p}} & e0lrg61pa8jctwey_k)
                  | ({64{a7bzgrh}} & b6nv94op09myrtj3wy)



                  | ({64{n3w1kpphj}} & q02_ci8ru207_lx)



                   | ({64{1'b0}})




                  | ({64{hnf_wyxvz1jn9wt8}} & alitplyh4w0svbs48nie1m)
                  ;


  wire [64-1:0] a9bvrwjinrx843zuzb6j5rueh = 
                    ({64{~pz2bb_5njek}} & {{64-64{1'b0}},lojt0eer4uu4n07ak})
                  | ({64{pz2bb_5njek}} & vr1msvsauqfuz4s);

  assign kdpgigzs75vcc1d   = qbpmsk2
                  ;

  assign h8wu7unf_ixmxfeh  = a9bvrwjinrx843zuzb6j5rueh; 
  assign b84l246u4jmnu = fhhe7189lmum; 

  wire v2cyf3u556m3fjzy4; 

  wire t62tpit597ljt = ojbpo5z6urt;
























































  wire a16omkrimdk  = 1'b1
                   ;



  wire jn9dck0_w7__ = n3w1kpphj | ncphj0b 
                     | zwzzi2nr 
                   ; 


wire e45zjh64jxwnli64ak; 
wire ngiuqj2j6rsgfaeu27  ; 

generate
  if (hcl69mdlw0ykna4ue4_t1 == 1) begin:sy346h1s7rulrjo


    assign  e45zjh64jxwnli64ak = l7076zhst5;
    assign  ngiuqj2j6rsgfaeu27   = 1'b0; 
  end else begin:j6r2_lpg87d4bn07bk



    assign e45zjh64jxwnli64ak = sq6asp7q1ph0o1 & l7076zhst5 & (a16omkrimdk  ? od8eje0yjk8  : 1'b1);
    assign ngiuqj2j6rsgfaeu27   = t62tpit597ljt & (~gm39_778) & (~tywculgjyor8ndw);
  end
endgenerate

  assign v2cyf3u556m3fjzy4 = rxjuugktc38un; 
  assign jugi02ecegnos3 = e45zjh64jxwnli64ak;
  assign uh251o1pav   = ngiuqj2j6rsgfaeu27;

generate
  if (hcl69mdlw0ykna4ue4_t1 == 1) begin:zxqb74w0wu6kgtfxyg

    assign j6osee8dtbl =  rxjuugktc38un; 

    assign zu8yygom_ioh  = 1'b0;
  end else begin:ta_6d3t7dcz4xjg8
    assign j6osee8dtbl = 
           (a16omkrimdk  ? od8eje0yjk8  : 1'b1)  
         & (sq6asp7q1ph0o1 ? rxjuugktc38un : 1'b1); 
    assign zu8yygom_ioh  = a16omkrimdk  & l7076zhst5 & (sq6asp7q1ph0o1 ? rxjuugktc38un : 1'b1);
  end
endgenerate

generate
  if (hcl69mdlw0ykna4ue4_t1 == 1) begin:nq8zh79xxbecmmhdb9ft5y
    assign lrhkvgg4x13sq245  = l55er67nkdneeatw & rxjuugktc38un;
  end else begin:qe7uc419gj96zm0g9vjyur5d
    assign lrhkvgg4x13sq245  = a16omkrimdk & l55er67nkdneeatw & (sq6asp7q1ph0o1 ? rxjuugktc38un : 1'b1);
  end
endgenerate

  assign y45254ns5fjfjnwjiwr1_quk =  ldicihngwys9frt8r_q;
  assign sshjsyphxbyaqk3kr = ye3uidmavh9jbm9w4;      


  assign mbnh9clp6pd3t   = k0xug5g;  
  assign tsml_wqqwnty   = bktu0z1mk56;
  assign cv8rkirz   = bwjyqadn;  
  assign z091v3i7q4_rty4  = bvzc7t76o17;
  assign pdz01l48nt = nrebzehsuam;







  assign l_km9bow2ubqs5dtd      =







                              ipht6ss_sh6h;





  assign d7kpxfpyhil_2nt   = n1rp2mggtiknd88;














  assign l5zrepfg8it         = khaw8p & rb8jt7db79k4r076h;
  assign aq4b6s94dp0f        = khaw8p & g4gfgb2tm_ujg9dhex;
  assign dmg1a5xdc9         = khaw8p & vyp0v8hghszoph ;
  assign v1j50zesdgxioc         = khaw8p & uzn0rxbzurqxprl ;
  assign tkhm63y407b        = khaw8p & rz9jowsqb1lne29t6;
  assign nh1gz4628x89        = khaw8p & uo8rfftroteg2gy267f;
  assign l4anyablbw3gt        = khaw8p & h8j00pdvikgalx01_;
  assign qhkm8drwygkskh_        = khaw8p & fxpfb14s16dp6ihm;
  assign twjiv2hewisn6o    = khaw8p & f8c0swke1b88ml;
  assign l4i6kd5vs494chi    = khaw8p & hmbu9tiu4cl764c;
  assign w2gbqib7zable3o      = khaw8p & njgro75dfrjo_60y;
  assign zp24wdce6ufxkpbs      = khaw8p & djpeelru7ruovogpcwr;
  assign xxee65tc1tureck    = (hnf_wyxvz1jn9wt8 & bdmoj3mcktel1_qus3 & s1woka0byzgo); 

  assign vn5b662w76_a3npe       = ei82smlw45m & cqss2zfmm9gkyqrwf;
  assign wigtf10_bybfdpp_x      = ei82smlw45m & yamns_fbsulfpji691;
  assign wr1tfb0_sg9         = ei82smlw45m & hyram4bhtm3b2uv_2;
  assign enhpakthwj3e65vldt = piwiqvrjoq;
  assign mz47ksy6nekv1cbaq75  = al4xeg8mukgfg;
  assign egplp36i1ttcggdv2b0xo2e = ryc6z1c7rmzrnlno;
  assign rbsutocgtudusq3v  = rhufxsnopy0n;
  assign sgy1x259o9ltvsfe  = wbhvg_1r9435;
  assign tr2dgjt2yqfzjaos9o  = s1woka0byzgo;
  assign o8m475rdcb4y71zte3fbd30 =  binjv97px9r7dt04h0;
  assign nzm80hh72kwblbx4fcg = o_d157fc5_l;
  assign br6lhce3u3l01blvxzrqphj5svlum =  ajl4tppx98ihuirj_mxih;
  assign zq261z2pygzc0_h44fo   = q8977k41y4
                           | (w86hm036xqu9hguo & owq8xep05y1_39287n92) 
                           | (w86hm036xqu9hguo & scadliwzjp0l78srd9p) 
                           | (n3w1kpphj & scadliwzjp0l78srd9p) 
                           | (a7bzgrh & r0s7d8cr68i2qs1z)
                        ;
  assign g_w5s5kg5qk2w1gyo7odo2nubrxo0 = q8977k41y4 & (~ciiwo7qhifea);
  assign b1iduhkyfb7xynn3btxh6lhgev7_ = q8977k41y4 &   ciiwo7qhifea;
  assign ndtc71v47ribx6u_eqsx8tdk0   = a7bzgrh & r0s7d8cr68i2qs1z & kakelc68be0x7tdm9b9o;
  assign efp001u9ffq4ypu8uk4l8tbblt8   = a7bzgrh & r0s7d8cr68i2qs1z & j3j1czgoam48vhs8auo;
  assign fce921hmrlbrv4qdu4cb0pee   = a7bzgrh & r0s7d8cr68i2qs1z & gm1r5itc44uxw_y0_msk;







  assign suxmggt9hea4ao3r    = qherdpqlgbhx1;
  assign kwn45x5pjj_5mi    = esr71bul94s1v;
  assign lp9c9xlhbpjow4k    = bycddb3mhn1ga;
  assign ts1jnweqrdhomp    = j61lgkdibp_nr8n;

  assign ze26d9sog9r3thx = ft7ipo4vuxj;

generate
  if (hcl69mdlw0ykna4ue4_t1) begin: c6lnj8z1h74v17v822xl3x_9ix
    assign  phofig8d5zd_8v9g8       = q02_ci8ru207_lx[27-1+12 : 12];
    assign  js0ml55dtie8qenb4eoj2 = q02_ci8ru207_lx[64-1 : 27+12-1];
    assign  p343qo1j             = yqs98coa39vu7;
    assign  h8m3g7a             = cd0szp_7s1jnw;
    assign  r9ix0zzks6zej       = 1'b0;
    assign  l8xeqkc               = f02j1_1eastxoh[11:11] || f02j1_1eastxoh[6:6];
  end
  else begin: f7p4e703s8jwvygbwg7x9zfg
    assign  phofig8d5zd_8v9g8       = 27'b0;
    assign  js0ml55dtie8qenb4eoj2 = 26'b0;
    assign  p343qo1j             = 64'b0;
    assign  h8m3g7a             = 64'b0;
    assign  r9ix0zzks6zej       = 1'b0;
    assign  l8xeqkc               = 1'b0;
    assign  yqs98coa39vu7           = 64'b0;
    assign  cd0szp_7s1jnw           = 64'b0;
  end

endgenerate






  wire sdnnqw20be9le = zu8yygom_ioh & od8eje0yjk8;
  wire vg5fg43b18k = 
                   sdnnqw20be9le & ( 
                      (~pw3qcykea5ib_ieka & n3w1kpphj) 

                       
                    | (ncphj0b) 
                    | (zwzzi2nr) 
                    | (w86hm036xqu9hguo) 
                    | (mxn4wdlge)
                  ) ; 

endmodule                                      




































module sneku_08a9mn2xq1ql88_9w6 #(
    parameter xa6g65id = 65
)(
    input  [2:0]        x, 
    input  [xa6g65id-1:0]  y, 
    output [xa6g65id:0]    iyeq5, 
    output              ugjvcvd2l_
    );















    assign ugjvcvd2l_ = x[2];
    assign iyeq5 = {(xa6g65id+1){x == 3'b000}} & {(xa6g65id+1){1'b0}}
              | {(xa6g65id+1){x == 3'b001}} & {y[xa6g65id-1],y}
              | {(xa6g65id+1){x == 3'b010}} & {y[xa6g65id-1],y}
              | {(xa6g65id+1){x == 3'b011}} & {y,1'b0}
              | {(xa6g65id+1){x == 3'b100}} & {~y,1'b1}
              | {(xa6g65id+1){x == 3'b101}} & {~y[xa6g65id-1],~y}
              | {(xa6g65id+1){x == 3'b110}} & {~y[xa6g65id-1],~y}
              | {(xa6g65id+1){x == 3'b111}} & {(xa6g65id+1){1'b1}}
              ;





endmodule

module l3hw_f8igiui51siqdj #(
  parameter onr7l = 106 
)(
  input [onr7l-1:0] frgfco,
  input [onr7l-1:0] ii,
  input [onr7l-1:0] fij51v,
  output [onr7l-1:0] c,
  output [onr7l-1:0] s 
);

assign s = (frgfco ^ ii) ^ fij51v;

wire [onr7l-1:0] oz7_y5 = (frgfco & ii) | (frgfco & fij51v) | (ii & fij51v);

assign c = {oz7_y5[onr7l-2:0], 1'b0};

endmodule


module mm88fxnds62ofbh80 #(
    parameter onr7l = 106 
)(
  input [onr7l-1:0] frgfco,
  input [onr7l-1:0] ii,
  input [onr7l-1:0] fij51v,
  input [onr7l-1:0] cuzhl9,
  output [onr7l-1:0] c,
  output [onr7l-1:0] s 
);

   wire [onr7l-1:0] i885 = (frgfco & ii) | (ii & fij51v) | (frgfco & fij51v);
   wire [onr7l-1:0] smqrocit = {i885[onr7l-2:0], 1'b0};

   wire [onr7l-1:0] tqxp_8 = smqrocit ^ cuzhl9;
   wire [onr7l-1:0] ddaxu87 = (frgfco ^ ii) ^ fij51v;

   assign s = tqxp_8 ^ ddaxu87;

   wire [onr7l-1:0] hgtxv = (ddaxu87 & cuzhl9) |  (cuzhl9 & smqrocit) | (smqrocit & ddaxu87);

   assign c = {hgtxv[onr7l-2:0], 1'b0};

endmodule

























module lqqd_zj04p6o3_g6h1le(

  input  ip4b_cj6h98z45oey8l,

  input [2-1:0] r21i4by0bu3ks,

  input  lu3guz5hxinmv_i4vg2k,  
  input  [64-1:0] tbncz5fmqkrrvgqd9n8lz,
  input  m5qoggt2in4ie_llz91,
  input  d2cosjdh8e6u1zldf6kf09,
  output l9wonwtwviy4i8w6s, 
  input  nwpj2xvetia76ai6nkrnv5k8cpxq,
  output w5rbttl5mj11z,
  input  xlzi1qrfl8ef8u0,  
  input  bn3gk8oaq6g3ax,
  input  yec_1lu2ooyq,
  input  hhimu5qv7me_z,
  input  asl4zsbrnfn7,
  input  psf3mvojppotcy,
  input  obqt4l21562rgtgxh,
  input  uiqmdx8tnsb,  
  input  c9q9b8x3r05mpe5,  
  input  ntedv1bjeakd ,  
  input  i1a3ajcrp,  
  input  wokc20mug9u1gn,  
  input  otv3n61fdzkg6gt,
  input  bq_u11fb64d2bir3vxj,
  input  [64-1:0] sfs34sstg9pk,  
  input  [64-1:0] c_fnucn4hvf3g,

  input  l7r_xp04shn9v4n12,
  input  ouj04k7brubwkv_h9qhnkh,
  input  c00vdqa8yvwhd6r55g,
  output [64-1:0] lovkp0eqfnxtb7,


  input  [64-1:0] pldoasxyzlvx2,
  input  [64-1:0] bde41te346q515l,
  input  [64-1:0] hn85hkp2yav,

  input  aw82i964do,
  input  rvr30vvllni,
  input  z1cj655u31,
  input  y8_gkxsfle,
  input  lhu2z948o3n,
  input  pydatzxqqi,

  input  glime27x19feqrvvsa2nmeh5f,
  input  llyh4o81vzcbw0zjekct,
  output mnqkmoietusiwyf95g,


  output bq75f6k903dwxcstjv1wpw2cg09,  
  output m1yqe0cmaq2_frcfgf_1c1qtgm7,  
  output t2uejj01ae4b5d7shv4q2x,  
  output [64-1:0] sdsekm12iz4x32pwrh,  
  output tskef3o28v1jcu97th07m_,  
  output nd7mxlwd9xekhy2oqb88dre5,  


  output rrujrlc85mhm,
  output s_m3pbf5m2tr6v,
  output jw4fsjecr0u919fr7,
  output n4soswat5yihd74b,
  output gfod0nmy6eta29jeeg6mr2,
  output y8wz7aud_fd6dfiakjtx2i0g, 
  output a3xib90kwk4_hm1,
  output nfzexr8q9g893gi,
  output [64-1:0] opkkwp3eg8g3448t,
  output tv3_4qrynvnaoy4riz,


  input  gf33atgy,
  input  ru_wi
  );

  wire qvu7q5ec5s706083i7burd;
  wire brchmis_flush_req_pre;

  assign mnqkmoietusiwyf95g = brchmis_flush_req_pre ;
  assign qvu7q5ec5s706083i7burd = llyh4o81vzcbw0zjekct ;






  wire o6r2xec3_010m1kq = nwpj2xvetia76ai6nkrnv5k8cpxq &  m5qoggt2in4ie_llz91;
  wire xj5aw3zada2vzo7c = uiqmdx8tnsb & (otv3n61fdzkg6gt ^ bq_u11fb64d2bir3vxj);
  assign tv3_4qrynvnaoy4riz = uiqmdx8tnsb & bq_u11fb64d2bir3vxj;
  wire rc8qiqhp68leip00pn = c9q9b8x3r05mpe5 & (~i1a3ajcrp);
  assign nfzexr8q9g893gi = i1a3ajcrp & (~wokc20mug9u1gn) & lu3guz5hxinmv_i4vg2k; 
  assign a3xib90kwk4_hm1 = (~i1a3ajcrp) & wokc20mug9u1gn & lu3guz5hxinmv_i4vg2k; 
  assign y8wz7aud_fd6dfiakjtx2i0g = (i1a3ajcrp ^ wokc20mug9u1gn) & lu3guz5hxinmv_i4vg2k & mnqkmoietusiwyf95g;
  wire vmt1l92s4l4avu9hn6sw = rc8qiqhp68leip00pn & lu3guz5hxinmv_i4vg2k; 
  assign l9wonwtwviy4i8w6s = d2cosjdh8e6u1zldf6kf09 & rc8qiqhp68leip00pn;  
  assign gfod0nmy6eta29jeeg6mr2 = vmt1l92s4l4avu9hn6sw & o6r2xec3_010m1kq & d2cosjdh8e6u1zldf6kf09; 
  assign n4soswat5yihd74b = vmt1l92s4l4avu9hn6sw & (~d2cosjdh8e6u1zldf6kf09);
  wire zyy78w5a8r5d3zks5fys = (
         xj5aw3zada2vzo7c  

       | o6r2xec3_010m1kq 

       | asl4zsbrnfn7 
  
       | psf3mvojppotcy

       | yec_1lu2ooyq 
       | hhimu5qv7me_z 

       | bn3gk8oaq6g3ax 

       | obqt4l21562rgtgxh 
      );

  wire a57pg701_3knwklw = (
         uiqmdx8tnsb 
       | asl4zsbrnfn7 
       | psf3mvojppotcy
       | yec_1lu2ooyq 
       | hhimu5qv7me_z 
       | obqt4l21562rgtgxh 
       | bn3gk8oaq6g3ax 
      );

  assign brchmis_flush_req_pre = lu3guz5hxinmv_i4vg2k & zyy78w5a8r5d3zks5fys;
















  assign bq75f6k903dwxcstjv1wpw2cg09 = bn3gk8oaq6g3ax ? (r21i4by0bu3ks == 2'b11) :    
                                  yec_1lu2ooyq ? rvr30vvllni : 
                                  hhimu5qv7me_z ? 1'b0 :       
                                 (asl4zsbrnfn7 | otv3n61fdzkg6gt) ? aw82i964do : 
                                  psf3mvojppotcy ? aw82i964do :       
                                  obqt4l21562rgtgxh ? aw82i964do :       
                                      aw82i964do;

  assign m1yqe0cmaq2_frcfgf_1c1qtgm7 = bn3gk8oaq6g3ax ? (r21i4by0bu3ks == 2'b01) :    
                                  yec_1lu2ooyq ? z1cj655u31 : 
                                  hhimu5qv7me_z ? lhu2z948o3n : 
                                 (asl4zsbrnfn7 | otv3n61fdzkg6gt) ? y8_gkxsfle : 
                                  psf3mvojppotcy ? y8_gkxsfle :       
                                  obqt4l21562rgtgxh ? y8_gkxsfle :       
                                      y8_gkxsfle;


  assign t2uejj01ae4b5d7shv4q2x = bn3gk8oaq6g3ax ? 1'b0 :    
                                  yec_1lu2ooyq ? pydatzxqqi : 
                                  hhimu5qv7me_z ? pydatzxqqi : 
                                 (asl4zsbrnfn7 | otv3n61fdzkg6gt) ? pydatzxqqi : 
                                  psf3mvojppotcy ? pydatzxqqi :       
                                  obqt4l21562rgtgxh ? pydatzxqqi : 
                                      pydatzxqqi;

  assign opkkwp3eg8g3448t =  sfs34sstg9pk + (xlzi1qrfl8ef8u0 ? 64'd4 : 64'd2);
  assign lovkp0eqfnxtb7 =  
                        sfs34sstg9pk + (
                            (

                              l7r_xp04shn9v4n12 ? ( ouj04k7brubwkv_h9qhnkh ? 64'd0 : 64'd2) :
                             ( (xlzi1qrfl8ef8u0 
                               )
                             ) ? 64'd4 : 64'd2
                            )
                        );

      
  assign sdsekm12iz4x32pwrh = 
                                
                          (obqt4l21562rgtgxh) ? sfs34sstg9pk :
                          (asl4zsbrnfn7 | (uiqmdx8tnsb & (~c9q9b8x3r05mpe5) & otv3n61fdzkg6gt)) ? lovkp0eqfnxtb7 :
                          (psf3mvojppotcy) ? lovkp0eqfnxtb7 :
    
                          (uiqmdx8tnsb & (~c9q9b8x3r05mpe5) & (~otv3n61fdzkg6gt)) ? (sfs34sstg9pk + c_fnucn4hvf3g[64-1:0]) :
                          (uiqmdx8tnsb ) ?  tbncz5fmqkrrvgqd9n8lz :  
                          bn3gk8oaq6g3ax ? hn85hkp2yav :
                          hhimu5qv7me_z ? bde41te346q515l :
                                       pldoasxyzlvx2 ;
                          
                          
                          
                          
                                                  
  assign tskef3o28v1jcu97th07m_ = asl4zsbrnfn7; 
  assign nd7mxlwd9xekhy2oqb88dre5 = psf3mvojppotcy; 

  wire yc7lxuu8auz6j7jn908az73 = mnqkmoietusiwyf95g & llyh4o81vzcbw0zjekct;
  assign rrujrlc85mhm = yec_1lu2ooyq & yc7lxuu8auz6j7jn908az73 & (~ip4b_cj6h98z45oey8l);
  assign s_m3pbf5m2tr6v = hhimu5qv7me_z & yc7lxuu8auz6j7jn908az73 & (~ip4b_cj6h98z45oey8l);



  assign jw4fsjecr0u919fr7 = bn3gk8oaq6g3ax & yc7lxuu8auz6j7jn908az73 & (~ip4b_cj6h98z45oey8l);

  assign w5rbttl5mj11z = (~a57pg701_3knwklw) | 
                             (




                                qvu7q5ec5s706083i7burd  



                             );

endmodule                                      
























module ycwy7frvptowq59s2 (
  output btwmhh91h50d5flgwx4o6pwu,

  input   feq1g7m2cy1erl,

  input   se2buoxmq91dbic3y2m5hu,
  output  e9u0rtvt8jrygyc8s,
  input   a02zzbowpjn06h,

  input   [2-1:0] r21i4by0bu3ks,

  output  tywculgjyor8ndw,


  output  tw5xnp59d8x,
  output  af5qc04tmn51e4u2h1z,

  output  qo5p9t6s74zxpo,

  output [11:0] k3cmpuswk7in0u4,


  input   h7fseh5_df0hbx,

  input   uc5qxb4d2b28ye5,
  output  o2qkf90r783,

  input   w2fpnf5fg1byp6,

  output  y_0q8d40rrzolo1y6,
  output  qwcb6hcmvfqmf032z,
  input   ao17frh5wnr0wddz3,
  input   woon4h3ivznl_qiu7i_9,
  input   [4-1:0] p25dd0cxz7nmi6w9ebukmr,
  output  [4-1:0] uvgy9al0j8prciqsh,
  output  f8pn1x6gurodpy04d3j1ihn,
  output  mmludd_fnt2yevok8a1a0,
  input   buwj9_8l8bwj80kkinq9p,

  input   apid0ys34zyekptw7un,
  output  um8zsjyxn_4p,  

  output av1w8ld09cfofn,
  output im2b5l0h98avl6t4sj,
  output bw65wl7fvekfymd8vqx,
  output [64-1:0] pecbpcoa04vq,
  output [64-1:0] tb_snaxyfs,
  output [64-1:0] zc4mldgm25r,
  output [32-1:0] d23wb5yh1iyvf,
  output [1:0] srim3bfnzhve,
  output fvqwdz2hdbb,
  output cy3nuhzm_v2p73mt,


  input  fcjh1nct4r,
  input  [9:0] b4lwcgm6l21pi,
  input  zwcbp7zqfei5xz,
  input  dn8riluj40uunvq5,
  output dz0zrf512290tvcy4q,
  input [64-1:0] z0yhjfv_e0yaa2r,
  output z1l80uwh6vyyg34,
  input  rn1o3sl83,

  input   x6eltyshbu5,
  input   lt3v_fm0ipu,
  input   v3ne7glf8d8,
  input   v9dnbgjy6c0vf,
  input   hmzw4exmjn8k921c,

  input   siifnhwgancn8,
  input   mfzl2fqml69hx,
  input   aw0hbwfkx3f63s,
  input   u83p4flbuvkqt26z,
  input   tvglhc8o_izdq,


  input   s5f_36xvqrtq7,

  input                      gkjb6c98b5j1zsgbv26,
  input                      unntlrmfpzgdq8rnz3ug3_8,
  input                      asxvrob6s2_85u99em22,
  input                      bva3_s2oj2hgomj0eyrk,
  input                      n9q1kib2q28tfyzyue2j2or,
  input [64-1:0]  fbgda1d6z8gr725snyc2ylc,

  input  [31:0] qqlnmd2zlr98m5mdjyk,
  output [31:0] xq63jpu81drai3h0,
  input                      q23hngbyy69cc9ci9sjr8g4,
  input [64-1:0]  vqv5qr4a5j6difuyllem3ur_,
  input                      rnodgdrxyr_tulm0nnnign,

  input                      s_qow7tm_gendxgd,
  input [64-1:0]  j_v6uy8_pdqb7w,    
  input [4-1:0]t3xakjcvvthgm_v0,    

  input                      tb198r6lzk1sr77g4,
  input [64-1:0]  cvvsn7xc8qg5uk,    
  input [4-1:0]pc67uztpd_zg6bsal,    

  input                      d3n7pwgwcgze9cr4,
  output                     cphtk1_x8fwehad,
  input  [64-1:0] amc4c8vcbecv1i,  
  input  [32-1:0] qgp6cehpls743wtn0i,  
  input                      ama4p78xalq9j32,
  input                      zcldu5wj7n47pd36vbj,  
  input  [64-1:0]    d0e2kztse3ur2dt22q,
  input                      y4fasvbsps__6yzpqc7eymh,
  input                      k_5q95o2gjo1w_rk,

  input                      f_4x5ty4man9f87i,
  input                      uzhgx8hpcw0vcm6nfex,
  input                      ichypldcqgx_6hsv, 
  input                      mn3xo91xnxw486688t,
  input                      omxbj0blxqsqi9h,
  input                      yhg7so3hz941h,
  input                      qa04tbszp_crup1y4rvk,
  input                      p38eaxsiobphopbri,
  input                      c4mm5jszl6uvumay,
  input                      npbrk566oq0dkbf982i,
  input                      wyutdg78_ykde5xhd,
  input                      jw67do539fm4kvlowut9k62,
  input                      gqwf5n54sp4jlral,
  input                      eo9f914sbhga72uw1z,
  input                      xi8b7jmwma99a4gxgmri9v74 ,
  input                      g0esgcmgdknyveiq2t72xopfk ,
  input                      o4512597_0nxc_jrf287w8it ,
  input                      l4km4217yp2p969cwda8 ,
  input                      ugimrlqwlbs5gblkxuymto1h4 ,
  input                      xktv6472l59a_iqmuyhu ,

  input                      p27tnvqrliur1xjlr527b,
  output                     rx_c151de4k7bbwnwrak,
  input                      k3t4av4o2bjnmmpxdoqfumyxecc09u7q5h,
  input                      n3tpm7ps0ygbm4a_yr6ryn06egc1 ,
  input                      bnta1_ctyuyz6f0cs2zpyuy2nmfjv4 ,
  input                      rgf8gwy5mb_doix8zdjh30tiklwj ,
  input                      khjs1qtt_oec9bu6269tck93yo8gpdw ,
  input                      k7nmctokgpx6dz4ugb1i3zr9q20f ,
  input                      awq_rxiss6jp46gvm3g,
  input                      rgsv1cqeh7x_1ex_5tj,

  input                      kdofxulgpcpa9q310, 
  input                      e9g0sper1c9v_vmf,
  input                      xv88qbq7hr0lskm4cqrn,
  input                      zjuaef59fqixf4nfbc , 
  input                      yy8cmh_xtnis7nqw_60 , 
  input                      t73hv26oh7wdnclcbf5b6j9 ,      
  input                      zi6t1yvku2qc168r2cv9b4v10vi6ee7 , 
  input [5-1:0] fuvqsp044l3a4fk69bkuvqopz0 , 
  input [64-1:0]     pji7j1gx57ht5kwknem7at7 , 
  input [64-1:0]o09mrpo1o2k6w4jsat2_o,
  input                      dxvoc8nirjgo0by0yoex4l01a7 ,
  input                      cqlsgy50_6bt6xavc02vpsg9p,
  input                      iby9hp5grzp4ouc82c61kxa  , 
  input                      mpp5ftr3blzju24mrjjk4nv, 

  input  v1vwaj41ljxavm9366uapnar1zrk5,

  input                      gkhcosyb6da4dfdhh3,
  input                      qgf355r7t8juyfmkx9g,
  input  [64-1:0]    troptfm3sc9gj8rb  ,
  input  [64-1:0]    d_4gaf_5w4wygi9  ,




  input   pydatzxqqi,


  output  [64-1:0] wtd_nuaeb_mpye,
  output  x7eg618xaszd4f21cl_g,
  output  [64-1:0] elth4vimq_j,
  output  jlud6jeuxe0espga,






  output  [64-1:0] xd66pm611ai1dg,
  output  r9uxubpl2h2alj1q,
  output  ftp0juzjm2b587cyw5,

  output  sf0uuehfhfa,
  output  hvy2cpsp75f3,
  output  k3z202os,

  output  z35xlcc6bt4,
  output  [64-1:0] ew08uu2kn2p9e11s,
  output  xv08lot3vi9dag4vs0,
  output  [64-1:0] mtc04rctrfyb,
  output  if5jz8qk0aqefy3v35o,

  input   c4ughu0qm5sfai,


  output  [64-1:0] qeb3z0x5,
  output  ibhfuwrztbm8p4gg,
  output  [3-1:0] i8_5wt0vppx,
  output  osv2437qj_3nuf,


  output  b7g_vsn0zoewh6g1,
  output  [2-1:0] onnv64ydiajl,



  input   c5ewdqztjw9za,
  input   rn2mt6nngsc9w5cz,

  input   t5trf35s8vy,
  input   zbac123pv78sbz3,

  input   z4e_m564fxae0kpbjr,
  input   hixy2y36a1pn0,
  input   ozwene1gdpatk6g,

  input  [64*4-1:0] azll7rq5fab5ou,
  input  [64*4-1:0] n6a0r_0zddzrme8,
  output ns0i7siujgkrghjpqv6,

  output                     rrujrlc85mhm,



  output                     jw4fsjecr0u919fr7,
  output                     s_m3pbf5m2tr6v,
  input [64-1:0]  bde41te346q515l,
  output                     gfod0nmy6eta29jeeg6mr2,
  output                     n4soswat5yihd74b,
  output                     y8wz7aud_fd6dfiakjtx2i0g,
  output                     dgnjyd9xs8efyxm0tdlsvfq4eop,
  output                     a3xib90kwk4_hm1,
  output                     nfzexr8q9g893gi,
  output [64-1:0] opkkwp3eg8g3448t,
  output                     tv3_4qrynvnaoy4riz,

  input [64-1:0]  pldoasxyzlvx2,


  input [64-1:0]  hn85hkp2yav,
  input [64-1:0]     unbt3q05xijb,
  input [64-1:0]     hawbmpz6j7pzibqr,


  input   o7hoht1pqz01v7,
  input   [64-1:0] kbv2bs_lxmvu,

  output [64-1:0] lovkp0eqfnxtb7,




  input   w632tcbtqncn6,
  input   ai169tbqp4seb3,
  input   b0zz_ornhz010,
  input   yw4o4kdms07_32,
  input   ezl3jzeqhltgj7h,
  input   w529wbj853,
  input   i9xvsmm45fp0f58,
  input   [64-1:0]     r4bs4k_53n5wp,


  input   jqsukc5b5drcc1e78,
  input   gnn46rd7vvofruqij,
  input   vkyge0q4mfc5,
  input   [64-1:0]     cppkd01vpwwnlfy,
  input   [64-1:0]  d3hccrck1fl7jjf6,
  input   [64-1:0]     h_qwsgi7nk2,

  output  [64-1:0]     u25pqekq4df,
  output                       dhjwho76fa8hqc,
  output  [64-1:0]     xel6gw173w5x0,
  output                       icauf4l_12_c2xkj53lf,
  output  [64-1:0]     v8ydjtlz16x9tx,
  output                       e_z6d7r9kxqg32te,
  output  [64-1:0]  p5jpgn4rvarpo,
  output                       z2g63deibg1b1quqr,
  output  [64-1:0]     tlgcdv86voe9,
  output                       u_ufp_wg29ieoklxxz1,



  input   um28jgd2x4mbs,

  input   aw82i964do,
  input   cwwkpmk260lrt,
  input   rvr30vvllni,
  input   z1cj655u31,
  input   y8_gkxsfle,
  input   lhu2z948o3n,

  output                     i32x_jtt7bvmr9lu2p,
  input                      mxa77etukhs8o_5z6962l19,
  input                      cd4v4c_rw906kt5,
  input                      idat72abxke4z9s,
  input                      hv4wuttuo9jk_cqa8sxqwt , 
  input [64-1:0]r_8f7p3tznijza5y03ko,
  input                      ac8_dky9fhpbsxu0b9t88ag8,









  output  v35y3qnk7mx3l1695,

  input   zsgl59ydqwjln,
  output  b9yq2alidby7zgom1,
  output  tvqijouldcgiz2dxdco7,  
  output  zkxlkidschdubxpkpm,  
  output  xmcrni1qngfvh9pil9j,  
  output  btkcf2uqr61gkiqhde0lai,  
  output  [64-1:0] h01d94xsxbxe_req,  
  output  w1casjl7bz73brz,  
  output  hjri7cufo9ckntq,  
  output  yghffofulqa77bd7aw07badta1a,
  output  rrl7evvmayt1_vvp74iq9h6_cjf,
  output  [27-1:0] zddoxp22m1o11x30gbe,
  output  [16-1:0] hwfethpzkuauejcgtbl6o,  

  input   n3ak8l6cvn0s4,
  output  hsxh9536ho4bw8o,
  output  r_edve7v9jcr26q6zk,  
  output  vrqfzuog2k4pos133,  
  output  bmw2yi333716crywk,  
  output  k2sr7sw1plcmnki5ajtscw,  
  output  [64-1:0] jkzw_f9anx55,  
  output  t8muv9e6d7yk_whqa0,  
  output  hzdfp71n6g3f5fsg5,  
  output  lwdhmuzyvcvv14mjbl0h2a41z,
  output  xy48dugh009wtmazqug3kpy2a5h_,
  output  [27-1:0] l4ztejmt2__wxqm2rw,
  output  [16-1:0] s3ujdp2a8n69bm6engxok,  

  input   bisaqpu86vneunhkqtg,
  input   m3ar1m0lklmpw4oek2yjd3ev,  
  input   zk19lxmoqrzcdjx6rxuvc36,  
  input   a5_uct872oszxvfp4kn_,  
  input   pl2up5ze0wczfdx0ga70d,  
  input   [64-1:0] jathu3ui07hzkaq4g2z39,  

  input   psx330qmvh5so1to4iq,
  input   sefocn4wjn2k2f_zvlvnz,  
  input   qknomh2kbth19r1osddvzly,  
  input   bzz8x0np0dpmdjt1d0w7uf,  
  input   rl9a96pgy3troiao05jel,  
  input   [64-1:0] hzsp_nydab9ghw59v,  

  input   xsekawjaoeqedkdymhz6h,
  input   vsrfdna3ksbt8a__05sjdxr,  
  input   uttwdi1xwyv_l7uzt3x2ea,  
  input   d14swmczjaws9gr8uvx,  
  input   fg6gtaxnx8a0anercx,  
  input   [64-1:0] b0cs5n_1_q64sumeg,  

  output  qk0jm7flfzap,
  output  [4-1:0] fj4fje1ckitqjb_7,    
  output  nes78rg61lk5t2,

  input  dk2xhkj77a,
  input  gf33atgy,
  input  ru_wi
  );


  wire ip4b_cj6h98z45oey8l;


  wire                      cj4f17jo0s_z9vmi5htht;
  wire                      a0itdy0a5fts62ldu_woafqynzc;  
  wire                      zn5lc4nu61e0ms4p0u4v2siuxjz_6;  
  wire                      r0nx0iuols_4pg0z96k6ifhert;  
  wire [64-1:0] ztfuyixi1aw62ttyksukyd;
  wire d3vybluuijhl4u65a3wsn_n6i1;
  wire y0nferrzezge90_qml8ypux7i;

  wire                      v_4emtojw2fdkpaawwtjk4l;


  wire glime27x19feqrvvsa2nmeh5f;
  wire oyiml9jn3w6vt88yja9asjx;

  lqqd_zj04p6o3_g6h1le u_ux607_exu_branchslv(
    .r21i4by0bu3ks                   (r21i4by0bu3ks),
    .ip4b_cj6h98z45oey8l           (ip4b_cj6h98z45oey8l),
    .w5rbttl5mj11z                 (v_4emtojw2fdkpaawwtjk4l    ),
    .lu3guz5hxinmv_i4vg2k             (q23hngbyy69cc9ci9sjr8g4   ),  
    .tbncz5fmqkrrvgqd9n8lz        (vqv5qr4a5j6difuyllem3ur_),
    .m5qoggt2in4ie_llz91            (rnodgdrxyr_tulm0nnnign),

    .d2cosjdh8e6u1zldf6kf09           (p27tnvqrliur1xjlr527b),
    .l9wonwtwviy4i8w6s            (rx_c151de4k7bbwnwrak),
    .nwpj2xvetia76ai6nkrnv5k8cpxq   (k3t4av4o2bjnmmpxdoqfumyxecc09u7q5h),
    .xlzi1qrfl8ef8u0                  (k_5q95o2gjo1w_rk    ),  
    .uiqmdx8tnsb                   (f_4x5ty4man9f87i     ),  
    .c9q9b8x3r05mpe5                  (uzhgx8hpcw0vcm6nfex    ),  
    .ntedv1bjeakd                   (ichypldcqgx_6hsv     ),  
    .i1a3ajcrp                   (mn3xo91xnxw486688t     ),  
    .wokc20mug9u1gn                  (omxbj0blxqsqi9h    ),  
    .asl4zsbrnfn7                (qa04tbszp_crup1y4rvk  ),
    .psf3mvojppotcy                (p38eaxsiobphopbri  ),
    .yec_1lu2ooyq                  (c4mm5jszl6uvumay     ),
    .bn3gk8oaq6g3ax                  (npbrk566oq0dkbf982i     ),
    .hhimu5qv7me_z              (wyutdg78_ykde5xhd     ),
    .obqt4l21562rgtgxh              (jw67do539fm4kvlowut9k62),
    .otv3n61fdzkg6gt              (awq_rxiss6jp46gvm3g),
    .bq_u11fb64d2bir3vxj              (rgsv1cqeh7x_1ex_5tj),
    .sfs34sstg9pk                    (amc4c8vcbecv1i      ),
    .c_fnucn4hvf3g               (d0e2kztse3ur2dt22q),


    .l7r_xp04shn9v4n12        (g0esgcmgdknyveiq2t72xopfk    ),
    .ouj04k7brubwkv_h9qhnkh    (v1vwaj41ljxavm9366uapnar1zrk5),
    .c00vdqa8yvwhd6r55g      (ugimrlqwlbs5gblkxuymto1h4  ),
    .lovkp0eqfnxtb7            (lovkp0eqfnxtb7            ),

    .rrujrlc85mhm            (rrujrlc85mhm                  ),



    .jw4fsjecr0u919fr7            (jw4fsjecr0u919fr7                   ),
    .gfod0nmy6eta29jeeg6mr2      (gfod0nmy6eta29jeeg6mr2),
    .n4soswat5yihd74b         (n4soswat5yihd74b),
    .y8wz7aud_fd6dfiakjtx2i0g   (y8wz7aud_fd6dfiakjtx2i0g),  
    .a3xib90kwk4_hm1         (a3xib90kwk4_hm1),
    .nfzexr8q9g893gi          (nfzexr8q9g893gi),
    .opkkwp3eg8g3448t         (opkkwp3eg8g3448t),
    .pldoasxyzlvx2              (pldoasxyzlvx2         ),


    .hn85hkp2yav               (hn85hkp2yav         ),
    .s_m3pbf5m2tr6v            (s_m3pbf5m2tr6v      ),
    .bde41te346q515l              (bde41te346q515l        ),
    .tv3_4qrynvnaoy4riz           (tv3_4qrynvnaoy4riz     ),

    .pydatzxqqi                (pydatzxqqi),
    .aw82i964do                  (aw82i964do),
    .rvr30vvllni              (rvr30vvllni),
    .z1cj655u31              (z1cj655u31),
    .y8_gkxsfle                  (y8_gkxsfle),
    .lhu2z948o3n              (lhu2z948o3n),

    .glime27x19feqrvvsa2nmeh5f(glime27x19feqrvvsa2nmeh5f),
    .llyh4o81vzcbw0zjekct       (1'b1    ),
    .mnqkmoietusiwyf95g       (cj4f17jo0s_z9vmi5htht    ),


    .bq75f6k903dwxcstjv1wpw2cg09  (a0itdy0a5fts62ldu_woafqynzc),  
    .m1yqe0cmaq2_frcfgf_1c1qtgm7  (zn5lc4nu61e0ms4p0u4v2siuxjz_6),  
    .t2uejj01ae4b5d7shv4q2x  (r0nx0iuols_4pg0z96k6ifhert),  
    .sdsekm12iz4x32pwrh        (ztfuyixi1aw62ttyksukyd),  
    .tskef3o28v1jcu97th07m_    (d3vybluuijhl4u65a3wsn_n6i1),
    .nd7mxlwd9xekhy2oqb88dre5    (y0nferrzezge90_qml8ypux7i),

    .gf33atgy   (gf33atgy  ),
    .ru_wi (ru_wi)
  );

  wire ljd_sv9l5ykkrwitvxjydqd5n55;  
  wire wrg2t13vafz_5z44ejdmrpmnk1;  
  wire g7cxea_49xi94dndcklkkq;  
  wire vj6p6j6avq664060js8d_wit_7a;  


  wire [64-1:0] vfga_wjq02bdlelajwej;
  wire n8337lh9w_n6vby0gecd6esky;

  wire fh49u69v0he;


  qaszx6xv9r9g8927s  u_ux607_exu_excp(
    .a02zzbowpjn06h   (a02zzbowpjn06h),

    .se2buoxmq91dbic3y2m5hu (se2buoxmq91dbic3y2m5hu),
    .e9u0rtvt8jrygyc8s     (e9u0rtvt8jrygyc8s),

    .feq1g7m2cy1erl     (feq1g7m2cy1erl),

    .av1w8ld09cfofn     (av1w8ld09cfofn    ),
    .im2b5l0h98avl6t4sj (im2b5l0h98avl6t4sj),
    .bw65wl7fvekfymd8vqx  (bw65wl7fvekfymd8vqx ),
    .pecbpcoa04vq      (pecbpcoa04vq     ),
    .tb_snaxyfs       (tb_snaxyfs      ),
    .zc4mldgm25r      (zc4mldgm25r     ),
    .d23wb5yh1iyvf      (d23wb5yh1iyvf     ),
    .srim3bfnzhve       (srim3bfnzhve      ),
    .fvqwdz2hdbb      (fvqwdz2hdbb     ),
    .cy3nuhzm_v2p73mt  (cy3nuhzm_v2p73mt ),  

    .rvr30vvllni              (rvr30vvllni),

    .k3cmpuswk7in0u4   (k3cmpuswk7in0u4),
    .btwmhh91h50d5flgwx4o6pwu (btwmhh91h50d5flgwx4o6pwu),
    .tywculgjyor8ndw (tywculgjyor8ndw),







    .h7fseh5_df0hbx         (h7fseh5_df0hbx),

    .uc5qxb4d2b28ye5          (uc5qxb4d2b28ye5),
    .o2qkf90r783          (o2qkf90r783),





    .w2fpnf5fg1byp6      (w2fpnf5fg1byp6),


    .tw5xnp59d8x              (tw5xnp59d8x        ),
    .y_0q8d40rrzolo1y6      (y_0q8d40rrzolo1y6),
    .qwcb6hcmvfqmf032z      (qwcb6hcmvfqmf032z),
    .ao17frh5wnr0wddz3      (ao17frh5wnr0wddz3),
    .woon4h3ivznl_qiu7i_9      (woon4h3ivznl_qiu7i_9),
    .p25dd0cxz7nmi6w9ebukmr     (p25dd0cxz7nmi6w9ebukmr),
    .uvgy9al0j8prciqsh        (uvgy9al0j8prciqsh   ),
    .f8pn1x6gurodpy04d3j1ihn     (f8pn1x6gurodpy04d3j1ihn   ),
    .mmludd_fnt2yevok8a1a0      (mmludd_fnt2yevok8a1a0),
    .buwj9_8l8bwj80kkinq9p      (buwj9_8l8bwj80kkinq9p),
    .apid0ys34zyekptw7un       (apid0ys34zyekptw7un),
    .um8zsjyxn_4p             (um8zsjyxn_4p      ),  

    .wtd_nuaeb_mpye           (wtd_nuaeb_mpye    ), 
    .x7eg618xaszd4f21cl_g       (x7eg618xaszd4f21cl_g),
    .elth4vimq_j              (elth4vimq_j        ),
    .jlud6jeuxe0espga          (jlud6jeuxe0espga    ),
    .pldoasxyzlvx2           (pldoasxyzlvx2),
    .bde41te346q515l           (bde41te346q515l),






    .xd66pm611ai1dg             (xd66pm611ai1dg      ),
    .r9uxubpl2h2alj1q         (r9uxubpl2h2alj1q  ),

    .sf0uuehfhfa              (sf0uuehfhfa       ),
    .hvy2cpsp75f3               (hvy2cpsp75f3        ),
    .k3z202os              (k3z202os       ),
    .z35xlcc6bt4               (z35xlcc6bt4        ),
    .ew08uu2kn2p9e11s           (ew08uu2kn2p9e11s    ),
    .xv08lot3vi9dag4vs0       (xv08lot3vi9dag4vs0),
    .mtc04rctrfyb          (mtc04rctrfyb    ),
    .if5jz8qk0aqefy3v35o      (if5jz8qk0aqefy3v35o),


    .jw4fsjecr0u919fr7          (jw4fsjecr0u919fr7   ),
    .fh49u69v0he               (fh49u69v0he        ),
    .af5qc04tmn51e4u2h1z      (af5qc04tmn51e4u2h1z),

    .w632tcbtqncn6         (w632tcbtqncn6    ),
    .ai169tbqp4seb3            (ai169tbqp4seb3       ),
    .b0zz_ornhz010            (b0zz_ornhz010       ),
    .yw4o4kdms07_32            (yw4o4kdms07_32       ),
    .ezl3jzeqhltgj7h            (ezl3jzeqhltgj7h       ),
    .w529wbj853            (w529wbj853       ),
    .i9xvsmm45fp0f58            (i9xvsmm45fp0f58       ),
    .r4bs4k_53n5wp         (r4bs4k_53n5wp    ),
    .jqsukc5b5drcc1e78        (jqsukc5b5drcc1e78   ),
    .gnn46rd7vvofruqij        (gnn46rd7vvofruqij   ),
    .vkyge0q4mfc5          (vkyge0q4mfc5     ),
    .cppkd01vpwwnlfy           (cppkd01vpwwnlfy      ),
    .d3hccrck1fl7jjf6          (d3hccrck1fl7jjf6     ),
    .h_qwsgi7nk2           (h_qwsgi7nk2      ),
    .u25pqekq4df            (u25pqekq4df       ),
    .dhjwho76fa8hqc        (dhjwho76fa8hqc   ),
    .xel6gw173w5x0           (xel6gw173w5x0      ),
    .icauf4l_12_c2xkj53lf       (icauf4l_12_c2xkj53lf  ),
    .v8ydjtlz16x9tx          (v8ydjtlz16x9tx     ),
    .e_z6d7r9kxqg32te      (e_z6d7r9kxqg32te ),
    .p5jpgn4rvarpo              (p5jpgn4rvarpo         ),
    .z2g63deibg1b1quqr          (z2g63deibg1b1quqr     ),
    .tlgcdv86voe9          (tlgcdv86voe9     ),
    .u_ufp_wg29ieoklxxz1      (u_ufp_wg29ieoklxxz1 ),

    .p7rj2v1hvh0nab6ei      (d3n7pwgwcgze9cr4  ),
    .c8w01x5rfmr6shqzb      (n8337lh9w_n6vby0gecd6esky    ),
    .u3qmzjrm6inkod3m3ghp    (kdofxulgpcpa9q310),
    .fe8u85vitwnfnuszhl         (e9g0sper1c9v_vmf     ),
    .stx6pefjqd_oqqg5gej9      (xv88qbq7hr0lskm4cqrn  ),
    .qsn_nfmbj97wz1r3s59t2     (zjuaef59fqixf4nfbc ),
    .uuvo0ter1b1y6j1xfc     (yy8cmh_xtnis7nqw_60 ),
    .hjysp7ahvean99t41k89pt    (t73hv26oh7wdnclcbf5b6j9),
    .ggvuzlnuknlvg4a50n4hy7ok(zi6t1yvku2qc168r2cv9b4v10vi6ee7),
    .frfbo512g1_94ncrem_be859f  (fuvqsp044l3a4fk69bkuvqopz0),
    .lt3biawnyshgr5rw4q5chcg6u7rc(pji7j1gx57ht5kwknem7at7),
    .wql66zm9cb_1pzbk         (amc4c8vcbecv1i     ),
    .skcwu9hiw7zl59wu      (qgp6cehpls743wtn0i  ),
    .ij7ql6t124xbofcx      (ama4p78xalq9j32  ),
    .fof2qu1zf51j1nid7vs4       (k_5q95o2gjo1w_rk   ),
    .umg0x8yb1yqjkaw34l6t     (zcldu5wj7n47pd36vbj ),
    .z2574r4ajgr7u7mtpb_wpetx  (y4fasvbsps__6yzpqc7eymh),
    .k84xk2u4clez          (j_v6uy8_pdqb7w     ),
    .jd2_q1xken6mnd8v      (s_qow7tm_gendxgd ),
    .tb198r6lzk1sr77g4      (tb198r6lzk1sr77g4 ), 
    .cvvsn7xc8qg5uk          (cvvsn7xc8qg5uk     ), 
    .jp82o1hu0f41an        (zcldu5wj7n47pd36vbj ), 
    .n7orghfl8x_7wsaisuhpw9o    (o09mrpo1o2k6w4jsat2_o ),
    .j6g8r7rblr88am07jc3i5      (gqwf5n54sp4jlral   ),
    .klz7l8_75czqn63zb     (eo9f914sbhga72uw1z  ),
    .esb6gep_3iit0w        (yhg7so3hz941h  ),
    .iq2e_b4p5qjp2ryy5sktbl6kd0(xi8b7jmwma99a4gxgmri9v74),
    .om206h86cfrb69iqc9pzq3fq1 (g0esgcmgdknyveiq2t72xopfk ),
    .yk85cwkls6hcvp4_g70j2 (o4512597_0nxc_jrf287w8it ),
    .cj2z8_7e4hw2s1u6mhckmpm4i (l4km4217yp2p969cwda8 ),
    .rpt826mhm0kwty9qlty6rt1  (xktv6472l59a_iqmuyhu  ),
    .pmcsf3olv_ztinoakqw67nno42plkv(n3tpm7ps0ygbm4a_yr6ryn06egc1),
    .dgigaix0xkzcg64kbmiqjlagh1cqid2(bnta1_ctyuyz6f0cs2zpyuy2nmfjv4),
    .m2av7b78yjzgy1j3a9inerkjyzrkdg9  (rgf8gwy5mb_doix8zdjh30tiklwj  ),
    .z2tyajok7rez0sc5ugh28p8o0rsrq  (khjs1qtt_oec9bu6269tck93yo8gpdw  ),
    .o2rr0tomxjme9ua4btx71i4hsfz  (k7nmctokgpx6dz4ugb1i3zr9q20f  ),
    .wkyo2nrlaz9sq3m1chcysnofuenz  (dxvoc8nirjgo0by0yoex4l01a7  ),
    .vmkmkz3cm8cgbet959d4pw_0ti(cqlsgy50_6bt6xavc02vpsg9p),
    .gnn94t_31a_j59f483ym5f68sb    (iby9hp5grzp4ouc82c61kxa  ),     
    .zb322_7v29pmo4jvmvow3qi8  (mpp5ftr3blzju24mrjjk4nv),

    .lovkp0eqfnxtb7            (lovkp0eqfnxtb7            ),

    .fi9wz0kme0ey_bxavdqx_9      (gkjb6c98b5j1zsgbv26),
    .tmhbzyv2b510vt_9qkb16hdwa   (unntlrmfpzgdq8rnz3ug3_8),
    .nqoqg40hg82wgdbsfubvu4fg  (asxvrob6s2_85u99em22),
    .hcx0jkab_j87_6j7phxnsz  (bva3_s2oj2hgomj0eyrk),
    .t0zuyah73tpfg_dtxy56ug9ej  (n9q1kib2q28tfyzyue2j2or),
    .sq0y2gv0vwpq_6ckk9b89gybz (fbgda1d6z8gr725snyc2ylc),

    .i32x_jtt7bvmr9lu2p    (i32x_jtt7bvmr9lu2p  ),
    .mxa77etukhs8o_5z6962l19    (mxa77etukhs8o_5z6962l19  ),
    .cd4v4c_rw906kt5       (cd4v4c_rw906kt5     ),
    .idat72abxke4z9s       (idat72abxke4z9s     ),
    .hv4wuttuo9jk_cqa8sxqwt   (hv4wuttuo9jk_cqa8sxqwt ),
    .ac8_dky9fhpbsxu0b9t88ag8   (ac8_dky9fhpbsxu0b9t88ag8 ),
    .r_8f7p3tznijza5y03ko  (r_8f7p3tznijza5y03ko),

    .unbt3q05xijb           (unbt3q05xijb       ),

    .hawbmpz6j7pzibqr           (hawbmpz6j7pzibqr       ),

    .o7hoht1pqz01v7          (o7hoht1pqz01v7),
    .kbv2bs_lxmvu           (kbv2bs_lxmvu ),

    .fcjh1nct4r(fcjh1nct4r),
    .b4lwcgm6l21pi(b4lwcgm6l21pi),
    .zwcbp7zqfei5xz(zwcbp7zqfei5xz),
    .dn8riluj40uunvq5(dn8riluj40uunvq5),
    .dz0zrf512290tvcy4q(dz0zrf512290tvcy4q),
    .z0yhjfv_e0yaa2r(z0yhjfv_e0yaa2r),

    .z1l80uwh6vyyg34         (z1l80uwh6vyyg34),
    .rn1o3sl83             (rn1o3sl83),


    .x6eltyshbu5            (x6eltyshbu5        ),
    .lt3v_fm0ipu            (lt3v_fm0ipu        ),
    .v3ne7glf8d8            (v3ne7glf8d8        ),
    .v9dnbgjy6c0vf          (v9dnbgjy6c0vf      ),
    .hmzw4exmjn8k921c           (hmzw4exmjn8k921c       ),

    .siifnhwgancn8            (siifnhwgancn8        ),
    .mfzl2fqml69hx            (mfzl2fqml69hx        ),
    .aw0hbwfkx3f63s            (aw0hbwfkx3f63s        ),
    .u83p4flbuvkqt26z          (u83p4flbuvkqt26z      ),
    .tvglhc8o_izdq           (tvglhc8o_izdq       ),

    .s5f_36xvqrtq7          (s5f_36xvqrtq7),

    .c4ughu0qm5sfai          (c4ughu0qm5sfai),

    .qeb3z0x5               (qeb3z0x5        ),
    .ibhfuwrztbm8p4gg           (ibhfuwrztbm8p4gg    ),
    .i8_5wt0vppx            (i8_5wt0vppx     ),
    .osv2437qj_3nuf        (osv2437qj_3nuf ),


    .b7g_vsn0zoewh6g1          (b7g_vsn0zoewh6g1),
    .onnv64ydiajl              (onnv64ydiajl    ),

    .c5ewdqztjw9za              (c5ewdqztjw9za),
    .rn2mt6nngsc9w5cz      (rn2mt6nngsc9w5cz),

    .azll7rq5fab5ou      (azll7rq5fab5ou      ),
    .n6a0r_0zddzrme8      (n6a0r_0zddzrme8      ),
    .ns0i7siujgkrghjpqv6(ns0i7siujgkrghjpqv6),

    .t5trf35s8vy            (t5trf35s8vy),
    .zbac123pv78sbz3         (zbac123pv78sbz3),
    .z4e_m564fxae0kpbjr         (z4e_m564fxae0kpbjr),
    .hixy2y36a1pn0         (hixy2y36a1pn0),
    .ozwene1gdpatk6g            (ozwene1gdpatk6g),

    .pydatzxqqi              (pydatzxqqi),

    .um28jgd2x4mbs            (um28jgd2x4mbs),

    .aw82i964do                (aw82i964do),
    .y8_gkxsfle                (y8_gkxsfle),
    .cwwkpmk260lrt                (cwwkpmk260lrt),


    .ip4b_cj6h98z45oey8l        (ip4b_cj6h98z45oey8l       ),
    .ljd_sv9l5ykkrwitvxjydqd5n55   (ljd_sv9l5ykkrwitvxjydqd5n55),
    .wrg2t13vafz_5z44ejdmrpmnk1   (wrg2t13vafz_5z44ejdmrpmnk1),
    .g7cxea_49xi94dndcklkkq   (g7cxea_49xi94dndcklkkq),
    .vj6p6j6avq664060js8d_wit_7a   (vj6p6j6avq664060js8d_wit_7a),
    .vfga_wjq02bdlelajwej         (vfga_wjq02bdlelajwej),

    .glime27x19feqrvvsa2nmeh5f(glime27x19feqrvvsa2nmeh5f),
    .oyiml9jn3w6vt88yja9asjx   (oyiml9jn3w6vt88yja9asjx),

    .qo5p9t6s74zxpo (qo5p9t6s74zxpo),

    .dk2xhkj77a (dk2xhkj77a),
    .gf33atgy   (gf33atgy  ),
    .ru_wi (ru_wi)
  );





  wire hgx15j0zue2pefkufzq = b9yq2alidby7zgom1 | hsxh9536ho4bw8o;
  assign dgnjyd9xs8efyxm0tdlsvfq4eop = hgx15j0zue2pefkufzq; 

  assign cphtk1_x8fwehad = n8337lh9w_n6vby0gecd6esky & v_4emtojw2fdkpaawwtjk4l;


  wire ye5_uo_8dtdw3, pl_2g1e8267skhkk; 
  wire tcul30o723hqzs8i, l4mlt7so_hfc82en;

  wire [4-1:0] hno_lpz_7d804vv;
  wire [4-1:0] pw5op4ktw7ff093ctpjt6 = oyiml9jn3w6vt88yja9asjx ? pc67uztpd_zg6bsal : (qwcb6hcmvfqmf032z ? pc67uztpd_zg6bsal : t3xakjcvvthgm_v0);

  assign b9yq2alidby7zgom1      = 1'b0;
  assign tvqijouldcgiz2dxdco7 = 1'b0;
  assign zkxlkidschdubxpkpm = 1'b0;
  assign xmcrni1qngfvh9pil9j = 1'b0;
  assign btkcf2uqr61gkiqhde0lai = 1'b0;
  assign h01d94xsxbxe_req       = 64'b0;
  assign w1casjl7bz73brz   = 1'b0;
  assign hjri7cufo9ckntq           = 1'b0;
  assign yghffofulqa77bd7aw07badta1a    = 1'b0;
  assign rrl7evvmayt1_vvp74iq9h6_cjf  = 1'b0;
  assign zddoxp22m1o11x30gbe        = {27{1'b0}};
  assign hwfethpzkuauejcgtbl6o      = 16'b0;
  assign tcul30o723hqzs8i = 1'b0;
  assign ye5_uo_8dtdw3     = 1'b0;
  
  
  assign hsxh9536ho4bw8o     = bisaqpu86vneunhkqtg | psx330qmvh5so1to4iq | xsekawjaoeqedkdymhz6h | ip4b_cj6h98z45oey8l | cj4f17jo0s_z9vmi5htht;
  assign l4mlt7so_hfc82en = (bisaqpu86vneunhkqtg | psx330qmvh5so1to4iq) | (cj4f17jo0s_z9vmi5htht & (uzhgx8hpcw0vcm6nfex | ichypldcqgx_6hsv));
  assign pl_2g1e8267skhkk    = hsxh9536ho4bw8o & (~(l4mlt7so_hfc82en));

  
     
  assign r_edve7v9jcr26q6zk = bisaqpu86vneunhkqtg ? m3ar1m0lklmpw4oek2yjd3ev : psx330qmvh5so1to4iq ? sefocn4wjn2k2f_zvlvnz : xsekawjaoeqedkdymhz6h ? vsrfdna3ksbt8a__05sjdxr : ip4b_cj6h98z45oey8l ? ljd_sv9l5ykkrwitvxjydqd5n55 : a0itdy0a5fts62ldu_woafqynzc;   
  assign vrqfzuog2k4pos133 = bisaqpu86vneunhkqtg ? zk19lxmoqrzcdjx6rxuvc36 : psx330qmvh5so1to4iq ? qknomh2kbth19r1osddvzly : xsekawjaoeqedkdymhz6h ? uttwdi1xwyv_l7uzt3x2ea : ip4b_cj6h98z45oey8l ? wrg2t13vafz_5z44ejdmrpmnk1 : zn5lc4nu61e0ms4p0u4v2siuxjz_6;   
  assign bmw2yi333716crywk = bisaqpu86vneunhkqtg ? a5_uct872oszxvfp4kn_ : psx330qmvh5so1to4iq ? bzz8x0np0dpmdjt1d0w7uf : xsekawjaoeqedkdymhz6h ? d14swmczjaws9gr8uvx : ip4b_cj6h98z45oey8l ? g7cxea_49xi94dndcklkkq : r0nx0iuols_4pg0z96k6ifhert;   
  assign k2sr7sw1plcmnki5ajtscw = bisaqpu86vneunhkqtg ? pl2up5ze0wczfdx0ga70d : psx330qmvh5so1to4iq ? rl9a96pgy3troiao05jel : xsekawjaoeqedkdymhz6h ? fg6gtaxnx8a0anercx : ip4b_cj6h98z45oey8l ? vj6p6j6avq664060js8d_wit_7a : 1'b0;                         
  assign jkzw_f9anx55       = bisaqpu86vneunhkqtg ? jathu3ui07hzkaq4g2z39    : psx330qmvh5so1to4iq ? hzsp_nydab9ghw59v    : xsekawjaoeqedkdymhz6h ? b0cs5n_1_q64sumeg    : ip4b_cj6h98z45oey8l ? vfga_wjq02bdlelajwej       : ztfuyixi1aw62ttyksukyd;         
  assign t8muv9e6d7yk_whqa0   = bisaqpu86vneunhkqtg ? 1'b0                : psx330qmvh5so1to4iq ? 1'b0                : xsekawjaoeqedkdymhz6h ? 1'b0               : ip4b_cj6h98z45oey8l ? 1'b0                   : d3vybluuijhl4u65a3wsn_n6i1;     
  assign hzdfp71n6g3f5fsg5   = bisaqpu86vneunhkqtg ? 1'b0                : psx330qmvh5so1to4iq ? 1'b0                : xsekawjaoeqedkdymhz6h ? 1'b0               : ip4b_cj6h98z45oey8l ? 1'b0                   : y0nferrzezge90_qml8ypux7i;     
  assign lwdhmuzyvcvv14mjbl0h2a41z    = ~gkhcosyb6da4dfdhh3 & y0nferrzezge90_qml8ypux7i;
  assign xy48dugh009wtmazqug3kpy2a5h_  = ~qgf355r7t8juyfmkx9g & y0nferrzezge90_qml8ypux7i;
  assign l4ztejmt2__wxqm2rw        = gkhcosyb6da4dfdhh3 ? {27{1'b0}} : ({27{y0nferrzezge90_qml8ypux7i}} & troptfm3sc9gj8rb[27+12-1:12]);
  assign s3ujdp2a8n69bm6engxok      = qgf355r7t8juyfmkx9g ? {16{1'b0}}    : ({16{y0nferrzezge90_qml8ypux7i}}    & d_4gaf_5w4wygi9[16-1:0]);
  assign hno_lpz_7d804vv     = bisaqpu86vneunhkqtg ? pc67uztpd_zg6bsal      : psx330qmvh5so1to4iq ? pc67uztpd_zg6bsal      : xsekawjaoeqedkdymhz6h ? pc67uztpd_zg6bsal     : ip4b_cj6h98z45oey8l ? pw5op4ktw7ff093ctpjt6     : pc67uztpd_zg6bsal;         


  assign fh49u69v0he = d3n7pwgwcgze9cr4 & cphtk1_x8fwehad;



  assign ftp0juzjm2b587cyw5 = fh49u69v0he;



  assign af5qc04tmn51e4u2h1z = fh49u69v0he & (~hgx15j0zue2pefkufzq);



  assign v35y3qnk7mx3l1695 = glime27x19feqrvvsa2nmeh5f;







  assign xq63jpu81drai3h0[0] = 1'b0;

  assign xq63jpu81drai3h0[1] = 1'b1;







  assign xq63jpu81drai3h0[8:2] =  qqlnmd2zlr98m5mdjyk[8:2] & {7{ftp0juzjm2b587cyw5}};

  assign xq63jpu81drai3h0[9] = qqlnmd2zlr98m5mdjyk[9] & ftp0juzjm2b587cyw5 & rgsv1cqeh7x_1ex_5tj;
























  assign xq63jpu81drai3h0[31:10] = qqlnmd2zlr98m5mdjyk[31:10] & {22{ftp0juzjm2b587cyw5}};

  assign qk0jm7flfzap = hgx15j0zue2pefkufzq ; 

  assign fj4fje1ckitqjb_7 = hsxh9536ho4bw8o ? hno_lpz_7d804vv : pc67uztpd_zg6bsal; 
  assign nes78rg61lk5t2 = ye5_uo_8dtdw3 | pl_2g1e8267skhkk  ; 





endmodule                                      






















module nrcp90w_wy4yo (
  output pby60vfdze02,
  output [64-1:0] vm3pyzc9nt95,
  output rbz4pv_atxqopdwt,
  output [64-1:0] qs1xgat7r8xow,

  input  [64-1:0] lovkp0eqfnxtb7,

  input vdr9fi9zwq,

  output exltui35irvvmodu205vw,
  output s7eq8f6z1uyi2in,
  output qbsr1jytrqtsbk4ttb8nz,
  output w92a5o09fp9dg6   ,
  output eglor15f7p2ivpny5dc   ,
  output ous_emkpecrqhg5e7,
  output doh50j3p7c7yl7uk9,
  output bisaqpu86vneunhkqtg,
  output m3ar1m0lklmpw4oek2yjd3ev,  
  output zk19lxmoqrzcdjx6rxuvc36,  
  output a5_uct872oszxvfp4kn_,  
  output pl2up5ze0wczfdx0ga70d,  
  output [64-1:0] jathu3ui07hzkaq4g2z39,  

  output xsekawjaoeqedkdymhz6h,
  output vsrfdna3ksbt8a__05sjdxr,  
  output uttwdi1xwyv_l7uzt3x2ea,  
  output d14swmczjaws9gr8uvx,  
  output fg6gtaxnx8a0anercx,  
  output [64-1:0] b0cs5n_1_q64sumeg,  

  output w2fpnf5fg1byp6,
  output x_cq40qmp6a, 

  input [12-1:0] k3cmpuswk7in0u4,  

  input [64-1:0] nchi0_6mu,  

  input  [64-1:0] wd9dvepxj,

  input xx87vzbpchg,
  input pvfk1_6o89lmby,
  input zz5wo47gw146x4,
  input fgr486jx5kevbua,

  output habgbg2jn3qi,
  output apid0ys34zyekptw7un,
  output dg4hzu_,
  output h7fseh5_df0hbx,
  input wj5ypo5k,

  output o7hoht1pqz01v7,
  output [64-1:0] kbv2bs_lxmvu,


                   
                   
                   
                   
                   
                   
  output [8*32-1:0] pcr4upio7_tx37, 
  output [8*1-1:0] uzklqlncpqqm1rav,
  output [8*1-1:0] ortueunvnkx_l5m_j,
  output [8*1-1:0] hwuhtb7ucto_utk56,
  output [8*2-1:0] i1env2kmns7qvvuuc,
  output [8*1-1:0] g3s3vpafvy3i,


  input [31:0] xq63jpu81drai3h0,

  output       rm1dxjejhq7dh3q5m,




  input af5qc04tmn51e4u2h1z,

  input [64-1:0] guuvp01vkcryglsu1p3,
  output ix299qulxi5, 
  output jjj61w03m77lv,
  input enwn0u48p2_ls5az80,
  output[64-1:0]     z0yhjfv_e0yaa2r,
  output [7:0] f_i1959b4xizzq9jea,
  input [9:0] b4lwcgm6l21pi,
  input [7:0] hjrk_rwjkqj3zk_b,
  input zwcbp7zqfei5xz,
  input znzjygllppv1s0a8cqub3c, 
  output gfy3zost37aq8qmr,
  output dxi_ue3gf5zqqqxwgq2a,
  output dn8riluj40uunvq5,
  input [4:0] ciw6wwc7i33adp5,
  input       elspwgn4qhqqwg31epb,
  output [2:0] phk590vi2,
  output rnx27onf2lbe,
  input  ya8t4ev_aidf0t0x4or,
  input rb050tnl,
  input a94vd35etec4,
  input el7_p8jit09,
  input [12-1:0] e1go3iu,

  output x8rpm78rvvycis,
  input bwbmafs1inesgjyn,
  output [74-1:0] canacnkc7zibtkn418i, 
  input bkkiffh6ob85nh79doya_,
  input  [5:0] qhqqh0lyehgtfop1tc, 
  output [74-1:0] x03ux1utw4qem5kk3c, 
  output sxhicsqvufwfbnk0,
  input ydydp69z03wvr97,
  input pjic5x84bqxpvdduy4r2s,
  input w5az87bw32r0tjbo0tdrv2ouvx,  

  
  
  output                                   vs6ryzcr0bwqs5so, 
  output [32-1:0]                  j25ub196dc_agl8oovaex4, 
  output                                   pi2nokcm8qf7och7l4g, 
  output                                   c0i0hs5tz64_ce5f0z, 
  output                                   dmzdczrqcueolg3dzufj_by5rmf, 
  output                                   a1sqko6fok9qzpbtyuw0, 
  output                                   bquohubxiv2rsayn62v, 
  input                                    kqyojh1maxy0x834htg, 


  output                                   hpk3eafyque5ubt_c62flnny,       
  output [27-1:0]      sfezv1xz2ghvo8pkt,               
  output [1:0]                             vagaza053272juvmo59v8w20s,       
  output                                   rzf45534z36ejq96260,                        
  output [26-1:0]    frzfsbt7hp3n4aj3zvvumnh0s,         
  output [64-1:0]                  zkuxqezrmlhyyjjgx,              
  output [64-1:0]                  u3h5tvu1g2q93141j9o,              
  output                                   pjh0wad7t_5du3cync_0c,                        
  output                                   wmkgrgf631pbq,
  input                                    oyq1p3qa2iffjuqns0jkgg,

  input                                    qjw2q0j88rjr42lautsqnca,       
  input [26-1:0]     imkm56ujne9v4m6n08w1yf5622,     
  input [20-1:0]          txk1r9aiq_7l2nkw101w_,          
  input                                    ih4hmwugasiodbx5da9_40kx,        
  input                                    x5vjq7mshfwr0h3q514t7mhdt,        
  input                                    qrxtk7e03100_uwkx73sg7,        
  input                                    i7qiq2q9c6hbeful9qu9lb,         
  input                                    yr0s3skqk7cdqflsrbsxg9znu,         
  input                                    adqieke11qo0elfz93hlouwjc0,   
  input                                    w93gdpnnxuydy53eu0s9nxw7xdct7, 

  
  output                           cn8o3075eju6dycby, 
  output                           zi39s8s7rmgo_lyocr_, 
  output [5-1:0]g1cek93tezrlyyt, 
  output [64-1:0]          i22z6k7eo0it77lz2, 
  output                           ldj4m511gvpu12mdu1_, 
  output                           sl5f3k5g9ln8_zvzr, 
  input                            w2h8uh3l463qbgqmv, 











  output r0s7d8cr68i2qs1z,
  output kakelc68be0x7tdm9b9o,
  output j3j1czgoam48vhs8auo,
  output gm1r5itc44uxw_y0_msk,

  output [64-1:0] l9erxxpnphqd26vg9,
  output [64-1:0] hig2gwwbeuhnt65xrp,
  input  [64-1:0] vf5xcr67bqhzlo43_,

  input  [64-1:0] vmx1fh4kmh4c,

  input  [64-1:0] v09gw6e6rfjf05qg,

  output s5f_36xvqrtq7,

  output u83p4flbuvkqt26z,
  output tvglhc8o_izdq,
  output siifnhwgancn8,
  output mfzl2fqml69hx,
  output aw0hbwfkx3f63s,

  output v9dnbgjy6c0vf,
  output hmzw4exmjn8k921c,
  output x6eltyshbu5,
  output lt3v_fm0ipu,
  output v3ne7glf8d8,



  input btwmhh91h50d5flgwx4o6pwu,

  input [2-1:0] r21i4by0bu3ks,
  input zmwq3e9oijvo7d7,

  input  sxvvsxtbhyvt,
  
    
  output j0qaxhuqtdi,
  output pbzpk52jinfscit4mm,
  output gwj6ow6qvbhs0tc31,
  output [12-1:0] mm0ssgy582fv_j,
  output iwdkm52x_w4hpak_a2_w,
  output  [64-1:0] ir2913p9xpmq_1bvfd1,
  input  [64-1:0] bsjo0v5e0t556pph,
  input  mwegg_7inaca6povsw,
  input  wnkp7091zrsevkbl,


  input  pydatzxqqi,

  output aw82i964do,
  output cwwkpmk260lrt,
  output rvr30vvllni,
  output y8_gkxsfle,
  output z1cj655u31,
  output lhu2z948o3n,

  input [64-1:0] wtd_nuaeb_mpye,
  input x7eg618xaszd4f21cl_g,
  input [64-1:0] xd66pm611ai1dg,
  input r9uxubpl2h2alj1q,

  input [64-1:0] elth4vimq_j,




  input ftp0juzjm2b587cyw5,

  input jlud6jeuxe0espga,



  input sf0uuehfhfa,
  input z35xlcc6bt4,
  input hvy2cpsp75f3,
  input k3z202os,

  input [64-1:0] ew08uu2kn2p9e11s,
  input xv08lot3vi9dag4vs0,
  input [64-1:0] mtc04rctrfyb,
  input if5jz8qk0aqefy3v35o,

  input rrujrlc85mhm,

  input jw4fsjecr0u919fr7,

  output[64-1:0]  pldoasxyzlvx2,
  output[64-1:0]  p6rw9no76a3m,
  output[64-1:0]  vyxop00ua6vr,



  output[64-1:0]     unbt3q05xijb,
  output[64-1:0]     hawbmpz6j7pzibqr,



  output [64-1:0]     r4bs4k_53n5wp,
  output [64-1:0]     i7lgezdqu4bmka,

  output [64-1:0]     h_qwsgi7nk2,
  output [64-1:0]  bde41te346q515l,
  output [64-1:0]     tvh1llq2i3_y,
  output                      w632tcbtqncn6,

  output                      ai169tbqp4seb3,
  output                      b0zz_ornhz010,
  output                      yw4o4kdms07_32,
  output                      ezl3jzeqhltgj7h,
  output                      w529wbj853,
  output                      i9xvsmm45fp0f58,


  input  [64-1:0]     u25pqekq4df,
  input                       dhjwho76fa8hqc,
  input  [64-1:0]     xel6gw173w5x0,
  input                       icauf4l_12_c2xkj53lf,
  input  [64-1:0]     v8ydjtlz16x9tx,
  input                       e_z6d7r9kxqg32te,
  input  [64-1:0]  p5jpgn4rvarpo,
  input                       z2g63deibg1b1quqr,
  input  [64-1:0]     tlgcdv86voe9,
  input                       u_ufp_wg29ieoklxxz1,
  input                       s_m3pbf5m2tr6v,

  input  [64-1:0]     bj7h5jqg66r51jxki6emra,
  output [64-1:0]     zmfo8cca_77pc,

  input                       miax48k27o484e8a,

  output [7:0]                tcy_87vt9vet39knuw,
  input                       fc_4ns_w1nh4h02z_dgg, 
  output                      fzdb65fcrotwcaccus_cwo,

  output[64-1:0]   d3hccrck1fl7jjf6,
  output                      vkyge0q4mfc5,
  output [64-1:0]     cppkd01vpwwnlfy,

  output                      psx330qmvh5so1to4iq,
  output                      sefocn4wjn2k2f_zvlvnz,  
  output                      qknomh2kbth19r1osddvzly,  
  output                      bzz8x0np0dpmdjt1d0w7uf,  
  output                      rl9a96pgy3troiao05jel,  
  output [64-1:0]  hzsp_nydab9ghw59v,  


  input [31:0]           ij_sgq3rtvw2,
  input [31:0]           k9jntnqwqp,

  output                b0ry73kp6sc2,          
  output                hr64e6c3gy,          
  output                cz1hh6af7xp2,          
  output [1:0]          st2zalpx0uf,
  output [1:0]          w30ye15yns15,
  output                ni01kj42oob2x,          
  output                ah8kjlmvnaxzbi,          
  output                fkuqlh34r,          
  output [16-1:0] hnc10arn_rd,
  output [20-1:0]   b2ulqcjb,


  input  dk2xhkj77a,
  input  gf33atgy,
  input  ru_wi

  );
    
  localparam yka1tofub6dvhok = 12;

  localparam urjif1vu4pqgqxt4x8 = 51;
  localparam m_rz39tx6bnugdx = (urjif1vu4pqgqxt4x8<=2)?1:(urjif1vu4pqgqxt4x8<=4)?2:(urjif1vu4pqgqxt4x8<=8)?3:(urjif1vu4pqgqxt4x8<=16)?4:(urjif1vu4pqgqxt4x8<=32)?5:(urjif1vu4pqgqxt4x8<=64)?6:(urjif1vu4pqgqxt4x8<=128)?7:(urjif1vu4pqgqxt4x8<=256)?8:(urjif1vu4pqgqxt4x8<=512)?9:(urjif1vu4pqgqxt4x8<=1024)?10:(urjif1vu4pqgqxt4x8<=2048)?11:(urjif1vu4pqgqxt4x8<=4096)?12:-1;
  localparam v_1vibiyou7ysbpkunv = (urjif1vu4pqgqxt4x8  < 32) ? 8 : (m_rz39tx6bnugdx + 3);
  localparam ob0j3iecn59nr6s8ur   = (m_rz39tx6bnugdx < yka1tofub6dvhok) ? yka1tofub6dvhok : m_rz39tx6bnugdx;




      
wire ntlp7re07dp6nkb;

wire u2dvoyt5e7o_03z9z5;
wire f982i0gj5cmkoid;
wire iu2o274ax6rzokmi0;
wire l_jd4i6dsmcejyydh;
wire brfqcqo_b08lybzgt;
wire ve7t8hdsd1_tnt9v;

assign kakelc68be0x7tdm9b9o  = (~u2dvoyt5e7o_03z9z5) 
                           | ntlp7re07dp6nkb 
                           ;
assign gm1r5itc44uxw_y0_msk =   l_jd4i6dsmcejyydh 
                          | ve7t8hdsd1_tnt9v
                          | iu2o274ax6rzokmi0;
assign j3j1czgoam48vhs8auo = 
                      wnkp7091zrsevkbl 
                      | brfqcqo_b08lybzgt
                      | f982i0gj5cmkoid;

assign r0s7d8cr68i2qs1z = (a94vd35etec4 | el7_p8jit09) & (
                  kakelc68be0x7tdm9b9o 
                | j3j1czgoam48vhs8auo 
                | gm1r5itc44uxw_y0_msk
                );



wire izhvh9xxvwe2 =   a94vd35etec4 & rb050tnl & (~r0s7d8cr68i2qs1z) 
                    ;







wire [64-1:0] cause_r;

wire [1:0] status_priv_r;

assign aw82i964do = (status_priv_r == 2'b11); 

assign y8_gkxsfle = (status_priv_r == 2'b01); 

wire [1:0] gg_wcrbxzhh0uqxd;
wire d97fz0kv80e8so8  = (gg_wcrbxzhh0uqxd == 2'b01);
wire tjggo01j7rusjv3a9g_bx = (gg_wcrbxzhh0uqxd == 2'b10);
wire vqzw2od29tt6hat  = (gg_wcrbxzhh0uqxd == 2'b11);
assign cwwkpmk260lrt = vqzw2od29tt6hat;
wire w3ouq_ntb6lrj_6yi = cause_r[64-1];

wire cmt_irq_mret_ena;
assign cmt_irq_mret_ena = w3ouq_ntb6lrj_6yi & rrujrlc85mhm;
wire upp957fldz7r621ml4u = (~w3ouq_ntb6lrj_6yi) & rrujrlc85mhm;  




wire [1:0] dttzf_6vv87y;








wire vvp82oplb = (dttzf_6vv87y == 2'b11); 

assign rvr30vvllni = vvp82oplb;

wire uhz5i6ah7vc1b9 = (dttzf_6vv87y == 2'b01); 
assign z1cj655u31 = uhz5i6ah7vc1b9;





wire dxb0y6x6tzh8_cwt2 = (e1go3iu == 12'h4CF);
wire ye9b2qmw0l_hy0n28 = dxb0y6x6tzh8_cwt2 & el7_p8jit09;


wire fb_inlkctcnic = (e1go3iu == 12'h300);



wire m_l49l2tvr3sko = fb_inlkctcnic & el7_p8jit09;



wire q2k15_wd423_d = fb_inlkctcnic & a94vd35etec4;



wire to3k3giu627wb2b7yd = (q2k15_wd423_d & izhvh9xxvwe2) ;





wire vb113ohv_p_qvfsa7;

wire qo6gz18vzk6paj = to3k3giu627wb2b7yd;
wire gjwsoz8iiwm4asx0 = vf5xcr67bqhzlo43_[22];

assign b0ry73kp6sc2 = vb113ohv_p_qvfsa7;

ux607_gnrl_dfflr #(1) nu0jcvn681am4sr8f (qo6gz18vzk6paj, gjwsoz8iiwm4asx0, vb113ohv_p_qvfsa7, gf33atgy, ru_wi);



wire dii97bgu2z_fae0;

wire igq0yfxfh5kzs5xq = to3k3giu627wb2b7yd;
wire vxg5wx02fk2q089y = vf5xcr67bqhzlo43_[21];

assign hr64e6c3gy = dii97bgu2z_fae0;

ux607_gnrl_dfflr #(1) fdhiozl882zqxxr (igq0yfxfh5kzs5xq, vxg5wx02fk2q089y, dii97bgu2z_fae0, gf33atgy, ru_wi);



wire xt17qz_76v42;

wire oucmpl1vq2mmm06 = to3k3giu627wb2b7yd;
wire cy50u1stw46zgb = vf5xcr67bqhzlo43_[20];

assign cz1hh6af7xp2 = xt17qz_76v42;

ux607_gnrl_dfflr #(1) akh_979wckg50gchaz08 (oucmpl1vq2mmm06, cy50u1stw46zgb, xt17qz_76v42, gf33atgy, ru_wi);



wire hkl71xhnekm20fk;



wire rz377ucxvdy = s_m3pbf5m2tr6v;
wire glvudafm82gm = rrujrlc85mhm & ~rvr30vvllni;

wire d3ajn2bv7ru6veccs3 = 

        rz377ucxvdy |
        glvudafm82gm |
        to3k3giu627wb2b7yd;

wire g0v2ifpvvpr9zatcqgw = to3k3giu627wb2b7yd ? vf5xcr67bqhzlo43_[17] :
                       rz377ucxvdy     ? 1'b0             :
                                       1'b0             ;

ux607_gnrl_dfflr #(1) xshngwlz8dxgjgagpcfl (d3ajn2bv7ru6veccs3, g0v2ifpvvpr9zatcqgw, hkl71xhnekm20fk, gf33atgy, ru_wi);





wire maka6zd0las79r5dg5 = 
        
        z2g63deibg1b1quqr | 
        
        s_m3pbf5m2tr6v | 

        jlud6jeuxe0espga | 






        jw4fsjecr0u919fr7 |
        rrujrlc85mhm  






        ;


wire ogmro605vz43jd_a6;
wire [1:0] gah2y9c1ou_ln8ix8;

assign gah2y9c1ou_ln8ix8 = 

               jlud6jeuxe0espga ? 2'b11 :
        
               jw4fsjecr0u919fr7 ? r21i4by0bu3ks : 

               rrujrlc85mhm ? dttzf_6vv87y :
        
               z2g63deibg1b1quqr ? 2'b01 :     
        
               s_m3pbf5m2tr6v ? {1'b0,ogmro605vz43jd_a6} : 
                              status_priv_r;

              
ux607_gnrl_dfflrs #(2) jfld0h0k3gxyya7xz (maka6zd0las79r5dg5, gah2y9c1ou_ln8ix8, status_priv_r, gf33atgy, ru_wi);


assign rm1dxjejhq7dh3q5m = hkl71xhnekm20fk;


wire [1:0]     edu3vzxs7stp;
wire           idq_m7lglm;
wire           r1u74u2bcei1;
wire [2:1]     rlsnapd43j6;
wire           d63fiicib; 


wire cmt_irq_epc_ena;
assign cmt_irq_epc_ena= hvy2cpsp75f3 & jlud6jeuxe0espga;
wire ysdq7a_idp9m94_7qcva= cmt_irq_epc_ena & k3z202os;
wire wew7vt2_2h6k = (e1go3iu == 12'h345);
wire xcfnsabp39vvwn = (e1go3iu == 12'h7ED);
wire lg08w1fgrqdmj2trv50pi_; 
wire i8a3q6ebfamt1jmd4be2qh3;
wire aval5ewiun = ysdq7a_idp9m94_7qcva 
               | i8a3q6ebfamt1jmd4be2qh3
              ;
wire m5zfpzj06s9bxq;



wire d9w566umxhr1msc5h_;



wire tisldbai0191pm41m7  = 
    lg08w1fgrqdmj2trv50pi_ | 

       jlud6jeuxe0espga



     | rrujrlc85mhm 
     | to3k3giu627wb2b7yd
        ;

wire jxhi9cr3nbjdng6297  = 
    lg08w1fgrqdmj2trv50pi_ ? (
                        xcfnsabp39vvwn ? 1'b1 :
        guuvp01vkcryglsu1p3[3]) :






     jlud6jeuxe0espga ? 1'b0 :









    rrujrlc85mhm ? d9w566umxhr1msc5h_ :

    to3k3giu627wb2b7yd ? vf5xcr67bqhzlo43_[3] : 
                  s5f_36xvqrtq7; 

ux607_gnrl_dfflr #(1) smo2std8m7ao_oxeipz4 (tisldbai0191pm41m7, jxhi9cr3nbjdng6297, s5f_36xvqrtq7, gf33atgy, ru_wi);



















wire a96rxse5wp61642f61up;
wire kakkebd37ke18jyiv2sujpliozz = a96rxse5wp61642f61up & dn8riluj40uunvq5;
wire y0gytfbi3n3ba_mn  = 
       jlud6jeuxe0espga
     | rrujrlc85mhm 
     | kakkebd37ke18jyiv2sujpliozz   
     | to3k3giu627wb2b7yd;

wire gsuwcm3ksdxfts2_wgm = y0gytfbi3n3ba_mn;



wire [1:0] ial7ihq_lscsphgdii;













wire [1:0] r1cznjd8rub5fb1xpx1 =
                                      2'b00
                                  ;

wire  [64-1:0] uiulkx67fwpf7in8sde_kj;

assign ial7ihq_lscsphgdii = 

                jlud6jeuxe0espga ? status_priv_r : 


                rrujrlc85mhm ? 
                                  (w3ouq_ntb6lrj_6yi ? r1cznjd8rub5fb1xpx1 : rlsnapd43j6) :

                to3k3giu627wb2b7yd ? vf5xcr67bqhzlo43_[12:11] :
                 kakkebd37ke18jyiv2sujpliozz ?  uiulkx67fwpf7in8sde_kj[29:28]   : 
                                dttzf_6vv87y;


wire au4016pzmaqihyvwn6    = 





    jlud6jeuxe0espga ? s5f_36xvqrtq7 :






    rrujrlc85mhm  ? 
                                  (w3ouq_ntb6lrj_6yi ? 1'b1 : d63fiicib) :


    to3k3giu627wb2b7yd ? vf5xcr67bqhzlo43_[7] : 
      kakkebd37ke18jyiv2sujpliozz  ?  uiulkx67fwpf7in8sde_kj[27]:
                  d9w566umxhr1msc5h_; 

              
ux607_gnrl_dfflr #(2) at9q041uhsjnc881 (gsuwcm3ksdxfts2_wgm, ial7ihq_lscsphgdii, dttzf_6vv87y, gf33atgy, ru_wi);


ux607_gnrl_dfflr #(1) vbzyttr8v84p3dmckct8v (y0gytfbi3n3ba_mn, au4016pzmaqihyvwn6, d9w566umxhr1msc5h_, gf33atgy, ru_wi);






































































































































wire [1:0] yon43wm5u290o = 2'b10;








wire [1:0] nriqmhgyl2409 = 2'b10;







wire [1:0] l56q7o0hmnd98qc_;
wire [1:0] i8uou0fe4qb;
wire d6z8hz6u7gym = (l56q7o0hmnd98qc_ == 2'b11) | (i8uou0fe4qb == 2'b11);

wire b3lm_1ct7augo;








   
assign i8uou0fe4qb = 2'b0; 

wire [64-1:0] ilicr1czem8;
wire [64-1:0] klnr5w9m7dv5ejwl; 



wire f2n39xbpvn9k = a96rxse5wp61642f61up | r9uxubpl2h2alj1q;

wire [64-1:0] yrf31busye76;


assign kbv2bs_lxmvu = yrf31busye76;

wire [7:0] qrkpl4iy0;

wire [64-1:0] mintstatus_r;
wire [64-1:0] sintstatus_r;
assign gfy3zost37aq8qmr = (mintstatus_r != 64'b0) | (sintstatus_r != 64'b0);
wire i7e201yj = (e1go3iu == 12'h307);
wire kp2q6bh2 = el7_p8jit09 & i7e201yj;
wire yrwzf3cdms = a94vd35etec4 & i7e201yj;
wire g2y8t8mc94ns = (yrwzf3cdms & izhvh9xxvwe2);
wire [64-1:0] a93w0kejmfr0l =  {vf5xcr67bqhzlo43_[64-1:v_1vibiyou7ysbpkunv],{v_1vibiyou7ysbpkunv{1'b0}}}; 
wire [64-1:0] yc3tkcusq6;
ux607_gnrl_dfflr #(64) gy1tc7gb8fpv2xa (g2y8t8mc94ns, a93w0kejmfr0l, yc3tkcusq6, gf33atgy, ru_wi);
wire [64-1 :0] ptzmif3v0ur = yc3tkcusq6;
wire [64-1:0] tuh58_qx = yc3tkcusq6; 
assign z0yhjfv_e0yaa2r = {tuh58_qx[(64-1):(m_rz39tx6bnugdx+3)],b4lwcgm6l21pi[m_rz39tx6bnugdx-1:0],3'b0};

wire wsps0651m = (e1go3iu == 12'h7EC);
wire crgfb_c8n = el7_p8jit09 & wsps0651m;
wire uli1h7sbvq = a94vd35etec4 & wsps0651m;
wire wcukhy5hjx = (uli1h7sbvq & izhvh9xxvwe2);
  
wire [64-1:0] pty14rphd3 =  {vf5xcr67bqhzlo43_[64-1:2],1'b0,vf5xcr67bqhzlo43_[0]}; 
wire [64-1:0] nzfqkqop6l_a;
ux607_gnrl_dfflr #(64) p83skg7wjlx5dbsl (wcukhy5hjx, pty14rphd3, nzfqkqop6l_a, gf33atgy, ru_wi);
wire [64-1 :0] o3zhp2khg52i02 = nzfqkqop6l_a;
assign yrf31busye76 = nzfqkqop6l_a; 
assign o7hoht1pqz01v7 = yrf31busye76[0];



wire xpjx62p088i2vk_7ow4_acag;
wire mx6n8ae8twuk2mfjz_1 = (e1go3iu == 12'h346);
wire xlchao2g44p1tat_ = el7_p8jit09 & mx6n8ae8twuk2mfjz_1;
wire f1h7j_1pqx0g5v_ytwp =dn8riluj40uunvq5 & ( xpjx62p088i2vk_7ow4_acag
                                     | cmt_irq_epc_ena
                                     | cmt_irq_mret_ena); 

wire [64-1:0] jjb_1mrucinqpoy7nx4 = (xpjx62p088i2vk_7ow4_acag | cmt_irq_epc_ena) ? {{(64-32){1'b0}}, hjrk_rwjkqj3zk_b, 24'b0}   :
                                                                 cmt_irq_mret_ena ? {{(64-32){1'b0}}, qrkpl4iy0, 24'b0}         :
                                                                                    mintstatus_r;
ux607_gnrl_dfflr #(64) xtt6fx5zakc3pnmhdfy (f1h7j_1pqx0g5v_ytwp, jjb_1mrucinqpoy7nx4, mintstatus_r, gf33atgy, ru_wi);
wire [64-1:0] t7gzjhdzm9ftqnv7 = {mintstatus_r[64-1:24],8'h0,sintstatus_r[15:8],8'b0};
assign f_i1959b4xizzq9jea = mintstatus_r[31:24];

wire cgnhh8s1vo2cuntv = (e1go3iu == 12'h349);
wire zcege9lvdnn7d5f = el7_p8jit09 & cgnhh8s1vo2cuntv;
wire vto97yswc40s3 = (qrkpl4iy0 == 8'b0);
wire sokggdu75vi12fa2u3x9t2cq = (f_i1959b4xizzq9jea[7:0] == 8'b0);
wire myir1xya1lclgbvmhr = (vto97yswc40s3 != sokggdu75vi12fa2u3x9t2cq) & cgnhh8s1vo2cuntv & dn8riluj40uunvq5;
wire qphloyvbjzxcmxgms8sz9x7_5tk = izhvh9xxvwe2 & myir1xya1lclgbvmhr; 
wire [64-1:0] sotpl4qsv5jjhbht = myir1xya1lclgbvmhr ? klnr5w9m7dv5ejwl : vmx1fh4kmh4c;
wire [64-1:0] ixkez_bglcky89d58tfw3 = dn8riluj40uunvq5 ? sotpl4qsv5jjhbht : 64'b0; 


wire p7zidsgtr9q7bf81 = (e1go3iu == 12'h348);
wire ka2utev6jddufp7b9 = el7_p8jit09 & p7zidsgtr9q7bf81;
wire jywijmrdzis83sxzu = p7zidsgtr9q7bf81 & (dttzf_6vv87y != status_priv_r);
wire t_9kasosfl9_37azg4trv40ag0ch = izhvh9xxvwe2 & jywijmrdzis83sxzu; 
wire [64-1:0] hxxl4aq4sjdycyml2 = jywijmrdzis83sxzu ? klnr5w9m7dv5ejwl : vmx1fh4kmh4c;

wire gkxo6i5s875r = el7_p8jit09 & xcfnsabp39vvwn;

wire hcqw9t9s = el7_p8jit09 & wew7vt2_2h6k;

wire l9cidu8f0jn07fiqnf3i = wew7vt2_2h6k 
                       | xcfnsabp39vvwn 
                       ;

wire a6364gu6x8g_wiv = l9cidu8f0jn07fiqnf3i  
                        & znzjygllppv1s0a8cqub3c  
                        & gfy3zost37aq8qmr
                        & (hjrk_rwjkqj3zk_b > qrkpl4iy0)
                        & (~zwcbp7zqfei5xz) 
                        & dn8riluj40uunvq5;

assign xpjx62p088i2vk_7ow4_acag = a6364gu6x8g_wiv & izhvh9xxvwe2;
wire t758474hjb_u9x_qz5jrw2x = xpjx62p088i2vk_7ow4_acag;

wire [64-1:0] jlm7v1b79iuln;
assign  jlm7v1b79iuln = {ptzmif3v0ur[(64-1):(m_rz39tx6bnugdx+3)],b4lwcgm6l21pi[m_rz39tx6bnugdx-1:0],3'b0};


wire [64-1:0] cyxvmxf7k3h7 = a6364gu6x8g_wiv ? 
                                          jlm7v1b79iuln 
                                          : 64'b0;


assign dxi_ue3gf5zqqqxwgq2a = xpjx62p088i2vk_7ow4_acag;
assign lg08w1fgrqdmj2trv50pi_ = l9cidu8f0jn07fiqnf3i & izhvh9xxvwe2;

wire [64-1:0] igbraabs1 = a6364gu6x8g_wiv ? 
                                   nchi0_6mu
                                   : vmx1fh4kmh4c;

wire [64-1:0] pltp40lm289gs = dn8riluj40uunvq5 ?  igbraabs1 : 64'b0;

assign bisaqpu86vneunhkqtg = dxi_ue3gf5zqqqxwgq2a & xcfnsabp39vvwn;  
assign jathu3ui07hzkaq4g2z39  = jlm7v1b79iuln[64-1:0]; 
assign pl2up5ze0wczfdx0ga70d  = 1'b1;
assign a5_uct872oszxvfp4kn_  = pydatzxqqi;
assign m3ar1m0lklmpw4oek2yjd3ev  = aw82i964do;
assign zk19lxmoqrzcdjx6rxuvc36  = y8_gkxsfle;
assign i8a3q6ebfamt1jmd4be2qh3  = bisaqpu86vneunhkqtg & pl2up5ze0wczfdx0ga70d;

wire dfkhf0zzmeauwtqm3som;

wire iiq92rsh_v1ylb;

wire sim0gblc86voze3mam;
wire wft1k16f78xw2;


wire b00s0p78drh4z   = (e1go3iu == 12'h7a1);
wire lxcp51g29nqalv   = (e1go3iu == 12'h7a2);
wire tzfj8xp6rkw   = (e1go3iu == 12'h7a3);
wire mdl08rw1652e5 = b00s0p78drh4z | lxcp51g29nqalv | tzfj8xp6rkw;
wire c6lbvkska6qd     = (e1go3iu == 12'h7b0);


wire vqvbmvk4f_b_c;

assign xsekawjaoeqedkdymhz6h = izhvh9xxvwe2 & 








                          (   
                              1'b0
                              | mdl08rw1652e5
                              | sim0gblc86voze3mam
                              | dxb0y6x6tzh8_cwt2
                              
                              | dfkhf0zzmeauwtqm3som
                              | fb_inlkctcnic   
                              | c6lbvkska6qd
                              | vqvbmvk4f_b_c
                              | wft1k16f78xw2
                          )
                          ;
assign b0cs5n_1_q64sumeg  = lovkp0eqfnxtb7;
assign fg6gtaxnx8a0anercx  = 1'b0;
assign d14swmczjaws9gr8uvx  = pydatzxqqi;
assign vsrfdna3ksbt8a__05sjdxr  = aw82i964do;
assign uttwdi1xwyv_l7uzt3x2ea  = y8_gkxsfle;











   
   
   
   
   
   
   
   

wire zijl1miri7deso9se;
wire qy7n657jeoo8 = 
         ya8t4ev_aidf0t0x4or 
       | zijl1miri7deso9se;  

        
wire v5xf85uoa2mep  = 
        
        to3k3giu627wb2b7yd |
        b3lm_1ct7augo |
        
        (qy7n657jeoo8 & (~rnx27onf2lbe));

wire [1:0] mhlxmr2avg00i3aee5  = 
        
        to3k3giu627wb2b7yd ? vf5xcr67bqhzlo43_[14:13] : 
        b3lm_1ct7augo ? vf5xcr67bqhzlo43_[14:13] : 
        
        (qy7n657jeoo8 & (~rnx27onf2lbe)) ? 2'b11 :
                        l56q7o0hmnd98qc_;

ux607_gnrl_dfflr #(2) e2zyg2k5653e7w62s1t (v5xf85uoa2mep, mhlxmr2avg00i3aee5, l56q7o0hmnd98qc_, gf33atgy, ru_wi);





wire [64-1:0] csr_mstatus;
wire [64-1:0] csr_sstatus;
wire [64-1:0] csr_sie;
wire [64-1:0] csr_sip;




assign csr_mstatus[64-1]    = d6z8hz6u7gym;                        
assign csr_mstatus[64-2:36] = 27'b0;
assign csr_mstatus[35:34] = yon43wm5u290o;
assign csr_mstatus[33:32] = nriqmhgyl2409;
assign csr_mstatus[31]    = 1'b0; 

assign csr_mstatus[30:23] = 8'b0; 
assign csr_mstatus[22]    = vb113ohv_p_qvfsa7;                       
assign csr_mstatus[21]    = dii97bgu2z_fae0;                        
assign csr_mstatus[20]    = xt17qz_76v42;                       
assign csr_mstatus[19]    = csr_sstatus[19];                    
assign csr_mstatus[18]    = csr_sstatus[18];                    
assign csr_mstatus[17]    = hkl71xhnekm20fk;                      
assign csr_mstatus[16:15] = i8uou0fe4qb;                        
assign csr_mstatus[14:13] = l56q7o0hmnd98qc_;                        
assign csr_mstatus[12:11] = dttzf_6vv87y;                       
assign csr_mstatus[10:9]  = 2'b0; 
assign csr_mstatus[8]     = csr_sstatus[8];                     
assign csr_mstatus[7]     = d9w566umxhr1msc5h_;                      
assign csr_mstatus[6]     = 1'b0; 
assign csr_mstatus[5]     = csr_sstatus[5];                     
assign csr_mstatus[4]     = 1'b0;               
assign csr_mstatus[3]     = s5f_36xvqrtq7;                       
assign csr_mstatus[2]     = 1'b0; 
assign csr_mstatus[1]     = csr_sstatus[1];                     
assign csr_mstatus[0]     = 1'b0;               





















wire jan2q6micau0n4 = (e1go3iu == 12'h302);
wire ls8dsrnc8qwzmpg = (e1go3iu == 12'h303);

wire xd1ve1tqh9v = jan2q6micau0n4 & el7_p8jit09;
wire ekglglw24_squr = ls8dsrnc8qwzmpg & el7_p8jit09;

wire [64-1:0] csr_medeleg;
wire [64-1:0] csr_mideleg;






wire s5vf28d55rgucs = jan2q6micau0n4 & a94vd35etec4;
wire nreobds793ur = s5vf28d55rgucs & izhvh9xxvwe2;

wire [64-1:0] rut11ws_0t00uq;
wire [64-1:0] zmlt8meq9wrm0gym;

assign zmlt8meq9wrm0gym[8:0] = vf5xcr67bqhzlo43_[8:0];
assign zmlt8meq9wrm0gym[10:9]  = 2'b0; 

assign zmlt8meq9wrm0gym[11]  = 1'b0;
assign zmlt8meq9wrm0gym[12] = vf5xcr67bqhzlo43_[12];
assign zmlt8meq9wrm0gym[13] = vf5xcr67bqhzlo43_[13];
assign zmlt8meq9wrm0gym[14] = 1'b0;
assign zmlt8meq9wrm0gym[15] = vf5xcr67bqhzlo43_[15];
assign zmlt8meq9wrm0gym[16]  = 1'b0;
assign zmlt8meq9wrm0gym[64-1:17] = 15'b0;

ux607_gnrl_dfflr #(64) wlb1_8fd6dkg3fo (nreobds793ur, zmlt8meq9wrm0gym, rut11ws_0t00uq, gf33atgy, ru_wi);

assign csr_medeleg = rut11ws_0t00uq;
assign r4bs4k_53n5wp = csr_medeleg;    





wire bx1uul6oagk85s = ls8dsrnc8qwzmpg & a94vd35etec4;
wire igy7k5am9dh9hwt = (~dn8riluj40uunvq5) & bx1uul6oagk85s & izhvh9xxvwe2;

wire [64-1:0] cwtczyq3t3b;
wire [64-1:0] bz_fv6kksgjdp5;
assign bz_fv6kksgjdp5[1:0]   = vf5xcr67bqhzlo43_[1:0];
assign bz_fv6kksgjdp5[2]     = 1'b0;
assign bz_fv6kksgjdp5[5:3]   = vf5xcr67bqhzlo43_[5:3];
assign bz_fv6kksgjdp5[6]     = 1'b0;
assign bz_fv6kksgjdp5[9:7]   = vf5xcr67bqhzlo43_[9:7];
assign bz_fv6kksgjdp5[10]    = 1'b0;
assign bz_fv6kksgjdp5[11]    = vf5xcr67bqhzlo43_[11];
assign bz_fv6kksgjdp5[31:12] = 20'b0;

assign bz_fv6kksgjdp5[64-1:32] = {64-32{1'b0}};

ux607_gnrl_dfflr #(64) jpptf75jlhmmxymhc (igy7k5am9dh9hwt, bz_fv6kksgjdp5, cwtczyq3t3b, gf33atgy, ru_wi);

assign csr_mideleg = dn8riluj40uunvq5 ? 32'b0 : cwtczyq3t3b;
assign i7lgezdqu4bmka = csr_mideleg;     



wire ps869z4s = (e1go3iu == 12'h304);
wire wwc6g7 = ps869z4s & el7_p8jit09;
wire fx8mak0qu = ps869z4s & a94vd35etec4;
wire yw2rjoyrops = (~dn8riluj40uunvq5) & fx8mak0qu & izhvh9xxvwe2;
wire [64-1:0] aohjw;
wire [64-1:0] zlkg60c;
assign zlkg60c[64-1:22] = {(64-22){1'b0}};
assign zlkg60c[21] = 1'b0;
assign zlkg60c[20] = 1'b0;
assign zlkg60c[19] = 1'b0;
assign zlkg60c[18] = vf5xcr67bqhzlo43_[18];
assign zlkg60c[17] = vf5xcr67bqhzlo43_[17];
assign zlkg60c[16] = 1'b0;
assign zlkg60c[15:12] = 4'b0;
assign zlkg60c[11] = vf5xcr67bqhzlo43_[11];
assign zlkg60c[10:8] = 3'b0;
assign zlkg60c[ 7] = vf5xcr67bqhzlo43_[ 7];
assign zlkg60c[6:4] = 3'b0;
assign zlkg60c[ 3] = vf5xcr67bqhzlo43_[ 3];
assign zlkg60c[2:0] = 3'b0;
ux607_gnrl_dfflr #(64) tt3rnfqu_x7no (yw2rjoyrops, zlkg60c, aohjw, gf33atgy, ru_wi);
wire [64-1:0] csr_mie;
assign csr_mie = dn8riluj40uunvq5 ? 64'b0 : {aohjw[64-1:10],ai169tbqp4seb3,1'b0,aohjw[7:6],b0zz_ornhz010,1'b0,aohjw[3:2],yw4o4kdms07_32,1'b0};
assign tvglhc8o_izdq  = csr_mie[18];
assign u83p4flbuvkqt26z = csr_mie[16];
assign aw0hbwfkx3f63s = csr_mie[11];
assign siifnhwgancn8 = csr_mie[ 7];
assign mfzl2fqml69hx = csr_mie[ 3];






wire yoegchl8 = (e1go3iu == 12'h344);
wire oekhv_ = yoegchl8 & el7_p8jit09;
wire eunacz7 = (~dn8riluj40uunvq5) & yoegchl8 & a94vd35etec4;
wire gan2wxwq9 = eunacz7 & izhvh9xxvwe2;







wire l0hrd_ubxbkay3zy8yz;
assign ix299qulxi5 = l0hrd_ubxbkay3zy8yz;
wire mpe6p6hnhph9k_6d = (~dn8riluj40uunvq5) & ix299qulxi5;
wire cz0vkccbbonhv7 = cmt_irq_epc_ena & (k3cmpuswk7in0u4 == 12'd18);
wire pfztq9p448ixclu5fvp = mpe6p6hnhph9k_6d | (~cz0vkccbbonhv7);
wire vceay__vidby7u2pyk = gan2wxwq9 | mpe6p6hnhph9k_6d | cz0vkccbbonhv7;
wire zovis90gyknz23paxn = gan2wxwq9 ? vf5xcr67bqhzlo43_[18] : pfztq9p448ixclu5fvp;
ux607_gnrl_dfflr #(1) kj1ejs6kvfjb8e6p (vceay__vidby7u2pyk, zovis90gyknz23paxn, hmzw4exmjn8k921c, gf33atgy, ru_wi);



assign jjj61w03m77lv = 1'b0;
assign v9dnbgjy6c0vf = 1'b0;


wire xc_4r6ncv72 = cwtczyq3t3b[1];
wire m00o8sz4cyd_a9 = cwtczyq3t3b[5];
assign x_cq40qmp6a = cwtczyq3t3b[9];

assign x6eltyshbu5 = xx87vzbpchg & (~m00o8sz4cyd_a9);
assign lt3v_fm0ipu = pvfk1_6o89lmby & (~xc_4r6ncv72);
assign v3ne7glf8d8 = zz5wo47gw146x4;

wire [64-1:0] j4k2ts6t;
wire [64-1:0] csr_mip;

assign j4k2ts6t[64-1:22] = {(64-22){1'b0}};
assign j4k2ts6t[21] = 1'b0;
assign j4k2ts6t[20] = 1'b0;
assign j4k2ts6t[19] = 1'b0;
assign j4k2ts6t[18] = hmzw4exmjn8k921c;
assign j4k2ts6t[17] = 1'b0;
assign j4k2ts6t[16] = v9dnbgjy6c0vf;
assign j4k2ts6t[15:12] = 4'b0;
assign j4k2ts6t[11] = v3ne7glf8d8;
assign j4k2ts6t[10] = 1'b0;
assign j4k2ts6t[ 9] = ezl3jzeqhltgj7h;
assign j4k2ts6t[ 8] = 1'b0;
assign j4k2ts6t[ 7] = x6eltyshbu5;
assign j4k2ts6t[ 6] = 1'b0;
assign j4k2ts6t[ 5] = w529wbj853;
assign j4k2ts6t[ 4] = 1'b0;
assign j4k2ts6t[ 3] = lt3v_fm0ipu;
assign j4k2ts6t[ 2] = 1'b0;
assign j4k2ts6t[ 1] = i9xvsmm45fp0f58;
assign j4k2ts6t[ 0] = 1'b0;

assign csr_mip = dn8riluj40uunvq5 ? 64'b0 : j4k2ts6t;



wire etyac0jmfrzxm = (e1go3iu == 12'h305);
wire t4fpmjlqyt = el7_p8jit09 & etyac0jmfrzxm;
wire s415nowb_m = etyac0jmfrzxm & a94vd35etec4;
wire swsoaue2vpdpr = (s415nowb_m & izhvh9xxvwe2);
wire [64-1:0] jb2zldqg;
wire [64-1:0] gir1qkzddwv = vf5xcr67bqhzlo43_[64-1:0];
ux607_gnrl_dfflr #(64) v9a0wulyijcit4 (swsoaue2vpdpr, gir1qkzddwv, jb2zldqg, gf33atgy, ru_wi);
wire [64-1:0] p41zr5gkln = dn8riluj40uunvq5 ? jb2zldqg : {jb2zldqg[64-1:2],2'b0};
assign unbt3q05xijb = p41zr5gkln;



wire b9p2i13nz = (e1go3iu == 12'h7c3);
wire ycvvi2q5 = el7_p8jit09 & b9p2i13nz;


wire [64-1:0] glwac019m8pq = w2fpnf5fg1byp6 ? p41zr5gkln : wd9dvepxj;


assign hawbmpz6j7pzibqr = glwac019m8pq;



wire l52o_50oot2j6 = (e1go3iu == 12'h340);
wire rud1hmcy9tubf9k = l52o_50oot2j6 & el7_p8jit09;
wire ujw7_8d4aou = l52o_50oot2j6 & a94vd35etec4;
assign pby60vfdze02 = (ujw7_8d4aou & izhvh9xxvwe2) | t_9kasosfl9_37azg4trv40ag0ch | qphloyvbjzxcmxgms8sz9x7_5tk;
wire [64-1:0] mscratch_r;
assign vm3pyzc9nt95 = vf5xcr67bqhzlo43_;
ux607_gnrl_dfflr #(64) gri20em6huxaawv (pby60vfdze02, vm3pyzc9nt95, mscratch_r, gf33atgy, ru_wi);
assign klnr5w9m7dv5ejwl = mscratch_r;





















wire b8m44m4dqrd = (e1go3iu == 12'h341);
wire bk92fvsycux = b8m44m4dqrd & el7_p8jit09;
wire qj8fyo_ = b8m44m4dqrd & a94vd35etec4;
wire hagyoc47ea = (qj8fyo_ & izhvh9xxvwe2) | jlud6jeuxe0espga 
               | upp957fldz7r621ml4u
               ;
wire [64-1:0] czcawgfux3h7; 

wire [64-1:0] mzvpa_lx;
wire [64-1:0] bo81ykm6;


assign bo81ykm6[64-1:1] = 
        jlud6jeuxe0espga ? elth4vimq_j[64-1:1] :
        upp957fldz7r621ml4u ? czcawgfux3h7[64-1:1] :
        vf5xcr67bqhzlo43_[64-1:1];
assign bo81ykm6[0] = 1'b0;
ux607_gnrl_dfflr #(64) ghe2y0gfj2y (hagyoc47ea, bo81ykm6, mzvpa_lx, gf33atgy, ru_wi);
wire [64-1:0] csr_mepc;
assign csr_mepc = mzvpa_lx;
assign pldoasxyzlvx2 = mzvpa_lx;



























wire [1:0] a031mt59o9h2wubgw;






wire di2d3ktm1fz_8we = (e1go3iu == 12'h342);
wire k2zpid7lzqutl = di2d3ktm1fz_8we & el7_p8jit09;
assign m5zfpzj06s9bxq = di2d3ktm1fz_8we & a94vd35etec4;

assign a96rxse5wp61642f61up = 
               upp957fldz7r621ml4u |
               (m5zfpzj06s9bxq & izhvh9xxvwe2);

wire [64-1:0] qxyauqoyrj6kj; 
wire [64-1:0] t29y65qqvjjxvouca3; 
wire [64-1:0] emggndeggdfff68dw0; 

assign uiulkx67fwpf7in8sde_kj = 
               upp957fldz7r621ml4u ? qxyauqoyrj6kj :
               vf5xcr67bqhzlo43_;


assign ilicr1czem8[64-1]  = r9uxubpl2h2alj1q ? xd66pm611ai1dg[64-1] : uiulkx67fwpf7in8sde_kj[64-1];


assign ilicr1czem8[64-2:0] = {(64-1){1'b0}};
wire nbm3vo3_g;
assign dn8riluj40uunvq5 = (jb2zldqg[5:0] == 6'b11);
ux607_gnrl_dfflr  #(1) q5kg7vijybs7czw7jt (f2n39xbpvn9k, ilicr1czem8[64-1], cause_r[64-1], gf33atgy, ru_wi);
wire a44gbj7j9rxv0z8u = dn8riluj40uunvq5 & (a96rxse5wp61642f61up | aval5ewiun | enwn0u48p2_ls5az80);
wire cjeqbkzjih5bqe = aval5ewiun   ? 1'b1 :
                 enwn0u48p2_ls5az80 ? 1'b0 :
                 a96rxse5wp61642f61up   ? uiulkx67fwpf7in8sde_kj[30]:
                 nbm3vo3_g;
ux607_gnrl_dfflr  #(1) g2ioy27sv7mxe7u4c8auiv (a44gbj7j9rxv0z8u, cjeqbkzjih5bqe, nbm3vo3_g, gf33atgy, ru_wi);

wire yy3oakojfxha =  dn8riluj40uunvq5 & (cmt_irq_epc_ena | a96rxse5wp61642f61up);



wire [7:0] n6mca19y6u =   cmt_irq_epc_ena  ?  f_i1959b4xizzq9jea :
                        a96rxse5wp61642f61up   ?  uiulkx67fwpf7in8sde_kj[23:16] :
                        qrkpl4iy0;
ux607_gnrl_dfflr  #(8) ljde_yamnmmrrq8o (yy3oakojfxha, n6mca19y6u, qrkpl4iy0, gf33atgy, ru_wi);


wire xirflumwondxbesu = f2n39xbpvn9k | t758474hjb_u9x_qz5jrw2x;
wire [ob0j3iecn59nr6s8ur-1:0] yo5msmd5ht7wrj; 
wire [ob0j3iecn59nr6s8ur-1:0] i_mi6vrgn4y6y7bg = r9uxubpl2h2alj1q          ? xd66pm611ai1dg[ob0j3iecn59nr6s8ur-1:0] :
                                               t758474hjb_u9x_qz5jrw2x ? {{ob0j3iecn59nr6s8ur-m_rz39tx6bnugdx{1'b0}},b4lwcgm6l21pi[m_rz39tx6bnugdx-1:0]} 
                                             : uiulkx67fwpf7in8sde_kj[ob0j3iecn59nr6s8ur-1:0];

ux607_gnrl_dfflr  #(ob0j3iecn59nr6s8ur) fs6_dpydm_6h__gnmhnvz5 (xirflumwondxbesu,i_mi6vrgn4y6y7bg,yo5msmd5ht7wrj,gf33atgy,ru_wi);

assign cause_r[64-2:31] = {(64-32){1'b0}};
assign cause_r[30] = dn8riluj40uunvq5 ? nbm3vo3_g : 1'b0;
assign cause_r[29:28] =  dn8riluj40uunvq5 ? dttzf_6vv87y : 2'b0;
assign cause_r[27] =  dn8riluj40uunvq5 ? d9w566umxhr1msc5h_ : 1'b0;

assign cause_r[26:25] =  2'b0;
assign cause_r[24] = 1'b0;
assign cause_r[23:16] = dn8riluj40uunvq5 ? qrkpl4iy0 : 8'b0;
assign cause_r[15:ob0j3iecn59nr6s8ur] = {(16-ob0j3iecn59nr6s8ur){1'b0}};
assign cause_r[ob0j3iecn59nr6s8ur-1:0] = yo5msmd5ht7wrj;


assign p6rw9no76a3m = cause_r;





wire zavn9glbl0j62qi = (e1go3iu == 12'h343);
wire jbbx5w95zgs1 = zavn9glbl0j62qi & el7_p8jit09;
wire x19cn_wmb7i = zavn9glbl0j62qi & a94vd35etec4;
wire fsr4k75wyd83d46eyxmu1so = x7eg618xaszd4f21cl_g;
wire kg9jji1tok8zi = (x19cn_wmb7i & izhvh9xxvwe2) | fsr4k75wyd83d46eyxmu1so;
wire [64-1:0] ii7u725d3lqc;
wire [64-1:0] xp3cg4k96hrbwzi;
assign xp3cg4k96hrbwzi = fsr4k75wyd83d46eyxmu1so ? wtd_nuaeb_mpye : vf5xcr67bqhzlo43_[64-1:0];
ux607_gnrl_dfflr #(64) f6vtcg5uu4zjv5886b (kg9jji1tok8zi, xp3cg4k96hrbwzi, ii7u725d3lqc, gf33atgy, ru_wi);
wire [64-1:0] ga1zsr158e3cs9vru;
assign ga1zsr158e3cs9vru = ii7u725d3lqc;







wire by_qc3yb1cyytd = (e1go3iu == 12'h001);
wire fk5t4onucgv    = (e1go3iu == 12'h002);
wire lc6w646en   = (e1go3iu == 12'h003);


assign rnx27onf2lbe = (l56q7o0hmnd98qc_ == 2'b0);

assign ntlp7re07dp6nkb = 
    (a94vd35etec4 | el7_p8jit09) & 
    (by_qc3yb1cyytd | fk5t4onucgv | lc6w646en ) 
    & rnx27onf2lbe
    ;

    
assign zijl1miri7deso9se = 
        
    af5qc04tmn51e4u2h1z & 
        
    a94vd35etec4 & 
        
    (by_qc3yb1cyytd | fk5t4onucgv | lc6w646en ) 
    ;

wire [4:0] pmwb1r70;
wire [2:0] anewxg;
wire [7:0] oev4182515 = {anewxg, pmwb1r70};
wire [64-1:0] k427ik6bety0vdf = {27'b0, pmwb1r70};
wire [64-1:0] bw8e1bo__j  = {29'b0, anewxg};
wire [64-1:0] g8cty956i = {24'b0, anewxg, pmwb1r70};

wire xdxa3krj224xup = by_qc3yb1cyytd & el7_p8jit09;
wire tv1zx6i5y5 = by_qc3yb1cyytd & a94vd35etec4;
wire hx6va8sy    = fk5t4onucgv    & el7_p8jit09;
wire bngdktf858    = fk5t4onucgv    & a94vd35etec4;
wire t1muoi2gjx2o   = lc6w646en   & el7_p8jit09;
wire i8ijh5v   = lc6w646en   & a94vd35etec4;

wire fhfnt0icr_sh = ((tv1zx6i5y5 | i8ijh5v) & izhvh9xxvwe2) | elspwgn4qhqqwg31epb;
wire [5-1:0] d08eosf2kx4k;

assign d08eosf2kx4k = elspwgn4qhqqwg31epb ? (pmwb1r70 | ciw6wwc7i33adp5) : vf5xcr67bqhzlo43_[4:0];
ux607_gnrl_dfflr #(5) fnvzwsmxfbb651 (fhfnt0icr_sh, d08eosf2kx4k, pmwb1r70, gf33atgy, ru_wi);

wire j2e56lmg = ((bngdktf858 | i8ijh5v) & izhvh9xxvwe2);
wire [3-1:0] tshg8iwoxx1;
assign tshg8iwoxx1 =  i8ijh5v ? vf5xcr67bqhzlo43_[7:5] : vf5xcr67bqhzlo43_[2:0];
ux607_gnrl_dfflr #(3) r3z7rgj6p_20b0 (j2e56lmg, tshg8iwoxx1, anewxg, gf33atgy, ru_wi);
assign phk590vi2 = anewxg;


wire o9ci7gemz = (e1go3iu == 12'h301);
wire tqmr31e = o9ci7gemz & el7_p8jit09;

wire [64-1:0] a1sjkc9c8 = {
    2'b10 
   ,36'b0 
   ,1'b0 
   ,1'b0 
   ,1'b0 
   ,1'b0 
   ,1'b0 
   ,1'b1 
   ,1'b0 
   ,1'b1 
   ,1'b0 
   ,1'b0 
   ,1'b1 
   ,1'b0 
   ,1'b0 
   ,1'b1 
   ,1'b0 
   ,1'b0 
   ,1'b0 
   ,1'b1 
   ,1'b0 
   ,1'b0 
   ,1'b1 
   ,1'b0 
   ,1'b1 
   ,1'b1 
   ,1'b0 
   ,1'b1 
                           };








wire [64-1:0] hnd2jesdfkehin = 64'h0001c607 ;
wire [64-1:0] uonsn384se50 = 64'h01000200;
wire [64-1:0] mvsg2qxdmt29ncr9   = v09gw6e6rfjf05qg;


wire m8rmfuha0pch8g = (e1go3iu == 12'hF11);
wire os_f3xrbfr2or   = (e1go3iu == 12'hF12);
wire kp2w957z1v    = (e1go3iu == 12'hF13);
wire b18orstady8x36yc   = (e1go3iu == 12'hF14);
wire pjwkxwhqy7i    = (e1go3iu == 12'hFFF);

wire swp0cfl7pff8oo4 = el7_p8jit09 & m8rmfuha0pch8g;
wire e1j7flhjhq   = el7_p8jit09 & os_f3xrbfr2or  ;
wire tcpea5afm7of    = el7_p8jit09 & kp2w957z1v   ;
wire owcdacpz2mm   = el7_p8jit09 & b18orstady8x36yc  ;
wire ofj_z8n6541s    = el7_p8jit09 & pjwkxwhqy7i   ;


wire [64-1:0] p744ug1jil846r8g6p;


y123rdlyxl0o jbuwvh36bagusf09ex6(
    .rb050tnl       (rb050tnl      ),
    .a94vd35etec4     (a94vd35etec4    ),
    .el7_p8jit09     (el7_p8jit09    ),
    .e1go3iu       (e1go3iu      ),
    .vf5xcr67bqhzlo43_  (vf5xcr67bqhzlo43_ ),
    .l9erxxpnphqd26vg9  (p744ug1jil846r8g6p ),
    .izhvh9xxvwe2  (izhvh9xxvwe2),
    .u2dvoyt5e7o_03z9z5(dfkhf0zzmeauwtqm3som),

    .pcr4upio7_tx37     (pcr4upio7_tx37   ), 
    .uzklqlncpqqm1rav  (uzklqlncpqqm1rav),
    .ortueunvnkx_l5m_j  (ortueunvnkx_l5m_j),
    .hwuhtb7ucto_utk56  (hwuhtb7ucto_utk56),
    .i1env2kmns7qvvuuc  (i1env2kmns7qvvuuc),
    .g3s3vpafvy3i  (g3s3vpafvy3i),

    .gf33atgy  (gf33atgy  ),
    .ru_wi(ru_wi)

  );







wire nxhwdm9t8elx18;

wire xstatus_typ_ena;
assign xstatus_typ_ena = 
       jlud6jeuxe0espga
     | rrujrlc85mhm 
     | nxhwdm9t8elx18;

wire [1:0] xstatus_typ_nxt;
assign xstatus_typ_nxt  = 

               jlud6jeuxe0espga ? ( 
                   ( {2{sf0uuehfhfa}} & 2'b10) |
                   ( {2{hvy2cpsp75f3 }} & 2'b01 ) |
                   ( {2{z35xlcc6bt4 }} & 2'b11 )  
               ) :
               rrujrlc85mhm ? a031mt59o9h2wubgw :
               nxhwdm9t8elx18 ? vf5xcr67bqhzlo43_[7:6] :
                  gg_wcrbxzhh0uqxd; 

ux607_gnrl_dfflr #(2) at0_vr77bps1ovn6qyxr (xstatus_typ_ena, xstatus_typ_nxt, gg_wcrbxzhh0uqxd, gf33atgy, ru_wi);





wire a_i3bk5s12rg205nvokeu  = xstatus_typ_ena  



    ;

wire [1:0] asn4gw8dnmbzq_13f  = 
    jlud6jeuxe0espga ? (gg_wcrbxzhh0uqxd) :
    rrujrlc85mhm ? 
                 (w3ouq_ntb6lrj_6yi ? a031mt59o9h2wubgw  : edu3vzxs7stp) :
    nxhwdm9t8elx18 ? vf5xcr67bqhzlo43_[9:8] :



                  a031mt59o9h2wubgw; 

ux607_gnrl_dfflr #(2) zsip0goxtrf5w67xkl_ry (a_i3bk5s12rg205nvokeu, asn4gw8dnmbzq_13f, a031mt59o9h2wubgw, gf33atgy, ru_wi);



wire zj201cydmy_kb = (e1go3iu == 12'h7c4);
wire l0o8bky903 = zj201cydmy_kb & el7_p8jit09;
wire z92r7e_2xsqqb = zj201cydmy_kb & a94vd35etec4;
assign nxhwdm9t8elx18 = (z92r7e_2xsqqb & izhvh9xxvwe2) ;

wire fgc4ur8_m02 = (e1go3iu == 12'h7c9);
wire t3h801u9ezg0 = fgc4ur8_m02 & el7_p8jit09;
wire et2o3t3aus = fgc4ur8_m02 & a94vd35etec4;

wire b08e4aju4yb2 = (et2o3t3aus & izhvh9xxvwe2) | xv08lot3vi9dag4vs0  
               | upp957fldz7r621ml4u  
      ;
wire [64-1:0] nq512rs3pix;
wire [64-1:0] k_vcb1pm_phhq7k3;
assign k_vcb1pm_phhq7k3[64-1:3] = {64-3{1'b0}};
assign k_vcb1pm_phhq7k3[3-1:0] = 
                   xv08lot3vi9dag4vs0 ? ew08uu2kn2p9e11s[3-1:0] :
               upp957fldz7r621ml4u ? t29y65qqvjjxvouca3[3-1:0] :
                   vf5xcr67bqhzlo43_[3-1:0];

ux607_gnrl_dfflr  #(64) ea_5qmjjbjdx0htzfk (b08e4aju4yb2, k_vcb1pm_phhq7k3, nq512rs3pix, gf33atgy, ru_wi);
wire [64-1:0] it8le0crf9kmfqe = nq512rs3pix;


wire d521va8_2d6_c7j = 1'b0;
wire gbj6z3zlspk3_b9 = d521va8_2d6_c7j & el7_p8jit09;
wire r9oprq6okq6cw3dy = d521va8_2d6_c7j & a94vd35etec4;

wire cahpjkfqfy47 = (r9oprq6okq6cw3dy & izhvh9xxvwe2) | if5jz8qk0aqefy3v35o  
               | upp957fldz7r621ml4u  
      ;
wire [64-1:0] pt98qdy_96o0gqe;
wire [64-1:0] xlc5y90reewgujpre;
assign xlc5y90reewgujpre[64-1:3] = {64-3{1'b0}};
assign xlc5y90reewgujpre[3-1:0] = 
                   if5jz8qk0aqefy3v35o ? mtc04rctrfyb[3-1:0] :
               upp957fldz7r621ml4u ? emggndeggdfff68dw0[3-1:0] :

                   3'b0;

ux607_gnrl_dfflr  #(64) h_8be3yonuo1k0pyc6 (cahpjkfqfy47, xlc5y90reewgujpre, pt98qdy_96o0gqe, gf33atgy, ru_wi);
wire [64-1:0] viqilm0l71xjf5c = pt98qdy_96o0gqe;


  wire yntlnjuskcdz_iu5n9b  = 1'b0;
  wire x5cvi1amnkl04ey7vf_lr = 1'b0;








































  wire be3et1xn2x24urf  = 1'b0;
  wire mbxd32lvzvlnq_307s = 1'b0;







wire [64-1:0] vbw35s4mu01jg4;

assign vbw35s4mu01jg4[64-1:10] = {(64-10){1'b0}}; 
assign vbw35s4mu01jg4[ 9: 8] = a031mt59o9h2wubgw; 
assign vbw35s4mu01jg4[ 7: 6] = gg_wcrbxzhh0uqxd;  
assign vbw35s4mu01jg4[    5] = mbxd32lvzvlnq_307s ;   
assign vbw35s4mu01jg4[    4] = be3et1xn2x24urf;   
assign vbw35s4mu01jg4[    3] = 1'b0;
assign vbw35s4mu01jg4[    2] = 1'b0;
assign vbw35s4mu01jg4[    1] = x5cvi1amnkl04ey7vf_lr;
assign vbw35s4mu01jg4[    0] = yntlnjuskcdz_iu5n9b; 

assign vyxop00ua6vr = vbw35s4mu01jg4;



wire bun2s3y6z8vtjyxjzr9;
wire wfndbkyoc1wc094vwehhutg5krtg;
wire ad6d6ex80to7t3vvnc69u3pmz;
wire maynsergszxlh4jomqhce5ahk;
wire [64-1:0] o02hm9vkepj5rucwrif;
wire cry3qyaqkl89ztcpeizdmn2fj;
wire eil4t6r56iactzfh4_drmg7xv;
wire oi73ilapk89bv0c9d4nvacia05brp;

pcw8e2c5o1b_8 ozh_rtrqsuqd_ljv(

  .aw82i964do(aw82i964do),
  .y8_gkxsfle(y8_gkxsfle),

  .pydatzxqqi     (pydatzxqqi     ),
  .zmwq3e9oijvo7d7(zmwq3e9oijvo7d7),

  .btwmhh91h50d5flgwx4o6pwu(btwmhh91h50d5flgwx4o6pwu),

  .rb050tnl       (rb050tnl      ),
  .a94vd35etec4     (a94vd35etec4    ),
  .el7_p8jit09     (el7_p8jit09    ),
  .e1go3iu       (e1go3iu      ),
  .izhvh9xxvwe2  (izhvh9xxvwe2 ),
  .vf5xcr67bqhzlo43_  (vf5xcr67bqhzlo43_ ),
  .l9erxxpnphqd26vg9  (o02hm9vkepj5rucwrif ),

  .u2dvoyt5e7o_03z9z5     (bun2s3y6z8vtjyxjzr9     ),
  .um1_bmln_sf2i4vzbya_(maynsergszxlh4jomqhce5ahk),
  .chjt9v0na3idosi9_0j5fe  (wfndbkyoc1wc094vwehhutg5krtg  ),
  .i72_qcuo70vljgkcb0fbj  (ad6d6ex80to7t3vvnc69u3pmz  ),
  .gjyhd0u2t3wy11drm07 (oi73ilapk89bv0c9d4nvacia05brp ),
  .an0s8c6hcabd901wob_8zo  (cry3qyaqkl89ztcpeizdmn2fj  ),
  .e280ym1w614qoep160njy  (eil4t6r56iactzfh4_drmg7xv  ),

  .ftp0juzjm2b587cyw5(ftp0juzjm2b587cyw5),
  .fw4r5i27mgu0_(xq63jpu81drai3h0),

  .ij_sgq3rtvw2  (ij_sgq3rtvw2),
  .k9jntnqwqp (k9jntnqwqp),


  .l0hrd_ubxbkay3zy8yz(l0hrd_ubxbkay3zy8yz),

  .dk2xhkj77a  (dk2xhkj77a  ),
  .gf33atgy  (gf33atgy  ),
  .ru_wi(ru_wi)
  );

  wire s36z1abpqp;


wire [64-1:0] aur5f30tjm74ynd  ;  
wire [64-1:0] vxt5pb8sxldtxqw  ;  
wire [64-1:0] p3kutuvsyvsd  ;  




wire [64-1:0] mj56s1rlw1lf7pkf2icn8d;
wire vadpkdaztv820a8kvwp0;
wire ikq8fffiwai0wlaxzs4xfv08i;
wire wjtx1c23l6psom27nm_gsj1ljb2;

wire eu5gus8kcfxe2bn_5jpy90jbl;
wire nug315vy7hnf899pgdpd2t7oh8;






wire [64-1:0] ik3qrttb23ath92pyzd0i = vf5xcr67bqhzlo43_;

hprqrck8t9y3rksec  pkmwivzpaon0pdxx(

  .x8rpm78rvvycis                     (x8rpm78rvvycis                     ),
  .canacnkc7zibtkn418i                (canacnkc7zibtkn418i                ),
  .bwbmafs1inesgjyn                     (bwbmafs1inesgjyn                     ), 
  .bkkiffh6ob85nh79doya_                (bkkiffh6ob85nh79doya_                ), 
  .qhqqh0lyehgtfop1tc                (qhqqh0lyehgtfop1tc                ), 

  .sxhicsqvufwfbnk0                     (sxhicsqvufwfbnk0                     ),
  .x03ux1utw4qem5kk3c                (x03ux1utw4qem5kk3c                ),
  .ydydp69z03wvr97                     (ydydp69z03wvr97                     ), 
  .pjic5x84bqxpvdduy4r2s                (pjic5x84bqxpvdduy4r2s                ), 
  .w5az87bw32r0tjbo0tdrv2ouvx           (w5az87bw32r0tjbo0tdrv2ouvx           ), 

  .vs6ryzcr0bwqs5so                  (vs6ryzcr0bwqs5so                  ), 
  .j25ub196dc_agl8oovaex4                 (j25ub196dc_agl8oovaex4                 ), 
  .pi2nokcm8qf7och7l4g                 (pi2nokcm8qf7och7l4g                 ), 
  .c0i0hs5tz64_ce5f0z                (c0i0hs5tz64_ce5f0z                ), 
  .dmzdczrqcueolg3dzufj_by5rmf           (dmzdczrqcueolg3dzufj_by5rmf           ), 
  .a1sqko6fok9qzpbtyuw0                (a1sqko6fok9qzpbtyuw0                ), 
  .bquohubxiv2rsayn62v                (bquohubxiv2rsayn62v                ), 
  .kqyojh1maxy0x834htg               (kqyojh1maxy0x834htg               ), 

  .fkuqlh34r                         (fkuqlh34r                         ),                  
  .ni01kj42oob2x                       (ni01kj42oob2x                       ),                  
  .ah8kjlmvnaxzbi                       (ah8kjlmvnaxzbi                       ),           
  .st2zalpx0uf                       (st2zalpx0uf                       ),           
  .rm1dxjejhq7dh3q5m                      (rm1dxjejhq7dh3q5m                      ),           
  .sxvvsxtbhyvt                        (sxvvsxtbhyvt                        ),           
  .hpk3eafyque5ubt_c62flnny             (hpk3eafyque5ubt_c62flnny             ),        
  .sfezv1xz2ghvo8pkt                    (sfezv1xz2ghvo8pkt                    ),              
  .vagaza053272juvmo59v8w20s             (vagaza053272juvmo59v8w20s             ),       
  .rzf45534z36ejq96260                 (rzf45534z36ejq96260                 ),       
  .frzfsbt7hp3n4aj3zvvumnh0s              (frzfsbt7hp3n4aj3zvvumnh0s              ),        
  .zkuxqezrmlhyyjjgx                   (zkuxqezrmlhyyjjgx                   ),             
  .u3h5tvu1g2q93141j9o                   (u3h5tvu1g2q93141j9o                   ),             
  .pjh0wad7t_5du3cync_0c             (pjh0wad7t_5du3cync_0c             ),                        
  .wmkgrgf631pbq                     (wmkgrgf631pbq                     ),
  .oyq1p3qa2iffjuqns0jkgg                 (oyq1p3qa2iffjuqns0jkgg                 ),
  .qjw2q0j88rjr42lautsqnca             (qjw2q0j88rjr42lautsqnca             ),        
  .imkm56ujne9v4m6n08w1yf5622          (imkm56ujne9v4m6n08w1yf5622          ),    
  .txk1r9aiq_7l2nkw101w_               (txk1r9aiq_7l2nkw101w_               ),         
  .ih4hmwugasiodbx5da9_40kx              (ih4hmwugasiodbx5da9_40kx              ),        
  .x5vjq7mshfwr0h3q514t7mhdt              (x5vjq7mshfwr0h3q514t7mhdt              ),        
  .qrxtk7e03100_uwkx73sg7              (qrxtk7e03100_uwkx73sg7              ),        
  .i7qiq2q9c6hbeful9qu9lb              (i7qiq2q9c6hbeful9qu9lb              ),         
  .yr0s3skqk7cdqflsrbsxg9znu              (yr0s3skqk7cdqflsrbsxg9znu              ),         
  .adqieke11qo0elfz93hlouwjc0        (adqieke11qo0elfz93hlouwjc0        ),   
  .w93gdpnnxuydy53eu0s9nxw7xdct7      (w93gdpnnxuydy53eu0s9nxw7xdct7      ), 

  .ldj4m511gvpu12mdu1_                (ldj4m511gvpu12mdu1_                ), 
  .sl5f3k5g9ln8_zvzr                 (sl5f3k5g9ln8_zvzr                 ), 
  
  .cn8o3075eju6dycby                    (cn8o3075eju6dycby                    ), 
  .zi39s8s7rmgo_lyocr_               (zi39s8s7rmgo_lyocr_               ), 
  .g1cek93tezrlyyt                   (g1cek93tezrlyyt                   ), 
  .i22z6k7eo0it77lz2                    (i22z6k7eo0it77lz2                    ), 
  .w2h8uh3l463qbgqmv                      (w2h8uh3l463qbgqmv                      ), 
  

  .lodtxdqjnwvx                      (aw82i964do                            ),
  .cbbcxlflqkqoklckuekt                 (rvr30vvllni                        ),
  .n37wgp2u95gc5b_                      (y8_gkxsfle                            ),
  .ewe_b1wv9zhrc8rc6hhr                 (z1cj655u31                        ),
  .z28w9as50xav1c2ms                      (pydatzxqqi                          ),

  
  
  
  
  
  .s6ypv533tdywrez9dra               (izhvh9xxvwe2                      ),
  .wtxn5hz27d1ke0cp5p                    (a94vd35etec4                         ),
  .z_g_9tmwi_9phwpm                    (el7_p8jit09                         ),
  .zy04ur_r6ibez7                    (e1go3iu                           ),
  .tpenqez_048wjs0mji00                   (ik3qrttb23ath92pyzd0i                 ),
  .wg_nk5anc77k66ap                   (mj56s1rlw1lf7pkf2icn8d                 ),

  
  .m9i5nb3fpl7i1c2f7aqnda5a             (vadpkdaztv820a8kvwp0               ),
  .o9n8q26y9zbsj6n3w7zzdgn_d7n90v        (ikq8fffiwai0wlaxzs4xfv08i          ),
  .fc8jy9eix4zbo26a2l3mebjykj99y         (wjtx1c23l6psom27nm_gsj1ljb2           ),
  
  .zds0n3s_2vya92r6p0iu18ede83st        (eu5gus8kcfxe2bn_5jpy90jbl          ),
  .j_oxbujpaq4zahlaf42l9paa_kjbrj         (nug315vy7hnf899pgdpd2t7oh8           ),
  

  .gf33atgy                               (gf33atgy                               ),
  .ru_wi                             (ru_wi                             )


); 













wire vybduk_04wdx6z05 = (e1go3iu == 12'h811);


wire z49s15yop6m7rk = (e1go3iu == 12'h812);


wire k9p_ach = (e1go3iu == 12'h810);


wire x4_1imazttasol8  = el7_p8jit09 & vybduk_04wdx6z05    ;
wire hyvne9dzw       = el7_p8jit09 & z49s15yop6m7rk      ;
wire wuiysx          = el7_p8jit09 & k9p_ach      ;

wire zu0202y516s22nuo0fu  = a94vd35etec4 & vybduk_04wdx6z05    ;
wire ns4gff9tzi8lp       = a94vd35etec4 & z49s15yop6m7rk      ;
wire n_0isc          = a94vd35etec4 & k9p_ach      ;

wire xmvyqncdiz9_fgtwn342gu = (zu0202y516s22nuo0fu & izhvh9xxvwe2);
wire j2w9u9key57ykiqt2x      = (ns4gff9tzi8lp & izhvh9xxvwe2);
wire pcoac761dde         = (n_0isc & izhvh9xxvwe2);

wire [64-1:0] tkireqj3hero_;




wire wkkv54425fme32iu92j = xmvyqncdiz9_fgtwn342gu;
wire dfel3kb_gu9h9mvskf8q = wkkv54425fme32iu92j;
wire [64-1:0] o_7hbum_bc5xi2qa84 = {{(64-1){1'b0}},vf5xcr67bqhzlo43_[0]};
ux607_gnrl_dfflr #(64) yw06nxmp2cljc9wo0xgp (dfel3kb_gu9h9mvskf8q, o_7hbum_bc5xi2qa84, tkireqj3hero_, gf33atgy, ru_wi);

wire [64-1:0] uwpy_1502jyu8_t80s = tkireqj3hero_;
assign apid0ys34zyekptw7un = dfel3kb_gu9h9mvskf8q ? o_7hbum_bc5xi2qa84[0] : tkireqj3hero_[0];


wire [64-1:0] nv3epbls00sd;
wire xa4r96hs2__hj = j2w9u9key57ykiqt2x;
wire q4ksemahqzpmvli = nv3epbls00sd[0];
wire c2535e1_v_l01 = xa4r96hs2__hj | q4ksemahqzpmvli;
wire [64-1:0] udk340ssoag = xa4r96hs2__hj ? {{(64-1){1'b0}},vf5xcr67bqhzlo43_[0]} : 64'b0;

ux607_gnrl_dfflr #(64) s96jvi7a168qodw (c2535e1_v_l01, udk340ssoag, nv3epbls00sd, dk2xhkj77a, ru_wi);

wire [64-1:0] luex1cs6x7sa = nv3epbls00sd;


wire [64-1:0] hvvja;




wire xrop0ye = pcoac761dde;
wire l7lfxwvv = xrop0ye;
wire [64-1:0] fm13fd3bf = {{(64-1){1'b0}},vf5xcr67bqhzlo43_[0]};
ux607_gnrl_dfflr #(64) sd4t0wopt5 (l7lfxwvv, fm13fd3bf, hvvja, gf33atgy, ru_wi);

wire [64-1:0] inyyxdi9 = hvvja;


assign habgbg2jn3qi = tkireqj3hero_[0];
assign dg4hzu_ = nv3epbls00sd[0];
assign h7fseh5_df0hbx = hvvja[0];


      
wire f8nehtdp4c9jo5      = (e1go3iu == 12'h801);
wire lsbmvjc19i       = el7_p8jit09 & f8nehtdp4c9jo5;
wire suugkehjg       = a94vd35etec4 & f8nehtdp4c9jo5;
wire uh968q3yy1y3mfj0ra   = (suugkehjg & izhvh9xxvwe2);

wire [64-1:0] odwh1hqyx;
wire kjxnjvbr8s21 = wj5ypo5k | uh968q3yy1y3mfj0ra;
wire j82xc354drsqol41hms = wj5ypo5k | (uh968q3yy1y3mfj0ra & vf5xcr67bqhzlo43_[0]);  
wire [64-1:0] r_r1xl5n6o = {{64-1{1'b0}},j82xc354drsqol41hms};

ux607_gnrl_dfflr #(64) nljos7gcbpktdwlg (kjxnjvbr8s21, r_r1xl5n6o, odwh1hqyx, dk2xhkj77a, ru_wi);

wire [64-1:0] ywq7zmowlccfib = odwh1hqyx;


      
wire doorarnn829tt      = (e1go3iu == 12'hCFE);
wire vzxftoy0       = el7_p8jit09 & doorarnn829tt;
wire xmyr5k0r       = a94vd35etec4 & doorarnn829tt;
wire rj241pj6vx01ji   = xmyr5k0r & izhvh9xxvwe2;

wire [64-1:0] sp98l516;
wire bmh25fw9uqo6 =   jlud6jeuxe0espga
                  | z2g63deibg1b1quqr
                  | rj241pj6vx01ji
                  ;
wire [64-1:0] ntuqkqf6w76s = 
                    rj241pj6vx01ji ? vf5xcr67bqhzlo43_ : 
                    ~ftp0juzjm2b587cyw5 ? 'd0 :    
                    vdr9fi9zwq ? 64'd4 : 64'd2;

ux607_gnrl_dfflr #(64) ya4o7axl5df (bmh25fw9uqo6, ntuqkqf6w76s, sp98l516, dk2xhkj77a, ru_wi);

wire [64-1:0] vgcvjr8adr = sp98l516;



      
wire vu_8rttl4p4      = (e1go3iu == 12'hCFF);
wire mxqvlgcks       = el7_p8jit09 & vu_8rttl4p4;
wire behqufdlpd5o       = a94vd35etec4 & vu_8rttl4p4;
wire d55it488ay8jj7   = (behqufdlpd5o & izhvh9xxvwe2);

wire [64-1:0] qgu3m0jd6;
wire q7tjmm7esbmjes = d55it488ay8jj7;
wire [64-1:0] xd9tn1v151f5 = vf5xcr67bqhzlo43_;

ux607_gnrl_dfflr #(64) czqr6bwnmhb80z (q7tjmm7esbmjes, xd9tn1v151f5, qgu3m0jd6, dk2xhkj77a, ru_wi);

wire [64-1:0] cdiut_mads8ok7 = qgu3m0jd6;











wire gfy9n09ir7q8zrpld19 = (e1go3iu == 12'h7d6);
wire b2uwf6iur0a5ek5x9   = (e1go3iu == 12'h7d7);
wire x06wm7qebv8ymb   = (e1go3iu == 12'h7d9);
wire y_nu4e3x8595566bl = (e1go3iu == 12'h7d8);
wire od1i6efig3fvtth = (e1go3iu == 12'h7da);
wire zo5qd8wbwszeiqaye = (e1go3iu == 12'h7db);
wire rmx1zc2nonjyho98zpr_ = (e1go3iu == 12'h7dc);


wire tc3f_x03mu_vagb8bx2 = 1'b0;
wire ye2xj3py3c5f_h_b8f = 1'b0;

wire fw0ba932spu6w15bn  = el7_p8jit09 & gfy9n09ir7q8zrpld19    ;
wire b8ao64rq4cnci    = el7_p8jit09 & b2uwf6iur0a5ek5x9      ;
wire pssagx292xg6    = el7_p8jit09 & x06wm7qebv8ymb      ;
wire pa1_agmr_3hhej4  = el7_p8jit09 & y_nu4e3x8595566bl    ;
wire djtm53o1_m_3x_4o  = el7_p8jit09 & od1i6efig3fvtth    ;
wire kxurpsnfj171m_n2_3aq  = el7_p8jit09 & zo5qd8wbwszeiqaye    ;
wire pu3hs090altkbczlh  = el7_p8jit09 & rmx1zc2nonjyho98zpr_    ;
wire b0g_t6oj33jh4lf_l55  = el7_p8jit09 & tc3f_x03mu_vagb8bx2    ;
wire hvopxeap8rqft0nnorg  = el7_p8jit09 & ye2xj3py3c5f_h_b8f    ;

wire d28tf6v6wgut0ci191  = izhvh9xxvwe2 & gfy9n09ir7q8zrpld19    ;
wire ehr2ha7t48r288ggw    = izhvh9xxvwe2 & b2uwf6iur0a5ek5x9      ;
wire w7ugv9ru4_u97fifzqp3j    = izhvh9xxvwe2 & x06wm7qebv8ymb      ;
wire m0438k2k0dc44z1u3pq  = izhvh9xxvwe2 & y_nu4e3x8595566bl    ;
wire daikhhsxmcnerj_4e80ivqi  = izhvh9xxvwe2 & od1i6efig3fvtth    ;
wire bb6j64jqgyjkhe9ncqe086e  = izhvh9xxvwe2 & zo5qd8wbwszeiqaye    ;
wire kaevo5afr0fflt_v5kx4t  = izhvh9xxvwe2 & rmx1zc2nonjyho98zpr_    ;
wire p7wisvtobgzr9fhglsey  = izhvh9xxvwe2 & tc3f_x03mu_vagb8bx2    ;
wire t784v6a773lmvnqsbpo_e4d2  = izhvh9xxvwe2 & ye2xj3py3c5f_h_b8f    ;

wire [64-1:0] ct4b0esmktg1; 
wire [64-1:0] gommhcpwq192s; 
wire [64-1:0] jh7p08bkr6ub0y6; 
wire [64-1:0] fckpj6qj1ryebu5; 





wire [1:0]     lpfne7pyt67tz6;
wire           cyibxvd3ybhq;
wire           x8fa6tqc4bod0tu;
wire [2:1]     zmuxspq81yu;
wire           pk2thujd8c_2p; 

wire [1:0]     ratz7ui0huis;
wire           lr2553eqc4;
wire           voslv77u0qi90;
wire [2:1]     lzl3ye9q;
wire           wqhz17z2xwv; 

wire [1:0]     bzacx6dk;
wire           c6abnw7v4_4;
wire           ajexu7adnd9k_z;
wire [2:1]     ahdlwplx;
wire           uw21ysgbvd; 

wire  p70o11vw5nzktjjjxh1e8q = (~hvy2cpsp75f3) & jlud6jeuxe0espga;

wire okih598qdw9bggn60e  = 
       p70o11vw5nzktjjjxh1e8q
     | upp957fldz7r621ml4u
     | d28tf6v6wgut0ci191
     ;

assign {
     lpfne7pyt67tz6,
     cyibxvd3ybhq,
     x8fa6tqc4bod0tu,
     zmuxspq81yu,
     pk2thujd8c_2p, 

     ratz7ui0huis,
     lr2553eqc4,
     voslv77u0qi90,
     lzl3ye9q,
     wqhz17z2xwv}  = 
    p70o11vw5nzktjjjxh1e8q ? {
                    edu3vzxs7stp,
                    idq_m7lglm,
                    r1u74u2bcei1,
                    rlsnapd43j6,
                    d63fiicib,

                    a031mt59o9h2wubgw,
                    mbxd32lvzvlnq_307s,
                    x5cvi1amnkl04ey7vf_lr,
                    dttzf_6vv87y,
                    d9w566umxhr1msc5h_ 
                    } :
    upp957fldz7r621ml4u ?  {
                    bzacx6dk, 
                    c6abnw7v4_4, 
                    ajexu7adnd9k_z, 
                    r1cznjd8rub5fb1xpx1,
                    1'b1,

                    bzacx6dk, 
                    c6abnw7v4_4, 
                    ajexu7adnd9k_z, 
                    ahdlwplx, 
                    uw21ysgbvd 
                    }:
                        
     d28tf6v6wgut0ci191 ? {
                    vf5xcr67bqhzlo43_[15:14] ,
                    vf5xcr67bqhzlo43_[13] ,
                    vf5xcr67bqhzlo43_[11] ,
                    vf5xcr67bqhzlo43_[10:9] ,
                    vf5xcr67bqhzlo43_[8] ,

                    vf5xcr67bqhzlo43_[7:6],  
                    vf5xcr67bqhzlo43_[5],  
                    vf5xcr67bqhzlo43_[3] , 
                    vf5xcr67bqhzlo43_[2:1] , 
                    vf5xcr67bqhzlo43_[0]   
                    }:
                    {
                    bzacx6dk,
                    c6abnw7v4_4,
                    ajexu7adnd9k_z,
                    ahdlwplx,
                    uw21ysgbvd,

                    edu3vzxs7stp,
                    idq_m7lglm,
                    r1u74u2bcei1,
                    rlsnapd43j6,
                    d63fiicib
                    }; 

ux607_gnrl_dfflr #(2) y8egsunxctbci1wl(okih598qdw9bggn60e, lpfne7pyt67tz6, bzacx6dk, gf33atgy, ru_wi);
ux607_gnrl_dfflr #(1) byg9e5k3xelkqhmuo(okih598qdw9bggn60e, x8fa6tqc4bod0tu, ajexu7adnd9k_z, gf33atgy, ru_wi);
ux607_gnrl_dfflr #(1) am4axwh59yhu (okih598qdw9bggn60e, cyibxvd3ybhq, c6abnw7v4_4, gf33atgy, ru_wi);

ux607_gnrl_dfflr #(2) ojue1suz6k6yylcn(okih598qdw9bggn60e, ratz7ui0huis, edu3vzxs7stp, gf33atgy, ru_wi);
ux607_gnrl_dfflr #(1) wx1utku479ecgi84s(okih598qdw9bggn60e, voslv77u0qi90, r1u74u2bcei1, gf33atgy, ru_wi);
ux607_gnrl_dfflr #(1) bul54kxy43zgq (okih598qdw9bggn60e, lr2553eqc4, idq_m7lglm, gf33atgy, ru_wi);

   
ux607_gnrl_dfflrs #(1) b28tnracmria5e (okih598qdw9bggn60e, pk2thujd8c_2p, uw21ysgbvd, gf33atgy, ru_wi);
ux607_gnrl_dfflrs #(1) zkion4htku3e (okih598qdw9bggn60e, wqhz17z2xwv, d63fiicib, gf33atgy, ru_wi);

              
ux607_gnrl_dfflr #(2) db2xnamtwxjye(okih598qdw9bggn60e, zmuxspq81yu, ahdlwplx, gf33atgy, ru_wi);
ux607_gnrl_dfflr #(2) dyck1n2tuk(okih598qdw9bggn60e, lzl3ye9q, rlsnapd43j6, gf33atgy, ru_wi);

wire [64-1:0] v0k9xrr0s5wwex3;

assign v0k9xrr0s5wwex3[64-1:16] = {(64-16){1'b0}};  

assign v0k9xrr0s5wwex3[15:14] = bzacx6dk  ;  
assign v0k9xrr0s5wwex3[13]    = c6abnw7v4_4  ;
assign v0k9xrr0s5wwex3[12]    = 1'b0;
assign v0k9xrr0s5wwex3[11]    = ajexu7adnd9k_z;
assign v0k9xrr0s5wwex3[10:9]  = ahdlwplx   ;
assign v0k9xrr0s5wwex3[8]     = uw21ysgbvd  ;
assign v0k9xrr0s5wwex3[7:6]   = edu3vzxs7stp  ;
assign v0k9xrr0s5wwex3[5]     = idq_m7lglm  ;
assign v0k9xrr0s5wwex3[4]     = 1'b0;
assign v0k9xrr0s5wwex3[3]     = r1u74u2bcei1;
assign v0k9xrr0s5wwex3[2:1]   = rlsnapd43j6   ;
assign v0k9xrr0s5wwex3[0]     = d63fiicib  ;

wire [64-1:0] jrvynb6nwm9au6qy;
wire [64-1:0] ftl2bjw_0egby88_x;
wire [64-1:0] z6bcw7fftmftvdx_fz5;
wire [64-1:0] i__roj_o_7vaojofud;

wire e8klq193tz8bh  = 
       p70o11vw5nzktjjjxh1e8q
     | upp957fldz7r621ml4u
     | ehr2ha7t48r288ggw
     ;

assign z6bcw7fftmftvdx_fz5 = 
    p70o11vw5nzktjjjxh1e8q ?  mzvpa_lx :
    upp957fldz7r621ml4u ?  ct4b0esmktg1:
    ehr2ha7t48r288ggw ?  vf5xcr67bqhzlo43_ : 
                    czcawgfux3h7; 

assign jrvynb6nwm9au6qy[64-1:1] = z6bcw7fftmftvdx_fz5[64-1:1];
assign jrvynb6nwm9au6qy[0] = 1'b0;

ux607_gnrl_dfflr #(64) m2r9gyaf563g8r0tpxn (e8klq193tz8bh, jrvynb6nwm9au6qy, czcawgfux3h7, gf33atgy, ru_wi);

wire g59sx7ygjymrrfl  = 
       p70o11vw5nzktjjjxh1e8q
     | upp957fldz7r621ml4u
     | w7ugv9ru4_u97fifzqp3j
     ;

assign i__roj_o_7vaojofud = 
    p70o11vw5nzktjjjxh1e8q ?  czcawgfux3h7 :
    upp957fldz7r621ml4u ?  ct4b0esmktg1:
    w7ugv9ru4_u97fifzqp3j ?  vf5xcr67bqhzlo43_ :
                    ct4b0esmktg1; 

assign ftl2bjw_0egby88_x[64-1:1] = i__roj_o_7vaojofud[64-1:1];
assign ftl2bjw_0egby88_x[0] = 1'b0;
ux607_gnrl_dfflr #(64) nupw_222y0ly1ww3jmw (g59sx7ygjymrrfl, ftl2bjw_0egby88_x, ct4b0esmktg1, gf33atgy, ru_wi);

wire [64-1:0] ff8pmmjdb0np9ipt;
wire [64-1:0] rro5qnhi8bh2hueyg;
wire [64-1:0] l5r5ynf5reoln1b;
wire [64-1:0] pn08q28r7f2a40n;
wire [64-1:0] dr4_6e1yettrndsbt7a;
wire [64-1:0] x0nnpdtngclw_i7ci066;

wire qc5z5nk1jbslemtxz  = 
       p70o11vw5nzktjjjxh1e8q
     | upp957fldz7r621ml4u
     | m0438k2k0dc44z1u3pq
     ;

wire [64-1:0] yvnhi6v8964pj92_f2 = 
    p70o11vw5nzktjjjxh1e8q ?  cause_r :
    upp957fldz7r621ml4u ?  gommhcpwq192s:
    m0438k2k0dc44z1u3pq ?  vf5xcr67bqhzlo43_ :
                    qxyauqoyrj6kj; 


wire gcjjzvv_nuaq_4  = 
       p70o11vw5nzktjjjxh1e8q
     | upp957fldz7r621ml4u
     | daikhhsxmcnerj_4e80ivqi
     ;

wire [64-1:0] ca4msfd36ycj6_4u0huy = 
    p70o11vw5nzktjjjxh1e8q ?  qxyauqoyrj6kj :
    upp957fldz7r621ml4u ?  gommhcpwq192s:
    daikhhsxmcnerj_4e80ivqi ?  vf5xcr67bqhzlo43_ :
                    gommhcpwq192s; 


    
    
    
    
    
    
    


assign ff8pmmjdb0np9ipt[64-2:31] = {(64-32){1'b0}};
assign ff8pmmjdb0np9ipt[64-1] = yvnhi6v8964pj92_f2[64-1];
assign ff8pmmjdb0np9ipt[30:27]   = yvnhi6v8964pj92_f2[30:27]; 
assign ff8pmmjdb0np9ipt[26:24]   = 3'b0;
assign ff8pmmjdb0np9ipt[23:16]   = yvnhi6v8964pj92_f2[23:16]; 
assign ff8pmmjdb0np9ipt[15:ob0j3iecn59nr6s8ur] = {(16-ob0j3iecn59nr6s8ur){1'b0}};
assign ff8pmmjdb0np9ipt[ob0j3iecn59nr6s8ur-1:0]   = yvnhi6v8964pj92_f2[ob0j3iecn59nr6s8ur-1:0]; 

assign rro5qnhi8bh2hueyg[64-2:31] = {(64-32){1'b0}};
assign rro5qnhi8bh2hueyg[64-1] = ca4msfd36ycj6_4u0huy[64-1];
assign rro5qnhi8bh2hueyg[30:27]   = ca4msfd36ycj6_4u0huy[30:27]; 
assign rro5qnhi8bh2hueyg[26:24]   = 3'b0;
assign rro5qnhi8bh2hueyg[23:16]   = ca4msfd36ycj6_4u0huy[23:16]; 
assign rro5qnhi8bh2hueyg[15:ob0j3iecn59nr6s8ur] = {(16-ob0j3iecn59nr6s8ur){1'b0}};
assign rro5qnhi8bh2hueyg[ob0j3iecn59nr6s8ur-1:0]   = ca4msfd36ycj6_4u0huy[ob0j3iecn59nr6s8ur-1:0]; 


ux607_gnrl_dfflr #(64) xf3tgqf6ahng519eczp (qc5z5nk1jbslemtxz, ff8pmmjdb0np9ipt, qxyauqoyrj6kj, gf33atgy, ru_wi);
ux607_gnrl_dfflr #(64) k3swk6ftnqbxvdfmlyo7y (gcjjzvv_nuaq_4, rro5qnhi8bh2hueyg, gommhcpwq192s, gf33atgy, ru_wi);

wire sl4u3ym2f7n5zri3  = 
       p70o11vw5nzktjjjxh1e8q
     | upp957fldz7r621ml4u
     | bb6j64jqgyjkhe9ncqe086e
     ;

wire [64-1:0] gqap4hc5hxhdb8tux3r = 
    p70o11vw5nzktjjjxh1e8q ?  nq512rs3pix :
    upp957fldz7r621ml4u ?  jh7p08bkr6ub0y6:
    bb6j64jqgyjkhe9ncqe086e ?  vf5xcr67bqhzlo43_ :
                    t29y65qqvjjxvouca3; 


wire kvaqqoo5f3wds76pn  = 
       p70o11vw5nzktjjjxh1e8q
     | upp957fldz7r621ml4u
     | kaevo5afr0fflt_v5kx4t
     ;

wire [64-1:0] kebewvcsk52j1txhtae2z0oz = 
    p70o11vw5nzktjjjxh1e8q ?  t29y65qqvjjxvouca3 :
    upp957fldz7r621ml4u ?  jh7p08bkr6ub0y6:
    kaevo5afr0fflt_v5kx4t ?  vf5xcr67bqhzlo43_ :
                    jh7p08bkr6ub0y6; 

assign l5r5ynf5reoln1b[64-1:3] = {64-3{1'b0}};
assign l5r5ynf5reoln1b[3-1:0]  = gqap4hc5hxhdb8tux3r[3-1:0];

assign pn08q28r7f2a40n[64-1:3] = {64-3{1'b0}};
assign pn08q28r7f2a40n[3-1:0]  = kebewvcsk52j1txhtae2z0oz[3-1:0];

ux607_gnrl_dfflr #(64) sjn0d2kxvpgchgs6tnkfp (sl4u3ym2f7n5zri3, l5r5ynf5reoln1b, t29y65qqvjjxvouca3, gf33atgy, ru_wi);
ux607_gnrl_dfflr #(64) ptkfb13zy9hytc_iih (kvaqqoo5f3wds76pn, pn08q28r7f2a40n, jh7p08bkr6ub0y6, gf33atgy, ru_wi);

wire ewafuhl7_38m2pahx  = 
       p70o11vw5nzktjjjxh1e8q
     | upp957fldz7r621ml4u
     | p7wisvtobgzr9fhglsey
     ;

wire [64-1:0] binf7qexd2mm509c0_kg = 
    p70o11vw5nzktjjjxh1e8q ?  pt98qdy_96o0gqe :
    upp957fldz7r621ml4u ?  fckpj6qj1ryebu5:
    
    p7wisvtobgzr9fhglsey ?  64'b0 :
                    emggndeggdfff68dw0; 


wire osp3gc4ntjcj2f6zu827  = 
       p70o11vw5nzktjjjxh1e8q
     | upp957fldz7r621ml4u
     | t784v6a773lmvnqsbpo_e4d2
     ;

wire [64-1:0] y1w5yntfe9czo780c22zypg = 
    p70o11vw5nzktjjjxh1e8q ?  emggndeggdfff68dw0 :
    upp957fldz7r621ml4u ?  fckpj6qj1ryebu5:
    
    t784v6a773lmvnqsbpo_e4d2 ? 64'b0   :
                    fckpj6qj1ryebu5; 

assign dr4_6e1yettrndsbt7a[64-1:5] = {64-5{1'b0}};
assign dr4_6e1yettrndsbt7a[5-1:0]  = binf7qexd2mm509c0_kg[5-1:0];

assign x0nnpdtngclw_i7ci066[64-1:5] = {64-5{1'b0}};
assign x0nnpdtngclw_i7ci066[5-1:0]  = y1w5yntfe9czo780c22zypg[5-1:0];

ux607_gnrl_dfflr #(64) l7k41f21lupcg1nr8jfvk_m (ewafuhl7_38m2pahx, dr4_6e1yettrndsbt7a, emggndeggdfff68dw0, gf33atgy, ru_wi);
ux607_gnrl_dfflr #(64) vpg1jga391ljotl_kwi (osp3gc4ntjcj2f6zu827, x0nnpdtngclw_i7ci066, fckpj6qj1ryebu5, gf33atgy, ru_wi);


wire [64-1:0] wsr5asmu2rsl6a076 = czcawgfux3h7; 
wire [64-1:0] pealk1ny1w3zypaet = ct4b0esmktg1; 
wire [64-1:0] oxqig8tg9r_4az4sf = qxyauqoyrj6kj; 
wire [64-1:0] clr_f9f2zh_fkkespze = gommhcpwq192s; 
wire [64-1:0] t_7nv9a3lsvuzxmcw = t29y65qqvjjxvouca3; 
wire [64-1:0] bqp1xynoo31eoavfit1 = jh7p08bkr6ub0y6; 
wire [64-1:0] rziri8ijn84w3o8cp = emggndeggdfff68dw0; 
wire [64-1:0] f36cakmqdwzxjjajghlg = fckpj6qj1ryebu5; 









wire jjvcrtzj366t   = (e1go3iu == 12'hfc0);
wire a06ag5mfqc7b   = (e1go3iu == 12'hfc1);
wire skog6xw8aj1km8ost   = (e1go3iu == 12'hfc2);
wire ad2bzpfqdx      = (e1go3iu == 12'h7c0);
wire veysvh0g_5rkx      = (e1go3iu == 12'h7c1);
wire andomkgjr      = (e1go3iu == 12'h7f0);
wire wefdo3j2oa      = (e1go3iu == 12'h7f1);
assign sim0gblc86voze3mam = (e1go3iu == 12'h7ca);
assign wft1k16f78xw2  = (e1go3iu == 12'h7d0);

wire zmgxfaohma89cv5    = el7_p8jit09 & jjvcrtzj366t     ;
wire l7r01a30uiu    = el7_p8jit09 & a06ag5mfqc7b     ;
wire noizhmz52v5iwfm    = el7_p8jit09 & skog6xw8aj1km8ost     ;
wire k1j9zf14hj       = el7_p8jit09 & ad2bzpfqdx        ;
wire n4vaq5qq96wr       = el7_p8jit09 & veysvh0g_5rkx        ;
wire rvkrf8rv4n       = el7_p8jit09 & andomkgjr        ;
wire ydeihiywm       = el7_p8jit09 & wefdo3j2oa        ;
wire n1zvf0y1dwpep  = el7_p8jit09 & sim0gblc86voze3mam   ;
wire aaa3cgvzwhecdc46s   = el7_p8jit09 & wft1k16f78xw2    ;

wire w0huy5l6o9y8h      = izhvh9xxvwe2 & ad2bzpfqdx        ;
wire ux0qwuvuvrefd57r      = izhvh9xxvwe2 & veysvh0g_5rkx        ;


wire j1mr0hvfc5jpcnsoxt = izhvh9xxvwe2 & sim0gblc86voze3mam   ;
wire c824j4y2hi7huhtrq  = izhvh9xxvwe2 & wft1k16f78xw2    ;

wire [64-1:0] exmn1blzuoj779;  
wire [64-1:0] lz2fvl6kd9hk6v;  
wire [64-1:0] dalvbjr5v1ubv5s;  

wire [64-1:0] u86s55pt;     
wire [64-1:0] s7rqtmyt3;     
wire [64-1:0] h5pilu9pman;     
wire [64-1:0] ynzhbk4inf;     
wire [64-1:0] gq9vjo4xdonfw; 
























































































  
  
  
  
  localparam yap91qk_7w8isg6wcdjkyvwa6ip = (7 - 3);

assign exmn1blzuoj779[3:0] = yap91qk_7w8isg6wcdjkyvwa6ip[3:0];

  
assign exmn1blzuoj779[6:4] = 
                       3'd1;
                  
  
  
  
assign exmn1blzuoj779[9:7] = 3'd3;

assign exmn1blzuoj779[15:10] = 6'b0;


  
  
  
  
  localparam b9vmqo1964xsuc4qlaf7 = (16 - 7);
assign exmn1blzuoj779[20:16] = b9vmqo1964xsuc4qlaf7[4:0];



assign exmn1blzuoj779[21] = 1'b0;


assign exmn1blzuoj779[64-1:22] = {64-22{1'b0}};





















































  
  
  
  
  localparam x7sf_ikvk9begv1bhvk = (6 - 3);
assign lz2fvl6kd9hk6v[3:0] = x7sf_ikvk9begv1bhvk[3:0];

  
assign lz2fvl6kd9hk6v[6:4] = 
                       3'd1;
                  
  
  
  
assign lz2fvl6kd9hk6v[9:7] = 3'd3;
assign lz2fvl6kd9hk6v[15:10] = 6'b0;



  
  
  
  
  localparam akx7tq_cq5f4fux_0a3 = (16 - 7);
assign lz2fvl6kd9hk6v[20:16] = akx7tq_cq5f4fux_0a3[4:0];

assign lz2fvl6kd9hk6v[64-1:21] = {64-21{1'b0}};


























































































































assign dalvbjr5v1ubv5s[0] = 
                          1'b0;
assign dalvbjr5v1ubv5s[1] = 
                          1'b0;
assign dalvbjr5v1ubv5s[2] = 
                          1'b1;
assign dalvbjr5v1ubv5s[3] = 
                          1'b1;
assign dalvbjr5v1ubv5s[4] = 
                          1'b0;
assign dalvbjr5v1ubv5s[5] = 
                          1'b1;
assign dalvbjr5v1ubv5s[6] = 
                          1'b0;
assign dalvbjr5v1ubv5s[7] = 
                          1'b1;
assign dalvbjr5v1ubv5s[8] = 
                          1'b1;
assign dalvbjr5v1ubv5s[9] = 
                          1'b1;
assign dalvbjr5v1ubv5s[10] = 
                          1'b1;

assign dalvbjr5v1ubv5s[64-1:11] = {64-11{1'b0}};


ux607_gnrl_dfflrs #1 kcef52gdx0720f (w0huy5l6o9y8h, vf5xcr67bqhzlo43_[0], u86s55pt[0], gf33atgy, ru_wi);

assign u86s55pt[9:1] = 9'b0;

localparam bfe8r_4hym5e4k = 32'h80000000;
assign u86s55pt[64-1:10] =  {{64-32{1'b0}},bfe8r_4hym5e4k[32-1:10]};


ux607_gnrl_dfflrs #1 zp38b9ydpac1d (ux0qwuvuvrefd57r, vf5xcr67bqhzlo43_[0], s7rqtmyt3[0], gf33atgy, ru_wi);

assign s7rqtmyt3[9:1] = 9'b0;

localparam ygsl88a_l_hqz9y1 = 32'h90000000;
assign s7rqtmyt3[64-1:10] = {{64-32{1'b0}},ygsl88a_l_hqz9y1[32-1:10]};

assign w92a5o09fp9dg6 = u86s55pt[0];
assign eglor15f7p2ivpny5dc = s7rqtmyt3[0];

assign h5pilu9pman[0] = 1'b1;
  
  
  
  localparam po27sb8b_9aadq96po7 = (20 - 9);
assign h5pilu9pman[5:1] = po27sb8b_9aadq96po7[4:0];
assign h5pilu9pman[9:6] = 4'b0;

localparam xiiok7kjgjsa62nr4 = 32'h10000000;
assign h5pilu9pman[64-1:10] = {{64-32{1'b0}},xiiok7kjgjsa62nr4[32-1:10]};

assign ynzhbk4inf[64-1:0] = 64'b0;

wire [64-1:0] jna8pdej27pvms1;
wire yj29etiue6_lit = j1mr0hvfc5jpcnsoxt;
wire [64-1:0] ek9pjlslchx9kci8l7;
assign ek9pjlslchx9kci8l7[0] = vf5xcr67bqhzlo43_[0];
assign ek9pjlslchx9kci8l7[15:1] = 15'b0;
assign ek9pjlslchx9kci8l7[16] = vf5xcr67bqhzlo43_[16];
assign ek9pjlslchx9kci8l7[64-1:17] = {64-17{1'b0}};

ux607_gnrl_dfflr #(64) b8c7uxhyc3__vpsiay (yj29etiue6_lit, ek9pjlslchx9kci8l7, jna8pdej27pvms1, gf33atgy, ru_wi);

assign ous_emkpecrqhg5e7 = jna8pdej27pvms1[0];


assign doh50j3p7c7yl7uk9 = jna8pdej27pvms1[16];

wire s_hrrjehjigdw3pyc7 = c824j4y2hi7huhtrq;
wire [64-1:0] ep7d1zp90qxkm0;

assign ep7d1zp90qxkm0[64-1:10] = {(64-10){1'b0}};
assign gq9vjo4xdonfw[64-1:10] = {(64-10){1'b0}};

assign ep7d1zp90qxkm0[9] = vf5xcr67bqhzlo43_[9];
ux607_gnrl_dfflr #(1) c9k70p51f8uzk18zk1 (s_hrrjehjigdw3pyc7, ep7d1zp90qxkm0[9], gq9vjo4xdonfw[9], gf33atgy, ru_wi);

assign w2fpnf5fg1byp6 = gq9vjo4xdonfw[9];

assign ep7d1zp90qxkm0[8:7] = 2'b0;
assign gq9vjo4xdonfw[8:7] = 2'b0;

assign ep7d1zp90qxkm0[5:4] = 2'b0;
assign gq9vjo4xdonfw[5:4] = 2'b0;


assign ep7d1zp90qxkm0[2] = 1'b0;

assign ep7d1zp90qxkm0[1:0] = 2'b0;
assign gq9vjo4xdonfw[1:0] = 2'b0;

assign ep7d1zp90qxkm0[6] = vf5xcr67bqhzlo43_[6];
ux607_gnrl_dfflrs #(1) zng6iz8v748hw3r0dksw (s_hrrjehjigdw3pyc7, ep7d1zp90qxkm0[6], gq9vjo4xdonfw[6], gf33atgy, ru_wi);
assign exltui35irvvmodu205vw = gq9vjo4xdonfw[6];


assign ep7d1zp90qxkm0[3] = vf5xcr67bqhzlo43_[3];
ux607_gnrl_dfflrs #(1) dzt48khd0xm5wo6e7kw1 (s_hrrjehjigdw3pyc7, ep7d1zp90qxkm0[3], gq9vjo4xdonfw[3], gf33atgy, ru_wi);
assign s7eq8f6z1uyi2in = gq9vjo4xdonfw[3];


ux607_gnrl_dfflr  #(1) ajan31fzj51ulu7n18r7  (s_hrrjehjigdw3pyc7, ep7d1zp90qxkm0[2], gq9vjo4xdonfw[2], gf33atgy, ru_wi);



assign qbsr1jytrqtsbk4ttb8nz = gq9vjo4xdonfw[2];




assign aur5f30tjm74ynd   = exmn1blzuoj779  ; 
assign vxt5pb8sxldtxqw   = lz2fvl6kd9hk6v  ;
assign p3kutuvsyvsd   = dalvbjr5v1ubv5s  ;
wire [64-1:0] ove0jfc9_      = u86s55pt     ;
wire [64-1:0] ae1hd9imgwd      = s7rqtmyt3     ;
wire [64-1:0] b0en4jlm5ni5      = h5pilu9pman     ;
wire [64-1:0] arakgrjva32d      = ynzhbk4inf     ;
wire [64-1:0] htdx5bpibi4z9nvhfcy = jna8pdej27pvms1;
wire [64-1:0] epnwm13_bdyvjd  = gq9vjo4xdonfw ;


wire [64-1:0] skijzqww3h5f0m4sa60i5v = 64'h112;
wire [64-1:0] juemut6ntjn4jv9_j6mivuv = 64'h211;
wire [64-1:0] bl_mgp0p3lt5qt52uv9 = 64'h211;
wire [64-1:0] hkvtut3x96fj_tl = (skijzqww3h5f0m4sa60i5v + juemut6ntjn4jv9_j6mivuv + bl_mgp0p3lt5qt52uv9);



wire [64-1:0] qyirue3_ioqbr = 64'h8b9746fc;







wire il_e54l8ycmz2u;
wire bd9vwvml7qb;

wire qb5qu1p3;
wire myuno7j;
wire hil0xjb;
wire mdssp2oy8dtr0s;
wire qtf8of_u5z5iai;
wire ed9vgeh97yj;
wire yl_l2gn_qt7p7;
wire kiky8rqvpf1zkvtf;
wire ja2k8c_59wnmay5l;
wire ng7hgd38lorxo;
wire eo9lmvnadbu765;
wire tf6c6wjqdv5vvu4;
wire b4etkbmloh;
wire ven2nsl;
wire zy44s2bwza9;
wire m4xr4juqkq;
wire no4tukpi8i35;
wire elq67c0en7exei;
wire fzwoxh5vqm8;
wire syf4axzj9zyr;
wire xrbzeq_xg1z9;
wire e364tfszybtw35;
wire h9bg0vmhmf;
wire ls416x5_x21tvc;
wire d1bjdianldviz8;
wire e3t8l4w0xlvk50p;
wire bh9_1u0btegoxnhc_;
wire rmh20fa2i1zgb;
wire wy0jv5w_isf0qmqb;
wire pyczk46mr25dxfykg;
wire ha7fcf0ap;
wire uz6ke_lem;
wire ano1d1_31;
wire kkco_owc1;
wire dk878usgx2r;
wire vcsyiox9w;
wire lqzw29rbc73ulx;
wire ddx7351w3ukkafuh3;
wire rjju_oexoi2ozf1eo;
wire ymnk8i8eh3n9_ib7224;
wire hze_3v_qjwxi4mrbnkcnic;



assign iiq92rsh_v1ylb = (e1go3iu == 12'h100);
assign il_e54l8ycmz2u = iiq92rsh_v1ylb & el7_p8jit09;
assign bd9vwvml7qb = iiq92rsh_v1ylb & a94vd35etec4;
assign b3lm_1ct7augo = bd9vwvml7qb & izhvh9xxvwe2;


wire f4_gpy7hep0c0klauu;
wire h3i6eb2cvw_u0sk_9ap9 = 
                         f4_gpy7hep0c0klauu   
                       | z2g63deibg1b1quqr       
                       | s_m3pbf5m2tr6v
                       | b3lm_1ct7augo 
                       | to3k3giu627wb2b7yd 
                       ;

wire uy_j_dcfffe0;
wire ty64g8m1v81v7625;
wire tgbuoad1ggbbyep9jj = 
                        f4_gpy7hep0c0klauu ? (
                        uy_j_dcfffe0 ? 1'b1 :
                        bj7h5jqg66r51jxki6emra[1]) :  
    
    
    
    
    
                        z2g63deibg1b1quqr ? 1'b0 :
    
    
    
    
                        s_m3pbf5m2tr6v ? ty64g8m1v81v7625 :
    
                        b3lm_1ct7augo ? vf5xcr67bqhzlo43_[1] : 
    
                        to3k3giu627wb2b7yd ? vf5xcr67bqhzlo43_[1] : 
                        w632tcbtqncn6; 

ux607_gnrl_dfflr #(1) t2vdw4z0jhefqknpkp (h3i6eb2cvw_u0sk_9ap9, tgbuoad1ggbbyep9jj, w632tcbtqncn6, gf33atgy, ru_wi);



wire xu0fn1yd6ygtq_mfki4dzag = syf4axzj9zyr & dn8riluj40uunvq5;
wire xyue7r6hcp92wroepjp  = 
       z2g63deibg1b1quqr
     | s_m3pbf5m2tr6v 
     | xu0fn1yd6ygtq_mfki4dzag   
     | b3lm_1ct7augo
     | to3k3giu627wb2b7yd;

wire z68n7_ywkx_w9h75_f8    = 
    
    
    
    
                           z2g63deibg1b1quqr ? w632tcbtqncn6 :
    
    
    
    
    
                           s_m3pbf5m2tr6v  ? 
    
    
    
                           1'b1 :
    
    
                           b3lm_1ct7augo ? vf5xcr67bqhzlo43_[5] : 
    
                           to3k3giu627wb2b7yd ? vf5xcr67bqhzlo43_[5] : 
                           xu0fn1yd6ygtq_mfki4dzag  ?  vf5xcr67bqhzlo43_[27]:
                           ty64g8m1v81v7625; 
ux607_gnrl_dfflr #(1) qdv46qi2i4k3j2ygkp (xyue7r6hcp92wroepjp, z68n7_ywkx_w9h75_f8, ty64g8m1v81v7625, gf33atgy, ru_wi);


wire t9kr9mnvt6dgqdy = xyue7r6hcp92wroepjp;

wire io722b8lft61t4i4qf;

wire osdmvzo4uwr9pncckow = 1'b0;   
assign io722b8lft61t4i4qf = 
    
                z2g63deibg1b1quqr ? status_priv_r[0] : 
    
    
                s_m3pbf5m2tr6v ? 



                                  osdmvzo4uwr9pncckow :

    
                to3k3giu627wb2b7yd ? vf5xcr67bqhzlo43_[8] :
                b3lm_1ct7augo ? vf5xcr67bqhzlo43_[8] :
                xu0fn1yd6ygtq_mfki4dzag ?  uiulkx67fwpf7in8sde_kj[28] : 
                                ogmro605vz43jd_a6;

ux607_gnrl_dfflr #(1) f_sxefqwl22acwufph7e (t9kr9mnvt6dgqdy, io722b8lft61t4i4qf, ogmro605vz43jd_a6, gf33atgy, ru_wi);


wire q16znjqn1kyhkskoei8 = b3lm_1ct7augo | to3k3giu627wb2b7yd;

wire fg008o985ioh4pzxat;
wire m795w3j_3yxa2b;

assign fg008o985ioh4pzxat =   1'b0
                         | vf5xcr67bqhzlo43_[18] 
                         ;

ux607_gnrl_dfflr #(1) wm30b71f_88p66bgip (q16znjqn1kyhkskoei8, fg008o985ioh4pzxat, m795w3j_3yxa2b, gf33atgy, ru_wi);



wire r50jn2fllskmnayjdfum = b3lm_1ct7augo | to3k3giu627wb2b7yd;

wire nml5xap0t4llynz;
wire tsa6ms1s2xk2ql;

assign nml5xap0t4llynz = vf5xcr67bqhzlo43_[19];

ux607_gnrl_dfflr #(1) p9p80bgqt4a6pf7j_7 (r50jn2fllskmnayjdfum, nml5xap0t4llynz, tsa6ms1s2xk2ql, gf33atgy, ru_wi);

wire jzukd13j0mn1 = tsa6ms1s2xk2ql;

assign csr_sstatus[64-1] = d6z8hz6u7gym;                 
assign csr_sstatus[64-2:36] = 27'b0;
assign csr_sstatus[35:34] = 2'b0;
assign csr_sstatus[33:32] = nriqmhgyl2409;
assign csr_sstatus[31]    = 1'b0; 

assign csr_sstatus[30:23] = 8'b0;                               
assign csr_sstatus[22:20] = 3'b0;                               
assign csr_sstatus[19]    = tsa6ms1s2xk2ql;                      
assign csr_sstatus[18]    = m795w3j_3yxa2b;                      
assign csr_sstatus[17]    = 1'b0;                               
assign csr_sstatus[16:15] = i8uou0fe4qb;                        
assign csr_sstatus[14:13] = l56q7o0hmnd98qc_;                        
assign csr_sstatus[12:9]  = 4'b0;
assign csr_sstatus[8]     = ogmro605vz43jd_a6;
assign csr_sstatus[7:6]   = 2'b0;
assign csr_sstatus[5]     = ty64g8m1v81v7625;
assign csr_sstatus[4]     = 1'b0;
assign csr_sstatus[3:2]   = 2'b0;
assign csr_sstatus[1]     = w632tcbtqncn6; 
assign csr_sstatus[0]     = 1'b0; 

wire arxwb4avzd = ogmro605vz43jd_a6; 
assign lhu2z948o3n = arxwb4avzd;















assign qb5qu1p3 = (e1go3iu == 12'h104);
assign myuno7j = qb5qu1p3 & el7_p8jit09;
assign hil0xjb = qb5qu1p3 & a94vd35etec4;
assign mdssp2oy8dtr0s = (~dn8riluj40uunvq5) & hil0xjb & izhvh9xxvwe2; 
wire u7s_j2xak2h = yw2rjoyrops;
wire ky0wefrd_hy = 
                 mdssp2oy8dtr0s
               | u7s_j2xak2h
               ;
wire [64-1:0] y0o55;
wire [64-1:0] zr5sc2vs;

assign zr5sc2vs[64-1:22] = {(64-22){1'b0}};
assign zr5sc2vs[21] = 1'b0;
assign zr5sc2vs[20] = 1'b0;
assign zr5sc2vs[19] = 1'b0;
assign zr5sc2vs[18] = 1'b0;
assign zr5sc2vs[17] = 1'b0;
assign zr5sc2vs[16] = 1'b0;












assign zr5sc2vs[15:10] = 6'b0;
assign zr5sc2vs[9] = 
    
                     mdssp2oy8dtr0s ? vf5xcr67bqhzlo43_[9] :   
    
                     u7s_j2xak2h ? vf5xcr67bqhzlo43_[9] :   
                     y0o55[9]; 
assign zr5sc2vs[8:6] = 3'b0;
assign zr5sc2vs[ 5] = 
    
                     mdssp2oy8dtr0s ? vf5xcr67bqhzlo43_[5] :   
    
                     u7s_j2xak2h ? vf5xcr67bqhzlo43_[5] :   
                     y0o55[5]; 
assign zr5sc2vs[4:2] = 3'b0;
assign zr5sc2vs[ 1] = 
    
                     mdssp2oy8dtr0s ? vf5xcr67bqhzlo43_[1] :   
    
                     u7s_j2xak2h ? vf5xcr67bqhzlo43_[1] :   
                     y0o55[1]; 
assign zr5sc2vs[0] = 1'b0;
ux607_gnrl_dfflr #(64) o2jmc146x (ky0wefrd_hy, zr5sc2vs, y0o55, gf33atgy, ru_wi);
assign csr_sie = dn8riluj40uunvq5 ? 32'b0 : y0o55;
assign ai169tbqp4seb3 = csr_sie[ 9];
assign b0zz_ornhz010 = csr_sie[ 5];
assign yw4o4kdms07_32 = csr_sie[ 1];
 


assign qtf8of_u5z5iai = (e1go3iu == 12'h105);
assign ed9vgeh97yj = el7_p8jit09 & qtf8of_u5z5iai;
assign yl_l2gn_qt7p7 = qtf8of_u5z5iai & a94vd35etec4;
assign kiky8rqvpf1zkvtf= yl_l2gn_qt7p7 & izhvh9xxvwe2;
wire enjb050zotyx23 = kiky8rqvpf1zkvtf;
wire [64-1:0] a82ka7y2g;
wire [64-1:0] n51bu0uh_wb51w = vf5xcr67bqhzlo43_[64-1:0];
ux607_gnrl_dfflr #(64) p70h4qjkrnk (enjb050zotyx23, n51bu0uh_wb51w, a82ka7y2g, gf33atgy, ru_wi);
wire [64-1:0] uxphpj98_831n = dn8riluj40uunvq5 ? a82ka7y2g : {a82ka7y2g[64-1:2],2'b0};
assign h_qwsgi7nk2 = uxphpj98_831n; 







wire [64-1:0] kmwz7do01j; 

wire wz0g6uqf = (e1go3iu == 12'h107);
wire u38vpo6j2uw3 = el7_p8jit09 & wz0g6uqf;
wire aeo3kt4q_8k = a94vd35etec4 & wz0g6uqf;
wire yqktpgrj = (aeo3kt4q_8k & izhvh9xxvwe2);
wire [64-1:0] zotth5kymnff =  {vf5xcr67bqhzlo43_[64-1:v_1vibiyou7ysbpkunv],{v_1vibiyou7ysbpkunv{1'b0}}}; 
wire [64-1:0] wbv8vx7udw;
ux607_gnrl_dfflr #(64) eip2ref6zmye (yqktpgrj, zotth5kymnff, wbv8vx7udw, gf33atgy, ru_wi);
wire [64-1 :0] i88tw2wiyz = wbv8vx7udw;
assign kmwz7do01j = wbv8vx7udw; 
assign d3hccrck1fl7jjf6 = {kmwz7do01j[(64-1):(m_rz39tx6bnugdx+3)],b4lwcgm6l21pi[m_rz39tx6bnugdx-1:0],3'b0};



assign ja2k8c_59wnmay5l = (e1go3iu == 12'h140);
assign ng7hgd38lorxo = ja2k8c_59wnmay5l & el7_p8jit09;
assign eo9lmvnadbu765 = ja2k8c_59wnmay5l & a94vd35etec4;
assign tf6c6wjqdv5vvu4 = eo9lmvnadbu765 & izhvh9xxvwe2;
wire hu94wuklp3oosx9df12j75vb0dqh;
wire fxp6atgiv6o9l7nxqxskuxxdkknk;
assign rbz4pv_atxqopdwt = tf6c6wjqdv5vvu4 | hu94wuklp3oosx9df12j75vb0dqh | fxp6atgiv6o9l7nxqxskuxxdkknk;
wire [64-1:0] sscratch_r;
assign qs1xgat7r8xow = vf5xcr67bqhzlo43_;
ux607_gnrl_dfflr #(64) w3anjuevpxzh4v (rbz4pv_atxqopdwt, qs1xgat7r8xow, sscratch_r, gf33atgy, ru_wi);
wire [64-1:0] y2ore77f3hund = sscratch_r;



assign b4etkbmloh = (e1go3iu == 12'h141);
assign ven2nsl = b4etkbmloh & el7_p8jit09;
assign zy44s2bwza9 = b4etkbmloh & a94vd35etec4;
assign m4xr4juqkq = zy44s2bwza9 & izhvh9xxvwe2;
wire xziuk0cj = m4xr4juqkq | z2g63deibg1b1quqr;

wire [64-1:0] x0fgxfber0q;
wire [64-1:0] l8fb_7ff6g;


assign l8fb_7ff6g[64-1:1] = 
        z2g63deibg1b1quqr ? p5jpgn4rvarpo[64-1:1] :
        vf5xcr67bqhzlo43_[64-1:1];
assign l8fb_7ff6g[0] = 1'b0;
ux607_gnrl_dfflr #(64) zss_bvvm_m_b_0 (xziuk0cj, l8fb_7ff6g, x0fgxfber0q, gf33atgy, ru_wi);
wire [64-1:0] csr_sepc;
assign csr_sepc   = x0fgxfber0q;  
assign bde41te346q515l = x0fgxfber0q;  



assign no4tukpi8i35 = (e1go3iu == 12'h142);
assign elq67c0en7exei = no4tukpi8i35 & el7_p8jit09;
assign fzwoxh5vqm8 = no4tukpi8i35 & a94vd35etec4;
assign syf4axzj9zyr = fzwoxh5vqm8 & izhvh9xxvwe2;
wire [64-1:0] qw8gu_4ag_hhlvq;
wire [64-1:0] o9smu2vou412;

wire wzy38v6ckq5dzl2 = syf4axzj9zyr | dhjwho76fa8hqc;   

assign qw8gu_4ag_hhlvq[64-1]  = dhjwho76fa8hqc ? u25pqekq4df[64-1] : vf5xcr67bqhzlo43_[64-1];


assign qw8gu_4ag_hhlvq[64-2:0] = {(64-1){1'b0}};
wire qlvy5r_3uh;
wire xbuq7x2mqt1;
ux607_gnrl_dfflr  #(1) z_6o90lqn6kt_st5uwsm1 (wzy38v6ckq5dzl2, qw8gu_4ag_hhlvq[64-1], o9smu2vou412[64-1], gf33atgy, ru_wi);
wire qpp_vt8_ds5mvm97q = dn8riluj40uunvq5 & (syf4axzj9zyr | xbuq7x2mqt1 | miax48k27o484e8a);

wire r1_9e6hksw6buoti2e1nbxqm_k3;
assign xbuq7x2mqt1 = hze_3v_qjwxi4mrbnkcnic 
               | r1_9e6hksw6buoti2e1nbxqm_k3
              ;

wire ktncdud7tycqpy = xbuq7x2mqt1   ? 1'b1 :
                 miax48k27o484e8a ? 1'b0 :
                 syf4axzj9zyr ? vf5xcr67bqhzlo43_[30]:
                 qlvy5r_3uh;
ux607_gnrl_dfflr  #(1) d7gb5o0uz5oyak2dbyabgw (qpp_vt8_ds5mvm97q, ktncdud7tycqpy, qlvy5r_3uh, gf33atgy, ru_wi);

wire jl2f_lr3ax_x =  dn8riluj40uunvq5 & (ymnk8i8eh3n9_ib7224 | syf4axzj9zyr);   

wire [7:0] efq4x16;
wire [7:0] gy2l1zlyhr =   ymnk8i8eh3n9_ib7224  ?  tcy_87vt9vet39knuw :
                        syf4axzj9zyr   ?  vf5xcr67bqhzlo43_[23:16] :
                        efq4x16;
ux607_gnrl_dfflr  #(8) ri03gy6_ytvbl3754ewyww (jl2f_lr3ax_x, gy2l1zlyhr, efq4x16, gf33atgy, ru_wi);

wire iu3bci_z0jchb0ss9unjyripebx;
wire vsyco_yl80nt2jkmm = wzy38v6ckq5dzl2 | iu3bci_z0jchb0ss9unjyripebx;
wire [ob0j3iecn59nr6s8ur-1:0] jy8ubxm932qii1hd2p; 
wire [ob0j3iecn59nr6s8ur-1:0] nicsojva70v_rf803qb = dhjwho76fa8hqc          ? u25pqekq4df[ob0j3iecn59nr6s8ur-1:0] :
                                               iu3bci_z0jchb0ss9unjyripebx ? {{ob0j3iecn59nr6s8ur-m_rz39tx6bnugdx{1'b0}},b4lwcgm6l21pi[m_rz39tx6bnugdx-1:0]} 
                                             : vf5xcr67bqhzlo43_[ob0j3iecn59nr6s8ur-1:0];

ux607_gnrl_dfflr  #(ob0j3iecn59nr6s8ur) dn0jytq_z7yu0xe1dblot (vsyco_yl80nt2jkmm,nicsojva70v_rf803qb,jy8ubxm932qii1hd2p,gf33atgy,ru_wi);

assign o9smu2vou412[64-2:31] = {(64-32){1'b0}};
assign o9smu2vou412[30] = dn8riluj40uunvq5 ? qlvy5r_3uh : 1'b0;
assign o9smu2vou412[29] =  1'b0;
assign o9smu2vou412[28] =  dn8riluj40uunvq5 ? ogmro605vz43jd_a6 : 1'b0;
assign o9smu2vou412[27] =  dn8riluj40uunvq5 ? ty64g8m1v81v7625 : 1'b0;
assign o9smu2vou412[26:25] =  2'b0;
assign o9smu2vou412[24] = 1'b0;
assign o9smu2vou412[23:16] = dn8riluj40uunvq5 ? efq4x16 : 8'b0;
assign o9smu2vou412[15:ob0j3iecn59nr6s8ur] = {(16-ob0j3iecn59nr6s8ur){1'b0}};
assign o9smu2vou412[ob0j3iecn59nr6s8ur-1:0] = jy8ubxm932qii1hd2p;


assign tvh1llq2i3_y = o9smu2vou412;



assign bh9_1u0btegoxnhc_ = (e1go3iu == 12'h143);
assign rmh20fa2i1zgb = bh9_1u0btegoxnhc_ & el7_p8jit09;
assign wy0jv5w_isf0qmqb = bh9_1u0btegoxnhc_ & a94vd35etec4;
assign pyczk46mr25dxfykg = wy0jv5w_isf0qmqb & izhvh9xxvwe2;  
wire uywyh0w5bkruximyfbbnb8w62 = u_ufp_wg29ieoklxxz1;   
wire nnyi5v6gcq1de = pyczk46mr25dxfykg | uywyh0w5bkruximyfbbnb8w62;
wire [64-1:0] r00ij28c0dqg;
wire [64-1:0] ln9lpk9i_r3jnjtvo;
assign ln9lpk9i_r3jnjtvo = uywyh0w5bkruximyfbbnb8w62 ? tlgcdv86voe9 : vf5xcr67bqhzlo43_;
ux607_gnrl_dfflr #(64) tocvqteqn6pfvxx_ (nnyi5v6gcq1de, ln9lpk9i_r3jnjtvo, r00ij28c0dqg, gf33atgy, ru_wi);
wire [64-1:0] d9jmhohu_gk6;
assign d9jmhohu_gk6 = r00ij28c0dqg;



assign ha7fcf0ap = (e1go3iu == 12'h144);
assign uz6ke_lem = ha7fcf0ap & el7_p8jit09;
assign ano1d1_31 = (~dn8riluj40uunvq5) & ha7fcf0ap & a94vd35etec4;
assign kkco_owc1 = ano1d1_31 & izhvh9xxvwe2;

assign i9xvsmm45fp0f58 = pvfk1_6o89lmby & xc_4r6ncv72;
assign w529wbj853 = xx87vzbpchg & m00o8sz4cyd_a9;



assign ezl3jzeqhltgj7h = fgr486jx5kevbua;

wire [64-1:0] xzml2u6ee;
assign xzml2u6ee[64-1:22] = 10'b0;
assign xzml2u6ee[21] = 1'b0;
assign xzml2u6ee[20] = 1'b0;
assign xzml2u6ee[19] = 1'b0;
assign xzml2u6ee[18] = 1'b0;
assign xzml2u6ee[17] = 1'b0;
assign xzml2u6ee[16] = 1'b0;
assign xzml2u6ee[15:12] = 4'b0;
assign xzml2u6ee[11:10] = 2'b0;
assign xzml2u6ee[9]     = ezl3jzeqhltgj7h;
assign xzml2u6ee[8:6]   = 3'b0;
assign xzml2u6ee[ 5]    = w529wbj853;
assign xzml2u6ee[4:2]   = 3'b0;
assign xzml2u6ee[ 1]    = i9xvsmm45fp0f58;
assign xzml2u6ee[ 0]    = 1'b0;

assign csr_sip = dn8riluj40uunvq5 ? 64'b0 : xzml2u6ee;


assign ddx7351w3ukkafuh3 = o9smu2vou412[64-1];

assign rjju_oexoi2ozf1eo = ddx7351w3ukkafuh3 & s_m3pbf5m2tr6v;  
assign ymnk8i8eh3n9_ib7224 = hvy2cpsp75f3 & z2g63deibg1b1quqr;        
assign hze_3v_qjwxi4mrbnkcnic  = ymnk8i8eh3n9_ib7224 & k3z202os;







assign vqvbmvk4f_b_c = (e1go3iu == 12'h180);
assign dk878usgx2r = vqvbmvk4f_b_c & el7_p8jit09;
assign vcsyiox9w = vqvbmvk4f_b_c & a94vd35etec4;
assign lqzw29rbc73ulx = vcsyiox9w & izhvh9xxvwe2;
wire am4nk9up = lqzw29rbc73ulx;

wire [64-1:0]    eclvpk;
wire [64-1:0]    ivwaytj4;
wire [64-1:0]    hs867vkzot86;


assign hs867vkzot86[64-1] = vf5xcr67bqhzlo43_[64-1]; 
assign hs867vkzot86[64-2:64-4] = 3'b0;
assign hs867vkzot86[64-5:0] = vf5xcr67bqhzlo43_[64-5:0];

ux607_gnrl_dfflr #(64) gt4eho16x8 (am4nk9up, hs867vkzot86, eclvpk, gf33atgy, ru_wi);


assign ivwaytj4 = eclvpk;  



wire v4u8py6g9qm7nxnzm93vex;
wire xmlgz6ri7nmdy67 = (e1go3iu == 12'h146);  
wire yry8e0jbvce3okne = el7_p8jit09 & xmlgz6ri7nmdy67;
wire x9uju93rexa6wv =dn8riluj40uunvq5 & ( v4u8py6g9qm7nxnzm93vex
                                     | ymnk8i8eh3n9_ib7224
                                     | rjju_oexoi2ozf1eo); 

wire [64-1:0] p_rxkqn5_ysam3gaisn = (v4u8py6g9qm7nxnzm93vex | ymnk8i8eh3n9_ib7224) ? {{(64-16){1'b0}}, hjrk_rwjkqj3zk_b,8'h0} :
                                                                 rjju_oexoi2ozf1eo ? {{(64-16){1'b0}}, efq4x16,8'h0}       :
                                                                                    sintstatus_r;
ux607_gnrl_dfflr #(64) jjduwuoiy7w3s3dm5s2i (x9uju93rexa6wv, p_rxkqn5_ysam3gaisn, sintstatus_r, gf33atgy, ru_wi);
wire [64-1:0] b4f0p1edkro3ny90i8 = sintstatus_r;
assign tcy_87vt9vet39knuw = sintstatus_r[15:8];




assign xrbzeq_xg1z9 = (e1go3iu == 12'h9c0);
assign e364tfszybtw35 = xrbzeq_xg1z9 & el7_p8jit09;
assign h9bg0vmhmf = xrbzeq_xg1z9 & a94vd35etec4;

wire u74l6ss7cdyx = (h9bg0vmhmf & izhvh9xxvwe2) | icauf4l_12_c2xkj53lf;
wire [64-1:0] l15mfr53w;
wire [64-1:0] m8efbb1yrkp5o;
assign m8efbb1yrkp5o[64-1:3] = {64-3{1'b0}};
assign m8efbb1yrkp5o[3-1:0] = 
                   icauf4l_12_c2xkj53lf ? xel6gw173w5x0[3-1:0] 
                                   : vf5xcr67bqhzlo43_[3-1:0];

ux607_gnrl_dfflr  #(64) k3h4m6coan_zzdb0 (u74l6ss7cdyx, m8efbb1yrkp5o, l15mfr53w, gf33atgy, ru_wi);
wire [64-1:0] znodfv_85_bqx9 = l15mfr53w;




assign ls416x5_x21tvc = 1'b0;
assign d1bjdianldviz8 = ls416x5_x21tvc & el7_p8jit09;
assign e3t8l4w0xlvk50p = ls416x5_x21tvc & a94vd35etec4;

wire uhubewjnc1uej = (e3t8l4w0xlvk50p & izhvh9xxvwe2) | e_z6d7r9kxqg32te;
wire [64-1:0] qr88cvk3fc4h;
wire [64-1:0] g94vtj5nko43557;
assign g94vtj5nko43557[64-1:5] = {64-5{1'b0}};
assign g94vtj5nko43557[5-1:0] = 
                   e_z6d7r9kxqg32te ? v8ydjtlz16x9tx[5-1:0] 
                                   
                                   : 5'b0;

ux607_gnrl_dfflr  #(64) nb8yg09y2jqwr8 (uhubewjnc1uej, g94vtj5nko43557, qr88cvk3fc4h, gf33atgy, ru_wi);
wire [64-1:0] fk85rb7md5gw3sw = qr88cvk3fc4h;




wire j1ylmn_bzfrz_ = (e1go3iu == 12'h145); 
wire j5kvlkrjxy = el7_p8jit09 & j1ylmn_bzfrz_;











wire dgadiuf5wx3oc3q6fi = (e1go3iu == 12'h148);
wire jsnbl6829nsp81ae = el7_p8jit09 & dgadiuf5wx3oc3q6fi;
wire k5jua7kub3him5uq5tsz9 = dgadiuf5wx3oc3q6fi & (ogmro605vz43jd_a6 != 1'b1);  
assign hu94wuklp3oosx9df12j75vb0dqh = izhvh9xxvwe2 & k5jua7kub3him5uq5tsz9; 
wire [64-1:0] ui1hd0tbisqqo5glc4kc = k5jua7kub3him5uq5tsz9 ? y2ore77f3hund : vmx1fh4kmh4c;











wire a7xf2tgo_tq3co7fsn5l9 = (e1go3iu == 12'h149);
wire tgxhzbu4fzxohws9_0 = el7_p8jit09 & a7xf2tgo_tq3co7fsn5l9;
wire xru5c6rzjn = (efq4x16 == 8'b0);
wire sgf5ditx2uzyicptvtom = (tcy_87vt9vet39knuw[7:0] == 8'b0);
wire i1ubl3bjccmw7ajzl6n = (xru5c6rzjn != sgf5ditx2uzyicptvtom) & a7xf2tgo_tq3co7fsn5l9 & dn8riluj40uunvq5;
assign fxp6atgiv6o9l7nxqxskuxxdkknk = izhvh9xxvwe2 & i1ubl3bjccmw7ajzl6n; 
wire [64-1:0] wmaji4s5cfj1 = i1ubl3bjccmw7ajzl6n ? y2ore77f3hund : vmx1fh4kmh4c;
wire [64-1:0] fp2zbc8_89qlmg_v9 = dn8riluj40uunvq5 ? wmaji4s5cfj1 : 64'b0; 




assign uy_j_dcfffe0 = (e1go3iu == 12'h947);
wire bdhgj6khs_7ga3 = el7_p8jit09 & uy_j_dcfffe0;


wire f22sj2magiajlxzz1 = j1ylmn_bzfrz_ 
                       | uy_j_dcfffe0 
                       ;

wire rnt3vdbdjmztyc4 = f22sj2magiajlxzz1  
                        & y8_gkxsfle                   
                        & fc_4ns_w1nh4h02z_dgg       
                        & gfy3zost37aq8qmr
                        & (hjrk_rwjkqj3zk_b > efq4x16)  
                        & (~zwcbp7zqfei5xz) 
                        & dn8riluj40uunvq5;

assign v4u8py6g9qm7nxnzm93vex = rnt3vdbdjmztyc4 & izhvh9xxvwe2;
assign iu3bci_z0jchb0ss9unjyripebx = v4u8py6g9qm7nxnzm93vex;

wire [64-1:0] dogg7s_r84uw;
assign dogg7s_r84uw = {i88tw2wiyz[(64-1):(m_rz39tx6bnugdx+3)],b4lwcgm6l21pi[m_rz39tx6bnugdx-1:0],3'b0};

wire [64-1:0] yjhxn3cnn387p4 = rnt3vdbdjmztyc4 ? 
                                          dogg7s_r84uw 
                                          : 64'b0;


assign fzdb65fcrotwcaccus_cwo = v4u8py6g9qm7nxnzm93vex;
assign f4_gpy7hep0c0klauu = f22sj2magiajlxzz1 & izhvh9xxvwe2;

wire [64-1:0] zyi73htc0wk = rnt3vdbdjmztyc4 ?         
                                   nchi0_6mu
                                   : vmx1fh4kmh4c;

wire [64-1:0] m3d19g2wsmf9x2em = dn8riluj40uunvq5 ?  zyi73htc0wk : 64'b0;
assign psx330qmvh5so1to4iq = fzdb65fcrotwcaccus_cwo & uy_j_dcfffe0;  
assign hzsp_nydab9ghw59v  = dogg7s_r84uw[64-1:0]; 
assign rl9a96pgy3troiao05jel  = 1'b1;
assign bzz8x0np0dpmdjt1d0w7uf  = pydatzxqqi;
assign sefocn4wjn2k2f_zvlvnz  = aw82i964do;
assign qknomh2kbth19r1osddvzly  = y8_gkxsfle;
assign r1_9e6hksw6buoti2e1nbxqm_k3  = psx330qmvh5so1to4iq & rl9a96pgy3troiao05jel;



wire [64-1:0] shs9_ifu4; 

wire mb9dfbm5rqlncg = (e1go3iu == 12'h948);
wire d9i_mw1cltd = el7_p8jit09 & mb9dfbm5rqlncg;
wire i97eur_3x = a94vd35etec4 & mb9dfbm5rqlncg;
wire w8rx22hkc = (i97eur_3x & izhvh9xxvwe2);
  
wire [64-1:0] b2v38pbv2n =  {vf5xcr67bqhzlo43_[64-1:2],1'b0,vf5xcr67bqhzlo43_[0]}; 
wire [64-1:0] gb7osa4w9;
ux607_gnrl_dfflr #(64) bw73sxcx7l0 (w8rx22hkc, b2v38pbv2n, gb7osa4w9, gf33atgy, ru_wi);
assign shs9_ifu4 = gb7osa4w9; 
assign vkyge0q4mfc5 = shs9_ifu4[0];  

assign cppkd01vpwwnlfy = shs9_ifu4;  














assign zmfo8cca_77pc = csr_sstatus;    
assign hig2gwwbeuhnt65xrp = csr_mstatus;
assign {u2dvoyt5e7o_03z9z5, l9erxxpnphqd26vg9} = {1'b0,64'b0} 
               | {vybduk_04wdx6z05      , ({64{x4_1imazttasol8      }} & uwpy_1502jyu8_t80s)}
               | {z49s15yop6m7rk           , ({64{hyvne9dzw           }} & luex1cs6x7sa)}
               | {k9p_ach              , ({64{wuiysx              }} & inyyxdi9)}

               | {fb_inlkctcnic    , ({64{m_l49l2tvr3sko    }} & csr_mstatus  )     }
               | {gfy9n09ir7q8zrpld19  , ({64{fw0ba932spu6w15bn  }} & v0k9xrr0s5wwex3)     }
               | {b2uwf6iur0a5ek5x9    , ({64{b8ao64rq4cnci    }} & wsr5asmu2rsl6a076  )     }
               | {x06wm7qebv8ymb    , ({64{pssagx292xg6    }} & pealk1ny1w3zypaet  )     }
               | {y_nu4e3x8595566bl  , ({64{pa1_agmr_3hhej4  }} & oxqig8tg9r_4az4sf)     }
               | {od1i6efig3fvtth  , ({64{djtm53o1_m_3x_4o  }} & clr_f9f2zh_fkkespze)     }
               | {zo5qd8wbwszeiqaye  , ({64{kxurpsnfj171m_n2_3aq  }} & t_7nv9a3lsvuzxmcw)     }
               | {rmx1zc2nonjyho98zpr_  , ({64{pu3hs090altkbczlh  }} & bqp1xynoo31eoavfit1)     }
               | {tc3f_x03mu_vagb8bx2 , ({64{b0g_t6oj33jh4lf_l55 }} & rziri8ijn84w3o8cp)    }
               | {ye2xj3py3c5f_h_b8f , ({64{hvopxeap8rqft0nnorg }} & f36cakmqdwzxjjajghlg)    }

               | {wft1k16f78xw2   , ({64{aaa3cgvzwhecdc46s   }} & epnwm13_bdyvjd )     }
               | {jan2q6micau0n4    , ({64{xd1ve1tqh9v    }} & csr_medeleg  )     }
               | {ls8dsrnc8qwzmpg    , ({64{ekglglw24_squr    }} & csr_mideleg  )     }
               | {ps869z4s        , ({64{wwc6g7        }} & csr_mie      )     }
               | {etyac0jmfrzxm      , ({64{t4fpmjlqyt      }} & p41zr5gkln    )     }
               | {b9p2i13nz      , ({64{ycvvi2q5      }} & glwac019m8pq    )     }
               | {b8m44m4dqrd       , ({64{bk92fvsycux       }} & csr_mepc     )     }
               | {l52o_50oot2j6   , ({64{rud1hmcy9tubf9k   }} & klnr5w9m7dv5ejwl )     }
               | {di2d3ktm1fz_8we     , ({64{k2zpid7lzqutl     }} & p6rw9no76a3m   )     }
               | {fgc4ur8_m02    , ({64{t3h801u9ezg0    }} & it8le0crf9kmfqe  )     }
               | {d521va8_2d6_c7j   , ({64{gbj6z3zlspk3_b9   }} & viqilm0l71xjf5c )     }
               | {zavn9glbl0j62qi   , ({64{jbbx5w95zgs1   }} & ga1zsr158e3cs9vru )     }
               | {yoegchl8        , ({64{oekhv_        }} & csr_mip      )     }
               | {o9ci7gemz       , ({64{tqmr31e       }} & a1sjkc9c8      )    }
               | {m8rmfuha0pch8g  , ({64{swp0cfl7pff8oo4  }} & hkvtut3x96fj_tl)     }
               | {pjwkxwhqy7i     , ({64{ofj_z8n6541s     }} & qyirue3_ioqbr   )     }
               | {os_f3xrbfr2or    , ({64{e1j7flhjhq    }} & hnd2jesdfkehin  )     }
               | {kp2w957z1v     , ({64{tcpea5afm7of     }} & uonsn384se50   )     }
               | {b18orstady8x36yc    , ({64{owcdacpz2mm    }} & mvsg2qxdmt29ncr9  )     }
               | {bun2s3y6z8vtjyxjzr9, o02hm9vkepj5rucwrif                            }
               | {wew7vt2_2h6k      , ({64{hcqw9t9s      }} & cyxvmxf7k3h7   )     }
               | {i7e201yj       , ({64{kp2q6bh2       }} & tuh58_qx     )     }
               | {xcfnsabp39vvwn    , ({64{gkxo6i5s875r    }} & pltp40lm289gs )     }
               | {wsps0651m      , ({64{crgfb_c8n      }} & yrf31busye76   )     }
               | {mx6n8ae8twuk2mfjz_1 , ({64{xlchao2g44p1tat_  }} & t7gzjhdzm9ftqnv7)   }
               | {cgnhh8s1vo2cuntv, ({64{zcege9lvdnn7d5f}} & ixkez_bglcky89d58tfw3)}


               | {p7zidsgtr9q7bf81 , ({64{ka2utev6jddufp7b9}} & hxxl4aq4sjdycyml2)  }
               | {mwegg_7inaca6povsw, bsjo0v5e0t556pph                            }

               | {zj201cydmy_kb    , ({64{l0o8bky903    }} & vbw35s4mu01jg4  )     }

               | {vadpkdaztv820a8kvwp0, mj56s1rlw1lf7pkf2icn8d                            }
               | {iiq92rsh_v1ylb    , ({64{il_e54l8ycmz2u    }} & csr_sstatus  )     }
               | {qb5qu1p3        , ({64{myuno7j        }} & csr_sie      )     }
               | {qtf8of_u5z5iai      , ({64{ed9vgeh97yj      }} & uxphpj98_831n    )     }
               | {ja2k8c_59wnmay5l   , ({64{ng7hgd38lorxo   }} & y2ore77f3hund )     }
               | {b4etkbmloh       , ({64{ven2nsl       }} & csr_sepc     )     }
               | {no4tukpi8i35     , ({64{elq67c0en7exei     }} & tvh1llq2i3_y   )     }
               | {xrbzeq_xg1z9    , ({64{e364tfszybtw35    }} & znodfv_85_bqx9  )     }
               | {ls416x5_x21tvc   , ({64{d1bjdianldviz8   }} & fk85rb7md5gw3sw )     }
               | {bh9_1u0btegoxnhc_   , ({64{rmh20fa2i1zgb   }} & d9jmhohu_gk6 )     }
               | {ha7fcf0ap        , ({64{uz6ke_lem        }} & csr_sip      )     }
               | {vqvbmvk4f_b_c       , ({64{dk878usgx2r       }} & ivwaytj4     )     }
               | {xmlgz6ri7nmdy67 , ({64{yry8e0jbvce3okne }} & b4f0p1edkro3ny90i8)    }
               | {j1ylmn_bzfrz_      , ({64{j5kvlkrjxy      }} & yjhxn3cnn387p4    )     }
               | {wz0g6uqf       , ({64{u38vpo6j2uw3       }} & kmwz7do01j     )     }
               | {dgadiuf5wx3oc3q6fi,({64{jsnbl6829nsp81ae }} & ui1hd0tbisqqo5glc4kc)   }
               | {a7xf2tgo_tq3co7fsn5l9,({64{tgxhzbu4fzxohws9_0}}& fp2zbc8_89qlmg_v9)  }
               | {uy_j_dcfffe0    , ({64{bdhgj6khs_7ga3    }} & m3d19g2wsmf9x2em  )     }
               | {mb9dfbm5rqlncg      , ({64{d9i_mw1cltd      }} & shs9_ifu4    )     }
               | {vu_8rttl4p4     , ({64{mxqvlgcks     }} & cdiut_mads8ok7   )     }
               | {doorarnn829tt     ,  ({64{vzxftoy0      }} & vgcvjr8adr    )     }
               | {f8nehtdp4c9jo5           , ({64{lsbmvjc19i           }} & ywq7zmowlccfib)}
               | {jjvcrtzj366t  , ({64{zmgxfaohma89cv5  }} & aur5f30tjm74ynd)     }
               | {a06ag5mfqc7b  , ({64{l7r01a30uiu  }} & vxt5pb8sxldtxqw)     }
               | {skog6xw8aj1km8ost  , ({64{noizhmz52v5iwfm  }} & p3kutuvsyvsd)     }




               | {ad2bzpfqdx       , ({64{k1j9zf14hj       }} & ove0jfc9_     )     }
               | {veysvh0g_5rkx       , ({64{n4vaq5qq96wr       }} & ae1hd9imgwd     )     }
               | {andomkgjr       , ({64{rvkrf8rv4n       }} & b0en4jlm5ni5     )     }
               | {dfkhf0zzmeauwtqm3som, (p744ug1jil846r8g6p)                                 }
               | {by_qc3yb1cyytd, ({64{xdxa3krj224xup     }} & k427ik6bety0vdf)        }
               | {fk5t4onucgv   , ({64{hx6va8sy        }} & bw8e1bo__j   )        }
               | {lc6w646en  , ({64{t1muoi2gjx2o       }} & g8cty956i  )        }
               | {sim0gblc86voze3mam, ({64{n1zvf0y1dwpep }} & htdx5bpibi4z9nvhfcy  ) }
               | {dxb0y6x6tzh8_cwt2    , ({64{1'b0 }} ) } 
               ;



  assign l_jd4i6dsmcejyydh =  a94vd35etec4 & ( 







                 m8rmfuha0pch8g
               | os_f3xrbfr2or  
               | kp2w957z1v   
               | b18orstady8x36yc   
               | jjvcrtzj366t 
               | a06ag5mfqc7b 
               | skog6xw8aj1km8ost 
               | pjwkxwhqy7i 
               ) ;



  assign s36z1abpqp = (~aw82i964do) & (~y8_gkxsfle) & (~pydatzxqqi);

  wire al4ew6cc9jzsnvt2piq6 = ( 1'b0 
                  | by_qc3yb1cyytd    
                  | fk5t4onucgv       
                  | lc6w646en      
                  | k9p_ach
                  | z49s15yop6m7rk
                  | vybduk_04wdx6z05
                  | f8nehtdp4c9jo5
                  | vu_8rttl4p4
                  | doorarnn829tt
                  | ikq8fffiwai0wlaxzs4xfv08i
                  | dxb0y6x6tzh8_cwt2
                 );

  wire o1ofai8pfroxnslalvk3 = s36z1abpqp &
                   
                   
               (~( 1'b0
                  | maynsergszxlh4jomqhce5ahk     
                  | al4ew6cc9jzsnvt2piq6     
                  ))
               ;


  assign f982i0gj5cmkoid = o1ofai8pfroxnslalvk3 | wfndbkyoc1wc094vwehhutg5krtg
                         | wjtx1c23l6psom27nm_gsj1ljb2
                         ;
  assign iu2o274ax6rzokmi0 = ad6d6ex80to7t3vvnc69u3pmz;



  wire ub1xslm06r09rvx11 = ( 1'b0 
                  | iiq92rsh_v1ylb
                  | qb5qu1p3 
                  | qtf8of_u5z5iai
                  | ja2k8c_59wnmay5l
                  | b4etkbmloh
                  | no4tukpi8i35
                  | xrbzeq_xg1z9
                  | ls416x5_x21tvc
                  | bh9_1u0btegoxnhc_ 
                  | ha7fcf0ap
                  | vqvbmvk4f_b_c
                  | xmlgz6ri7nmdy67
                  | j1ylmn_bzfrz_
                  | wz0g6uqf
                  | dgadiuf5wx3oc3q6fi
                  | a7xf2tgo_tq3co7fsn5l9
                  | mb9dfbm5rqlncg
                  | uy_j_dcfffe0
                  | al4ew6cc9jzsnvt2piq6     
                  | eu5gus8kcfxe2bn_5jpy90jbl
                 );

  wire ub8hotlnbvgn8ttgzq = y8_gkxsfle & (~pydatzxqqi) &
                   
                   
               (~( 1'b0
                  | oi73ilapk89bv0c9d4nvacia05brp     
                  | ub1xslm06r09rvx11     
                  ))
               ;


  assign brfqcqo_b08lybzgt = ub8hotlnbvgn8ttgzq | cry3qyaqkl89ztcpeizdmn2fj
                         | nug315vy7hnf899pgdpd2t7oh8
                         ;
  assign ve7t8hdsd1_tnt9v = eil4t6r56iactzfh4_drmg7xv;
















  assign j0qaxhuqtdi      = rb050tnl     ;
  assign pbzpk52jinfscit4mm    = a94vd35etec4   ;
  assign gwj6ow6qvbhs0tc31    = el7_p8jit09   ;
  assign mm0ssgy582fv_j      = e1go3iu     ;
  assign iwdkm52x_w4hpak_a2_w = izhvh9xxvwe2;
  assign ir2913p9xpmq_1bvfd1 = vf5xcr67bqhzlo43_;


  assign st2zalpx0uf = dttzf_6vv87y;
  assign ni01kj42oob2x = csr_mstatus[19];
  assign ah8kjlmvnaxzbi = csr_mstatus[18];
  assign fkuqlh34r   = ivwaytj4[64-1]; 
  assign hnc10arn_rd   = ivwaytj4[20 + 16 -1 : 20];
  assign b2ulqcjb    = ivwaytj4[20 -1 : 0];
  assign w30ye15yns15    = status_priv_r;

endmodule




















module jgz9v2pi3n5adi7j41(



  input  [32-1:0] k0xug5g,
  input  qhyq467foflgyn5y, 
  input  sa2f4h4xeakpfnunl,           
  input  u2k4dyp52s_m,
  input  djvj1e_,
  input  bktu0z1mk56,
  input  qbsr1jytrqtsbk4ttb8nz,
  input  b0ry73kp6sc2,
  input  hr64e6c3gy ,
  input  cz1hh6af7xp2,

  input  s1woka0byzgo,
  input  al4xeg8mukgfg,
  input  piwiqvrjoq,
  input  wi_dfzp70x09hm1m,
  input  jdyqycv3wdp2sgy,


  input  rnx27onf2lbe, 


  output g_o2wra9n9s,
  output nykwng_3anppxi,
  output shpynlimbt55rj4,
  output jycwup76klyed6d2,
  output i7pubsxfsb4uys,
  output [5-1:0] jc4yg1pkylr2gonwcd,
  output [5-1:0] nd3cgvec1pogf2,
  output [5-1:0] f7crsrzernrwgmepy,
  output [5-1:0] pw085ct76po3c,
  output [48-1:0] g5usf8ixwjaxjs1m,
  output [64-1:0] pxhhgm9746n,
  output fgm5kq4y725x6yylw,
  output awld9ngcypgfxa,
  output v5m66onlnmxeejfhn,
  output kfz3mojvfh2fsfd,

  output                           d40y0va2l7xzj,
  output [48-1:0] hhj5975j18r0n,

  output m05tjqf24b1fabuu0e, 


  output mg0onistbzu9ys,
  output g3btysb7vvv,
  output yjgkn7vcv,
  output sb8ax73d3ud,
  output f9_w27gbcq__,
  output iq9sj_i8z1k712,
  output b6cv9yeaga7hf,
  output [5-1:0] rig48lgqgq8oxt,    
  output [5-1:0] zaub9z0lm4s93y,    
  output [5-1:0] kd6v2vk601xpnm,     
  output [5-1:0] j_69hsshtbv,    


  output [64-1:0] t05leas4w4r,
  output fpwql5ik7_sp0,
  output dwci8hbxok739,
  output fqizcmmfg,
  output tbuacpjktio,
  output ciftsjs2bvaxns,
  output k_y4yq3crp_zqtg,
  output [31:0] zk9uk90j08ogqpn,

  output [19-1:0] eaxqugrf_ryu5rxxw41,
  output tkm5u9dl8zav4,

  output [105-1:0] z8t7w6zr5woh649,
  output [50-1:0] mg4yq4mui7ruja,
  output sibtd2rf5j,
  output hgvdw0qnels8,

  output qzdlalytscynhz1,

  output vfye1vj155_k,
  output vujduks2o30,
  output y4zqru1tedm,
  output q1coyps2cz7xe,
  output oli3_udj80h6urj,
  output rphjsg75001l2,
  output ch8qv98q9xu469etyz8oj,
  output [48-1:0]  zj0wqwminaxn,

  output t9xs6bqphiru,
  output ls1dudpc   ,
  output tzjssx03b   ,
  output cni2453cuofb   ,
  output kt04okvuth  ,
  output kq9gup8pu2  ,

  output nnng_p6632p,
  output ld01d40_n3,
  output o8rwk067,
  output r1on2k03r,
  output gw7452ctd577,
  output b1roq8tr9r,
  output j_ku88w81rg,
  output jw1vgacy_r0vr,

  output [5-1:0] ng_pudjzgnamv0es,
  output [64-1:0] bdhv0j4zhtx9nxmz 
  );



  wire [32-1:0] pq5pe3yehrqxr = k0xug5g;
  wire [16-1:0] tm0dvbtguid67 = k0xug5g[15:0];

  wire [6:0]  dlmxb1 = pq5pe3yehrqxr[6:0];

  wire wgqy37zae8oexwv  = (dlmxb1[1:0] == 2'b00);
  wire f9k8e7skb6cw2pkw3w  = (dlmxb1[1:0] == 2'b01);
  wire mqwi5z31tkb1fz81y  = (dlmxb1[1:0] == 2'b10);
  wire bfp4chz8bvbs7e8m  = (dlmxb1[1:0] == 2'b11);

  wire vlfahv69 = bfp4chz8bvbs7e8m;

  wire [4:0]  adjmfzwj55ej     = pq5pe3yehrqxr[11:7];
  wire [2:0]  p2f86tlrac56  = pq5pe3yehrqxr[14:12];
  wire [4:0]  ga71__f5g1    = pq5pe3yehrqxr[19:15];
  wire [4:0]  aihiftly    = pq5pe3yehrqxr[24:20];
  wire [6:0]  uk0ahn6nnbba7  = pq5pe3yehrqxr[31:25];

  wire [4:0]  z7cl6tvk     = adjmfzwj55ej;
  wire [4:0]  ag9ylluguwcr    = z7cl6tvk; 
  wire [4:0]  tbilhd3n1v    = pq5pe3yehrqxr[6:2];

  wire [4:0]  oduuhk6i    = {2'b01,pq5pe3yehrqxr[4:2]};
  wire [4:0]  yq79t1_13   = {2'b01,pq5pe3yehrqxr[9:7]};
  wire [4:0]  cjywp5cfm   = oduuhk6i;

  wire [2:0]  xm60rmyor_3v  = pq5pe3yehrqxr[15:13];


  wire d6r44hi25ixatafeu1 = (dlmxb1[4:2] == 3'b000);
  wire cizl6_7mbo_awon = (dlmxb1[4:2] == 3'b001);
  wire vw5it7jugq0nfvd04v = (dlmxb1[4:2] == 3'b010);
  wire bpk53yitybm32g = (dlmxb1[4:2] == 3'b011);
  wire asuyn96in9e48ikear_ = (dlmxb1[4:2] == 3'b100);
  wire kn3z45bkwagekkw = (dlmxb1[4:2] == 3'b101);
  wire cdwv54beu2vbzvh = (dlmxb1[4:2] == 3'b110);
  wire w3imaozzd_v_wb6wo = (dlmxb1[4:2] == 3'b111);
  wire w0s41titqc28jdt  = (dlmxb1[6:5] == 2'b00);
  wire wx_8fko7wy_rmnew7l  = (dlmxb1[6:5] == 2'b01);
  wire sfpsjr_3ucgrnnl4f  = (dlmxb1[6:5] == 2'b10);
  wire f_575odq4qxl04  = (dlmxb1[6:5] == 2'b11);

  wire ezupw6o2yfm5ojugrc3 = (p2f86tlrac56 == 3'b000);
  wire d24iqtxvb2trplxk2m = (p2f86tlrac56 == 3'b001);
  wire t8jc64yc1l6q8eclq_c = (p2f86tlrac56 == 3'b010);
  wire w__ro7gwx6w331 = (p2f86tlrac56 == 3'b011);
  wire d0jauc9xnvhr53rq3 = (p2f86tlrac56 == 3'b100);
  wire tcks0htkit9weu = (p2f86tlrac56 == 3'b101);
  wire o6hnybbrbqkztojg = (p2f86tlrac56 == 3'b110);
  wire dwe8qnpoudm94xa = (p2f86tlrac56 == 3'b111);

  wire mg22fa39qkmi1381_ = (xm60rmyor_3v == 3'b000);
  wire swilkhsvy0ciqh = (xm60rmyor_3v == 3'b001);
  wire ft758uk96h0lere58vu = (xm60rmyor_3v == 3'b010);
  wire t3skb9q5zbu_q_fb = (xm60rmyor_3v == 3'b011);
  wire lkhy22ju1fth_z = (xm60rmyor_3v == 3'b100);
  wire atw4jjamnfmexzna29 = (xm60rmyor_3v == 3'b101);
  wire pw945i12_3q9tpbldo = (xm60rmyor_3v == 3'b110);
  wire f9zuwwm5sc91jd4 = (xm60rmyor_3v == 3'b111);

  wire lrptc0hyjyd7hdoypa0_g = (uk0ahn6nnbba7 == 7'b0000000);
  wire bepkj4gbb77isq3_v9 = (uk0ahn6nnbba7 == 7'b0100000);
  wire t6_6ypj94nny67ise0x9 = (uk0ahn6nnbba7 == 7'b0000001);
  wire xfrai8f3331hb4z5ww5_ = (uk0ahn6nnbba7 == 7'b0000101);
  wire fcpfa9hp28k7bapl82 = (uk0ahn6nnbba7 == 7'b0000110);
  wire hx3wrp4j8s1ov27syy = (uk0ahn6nnbba7 == 7'b0001110);
  wire naged_b50dbpmu745zp = (uk0ahn6nnbba7 == 7'b0010110);
  wire jhbiy5xf0ygws7apfg03 = (uk0ahn6nnbba7 == 7'b0000111);
  wire pvy429fepo5d_7j0eq5ky = (uk0ahn6nnbba7 == 7'b0001001);
  wire cvhx1ne2we07dkbzbpwakl = (uk0ahn6nnbba7 == 7'b0001101);
  wire toaowsb_5w3arwmyl2 = (uk0ahn6nnbba7 == 7'b0010101);
  wire uncepq376ovruspfffvl5 = (uk0ahn6nnbba7 == 7'b0100001);
  wire i0ahgxc7hvmvc1hsbq8 = (uk0ahn6nnbba7 == 7'b0010001);
  wire lipdgvrqr439y_cnsv = (uk0ahn6nnbba7 == 7'b0010010);
  wire veb9c0lxewgh_4qiy5 = (uk0ahn6nnbba7 == 7'b0010011);
  wire k3sfqtpqynzqda4xtugl4 = (uk0ahn6nnbba7 == 7'b0101101);
  wire o5frxem9qrhhps9sw7n = (uk0ahn6nnbba7 == 7'b1111110);
  wire yf083xcjpnohrzqky4 = (uk0ahn6nnbba7 == 7'b1111111);
  wire mso_1l7nnv4ac14pv6qh = (uk0ahn6nnbba7 == 7'b0000100); 
  wire e9hn3j9k88f8miq238hz1 = (uk0ahn6nnbba7 == 7'b0001000); 
  wire duf6qt_vm6jkmkv9xu9 = (uk0ahn6nnbba7 == 7'b0001100); 
  wire gu_2fhfulrttqq4e_fiax = (uk0ahn6nnbba7 == 7'b0101100); 
  wire i6fh1oflvwwzfgicny1c = (uk0ahn6nnbba7 == 7'b0010000); 
  wire f6kcevztmpqpnc8xp3_r4 = (uk0ahn6nnbba7 == 7'b0010100); 
  wire m33lelq8_5u26vfl7hl6z = (uk0ahn6nnbba7 == 7'b0011100);
  wire amf97jdmi0f4r4z2kmw = (uk0ahn6nnbba7 == 7'b0011101);
  wire l6zyb5b3_f8uuon8o3p = (uk0ahn6nnbba7 == 7'b1100000); 
  wire k_h8qestuhin60n5ckxmkfx = (uk0ahn6nnbba7 == 7'b1110000); 
  wire ei5le5r3u2ub_qlszr3u6lq = (uk0ahn6nnbba7 == 7'b1111100);
  wire c7npl5770szduubj6_grim = (uk0ahn6nnbba7 == 7'b1010000); 
  wire tx0e46vrruq3cgq9ghul4 = (uk0ahn6nnbba7 == 7'b1101000); 
  wire v3hylq_n52mziras6qen = (uk0ahn6nnbba7 == 7'b1111000); 
  wire qcpti7i25_4w_aexyk1 = (uk0ahn6nnbba7 == 7'b1100011);
  wire whvtopzve8q_t001lyx = (uk0ahn6nnbba7 == 7'b1010001);  
  wire d9gmx9ccvp0rgcy7n_ii = (uk0ahn6nnbba7 == 7'b1011000);
  wire vrn4ssw1i97fztoyaq5kq = (uk0ahn6nnbba7 == 7'b1011001);
  wire eu9j7rkhrocfjsewdf6mfvu = (uk0ahn6nnbba7 == 7'b1110001);  
  wire rf284mrjg_bqa1hj60swyf = (uk0ahn6nnbba7 == 7'b1111001);
  wire rgjf1vrs4iai2hif_09x = (uk0ahn6nnbba7 == 7'b1100010);
  wire ng7__qxmefe1xunqibay7zg = (uk0ahn6nnbba7 == 7'b1111101);
  wire c9xaw73uh3hmihrn801brf = (uk0ahn6nnbba7 == 7'b1100001);  
  wire mnd8c7lvcdtsypyiygspg = (uk0ahn6nnbba7 == 7'b1101001);  
  wire q8xucja6w9gzw4ujn6f7 = (uk0ahn6nnbba7 == 7'b1000011);
  wire zpue29q3_sghsyln86mp = (uk0ahn6nnbba7 == 7'b1011011);
  wire ef0qt3ctq84209xo8ti63mv = (uk0ahn6nnbba7 == 7'b1011010);
  wire bju5h0qfjwac44bgx65qbdh = (uk0ahn6nnbba7 == 7'b1010010);
  wire hhf4if064tv59lxifk = (uk0ahn6nnbba7 == 7'b1010011);
  wire gv_izfe7yqh4gkvf76e93ct = (uk0ahn6nnbba7 == 7'b1001011);
  wire hobxt8_ayp1au2dt6zmqdcc = (uk0ahn6nnbba7 == 7'b1001010);
  wire wbsrjrrr8rt_27m9rwnm_ = (uk0ahn6nnbba7 == 7'b1010100);
  wire l9_rbvynoe7x8o0_n_27icr = (uk0ahn6nnbba7 == 7'b1010101);
  wire puc5pybv0exsbi1jenrc = (uk0ahn6nnbba7 == 7'b1011100);
  wire uzvf9tjdfep6fv53xc6uakt = (uk0ahn6nnbba7 == 7'b1011101);
  wire iye23utobc0hah06xcesc14 = (uk0ahn6nnbba7 == 7'b1000111);
  wire tqsbmvgi1q8l40_d8_5 = (uk0ahn6nnbba7 == 7'b1001111);
  wire i3yg5uqgsrfhxxu1pt4o3 = (uk0ahn6nnbba7 == 7'b0110000);
  wire po6ddes535c20_mmy_2u85p = (uk0ahn6nnbba7 == 7'b0111000);
  wire q1g4g81fl48iq3ndywfle3 = (uk0ahn6nnbba7 == 7'b1101010);
  wire a70w9nx14ytij6ok0iq = (uk0ahn6nnbba7 == 7'b1111011);
  wire tgij_tz20n4mlmn8gc = (uk0ahn6nnbba7 == 7'b1101011);



  wire jnhdayjoseb = (ga71__f5g1 == 5'b00000);
  wire l0b5ckml_h1err = (ga71__f5g1 == 5'b00001);
  wire o7pg9yox7y22 = (ga71__f5g1 == 5'b00101);
  wire y2hcqn22lsrsl = (aihiftly == 5'b00000);
  wire e66cg2_0h2b4 = (aihiftly == 5'b00001);
  wire k6belu_b9x2ayw = (aihiftly == 5'b00010);
  wire qkb4tougtjjwxs = (aihiftly == 5'b00011);
  wire adw7hffbin  = (adjmfzwj55ej  == 5'b00000);
  wire szrsuj92ztkk  = (adjmfzwj55ej  == 5'b00001);
  wire lrmd0wxme24  = (adjmfzwj55ej  == 5'b00010);
  wire gu8ts9t4tk1qht  = (adjmfzwj55ej  == 5'b00101);
  wire e_4dvc17j4r_lnf = l0b5ckml_h1err | o7pg9yox7y22; 
  wire omz3uztjy6xo0_l = szrsuj92ztkk | gu8ts9t4tk1qht;   

  wire [5-1:0] u2apzx0s0_ms;
  wire [5-1:0] cyoz2x_qbs1p;
  wire [5-1:0] h_3trq2o2w5gb ;

  wire yv7txmfn9ad8dt = (ag9ylluguwcr == 5'b00000);
  wire y3zkr5mp7y4 = (tbilhd3n1v == 5'b00000);
  wire zczkznydxqjksv  = (z7cl6tvk  == 5'b00000);
  wire lrpfnua6cii2bexrk = (u2apzx0s0_ms == 5'b00001);
  wire ds_ismxbia7ajfooum2 = (u2apzx0s0_ms == 5'b00101);
  wire evab9y_1jyv5cuf0 = (h_3trq2o2w5gb == 5'b00001);
  wire q3cprf7oa8pdc = (h_3trq2o2w5gb == 5'b00101);
  wire m0ra34i4no544w2gpb = lrpfnua6cii2bexrk | ds_ismxbia7ajfooum2; 
  wire qco8v_7vshusc9 = evab9y_1jyv5cuf0 | q3cprf7oa8pdc;   

  wire oezgh2bhqupmgh2 = (ga71__f5g1 == 5'b11111);
  wire sauhc6ef6pqjm_w4 = (aihiftly == 5'b11111);
  wire bgecyjs80sbc  = (adjmfzwj55ej  == 5'b11111);

  wire s3qnk2twp6     = w0s41titqc28jdt & d6r44hi25ixatafeu1 & bfp4chz8bvbs7e8m & ~(o6hnybbrbqkztojg | w__ro7gwx6w331);
  wire id7i5ufppar8     = w0s41titqc28jdt & d6r44hi25ixatafeu1 & bfp4chz8bvbs7e8m &  (o6hnybbrbqkztojg | w__ro7gwx6w331);
  wire g07txhn20bwh3as    = wx_8fko7wy_rmnew7l & d6r44hi25ixatafeu1 & bfp4chz8bvbs7e8m &  ~w__ro7gwx6w331; 
  wire hjxhtr2pfh    = wx_8fko7wy_rmnew7l & d6r44hi25ixatafeu1 & bfp4chz8bvbs7e8m &   w__ro7gwx6w331; 

  wire qwppxd4zz     = sfpsjr_3ucgrnnl4f & d6r44hi25ixatafeu1 & bfp4chz8bvbs7e8m; 
  wire cgfh21c1qcp   = f_575odq4qxl04 & d6r44hi25ixatafeu1 & bfp4chz8bvbs7e8m; 

  wire glv8ztvxphxctm  = w0s41titqc28jdt & cizl6_7mbo_awon & bfp4chz8bvbs7e8m; 
  wire kvnjxxg7anei8786qg = wx_8fko7wy_rmnew7l & cizl6_7mbo_awon & bfp4chz8bvbs7e8m; 
  wire wh7hmrmzlb     = sfpsjr_3ucgrnnl4f & cizl6_7mbo_awon & bfp4chz8bvbs7e8m; 
  wire sa6649too5v5     = f_575odq4qxl04 & cizl6_7mbo_awon & bfp4chz8bvbs7e8m & ezupw6o2yfm5ojugrc3; 

  wire oaeo4esxhvfuvt5j  = w0s41titqc28jdt & vw5it7jugq0nfvd04v & bfp4chz8bvbs7e8m; 
  wire kucqnffs6yyq22tu  = wx_8fko7wy_rmnew7l & vw5it7jugq0nfvd04v & bfp4chz8bvbs7e8m; 
  wire eueft5qh43m7e    = sfpsjr_3ucgrnnl4f & vw5it7jugq0nfvd04v & bfp4chz8bvbs7e8m; 
  wire l4z4jadnl59_a6  = f_575odq4qxl04 & vw5it7jugq0nfvd04v & bfp4chz8bvbs7e8m; 

  wire ifooo477tmr9ucsnr  = w0s41titqc28jdt & bpk53yitybm32g & bfp4chz8bvbs7e8m; 
  wire j3paeay4496m      = wx_8fko7wy_rmnew7l & bpk53yitybm32g & bfp4chz8bvbs7e8m & t8jc64yc1l6q8eclq_c;

  wire rt2gdnok8      = wx_8fko7wy_rmnew7l & bpk53yitybm32g & bfp4chz8bvbs7e8m & w__ro7gwx6w331;

  wire jn7op2_63ozfv    = sfpsjr_3ucgrnnl4f & bpk53yitybm32g & bfp4chz8bvbs7e8m; 
  wire h20g0j2jt      = f_575odq4qxl04 & bpk53yitybm32g & bfp4chz8bvbs7e8m; 

  wire it3sb6rq7z2i67   = w0s41titqc28jdt & asuyn96in9e48ikear_ & bfp4chz8bvbs7e8m; 
  wire v9zbczh8       = wx_8fko7wy_rmnew7l & asuyn96in9e48ikear_ & bfp4chz8bvbs7e8m; 
  wire aiuo7glh4vp0    = sfpsjr_3ucgrnnl4f & asuyn96in9e48ikear_ & bfp4chz8bvbs7e8m; 
  wire sm_lqinid6ej   = f_575odq4qxl04 & asuyn96in9e48ikear_ & bfp4chz8bvbs7e8m; 

  wire ccbtxbyh0qmcdfa    = w0s41titqc28jdt & kn3z45bkwagekkw & bfp4chz8bvbs7e8m; 
  wire hwj750kj      = wx_8fko7wy_rmnew7l & kn3z45bkwagekkw & bfp4chz8bvbs7e8m; 
  wire s04xhr460jiza2  = sfpsjr_3ucgrnnl4f & kn3z45bkwagekkw & bfp4chz8bvbs7e8m; 
  wire hka5a9rzat7j3ku  = f_575odq4qxl04 & kn3z45bkwagekkw & bfp4chz8bvbs7e8m; 

  wire extkhgjdeiqeyj85= w0s41titqc28jdt & cdwv54beu2vbzvh & bfp4chz8bvbs7e8m; 
  wire f8s0zhsklb7tg3m    = wx_8fko7wy_rmnew7l & cdwv54beu2vbzvh & bfp4chz8bvbs7e8m;

  wire h877ps0r0cih1_w_= extkhgjdeiqeyj85;
  wire aug3vtovlhu39z    = f8s0zhsklb7tg3m;

  wire g5vgckumk9u4krx99  = sfpsjr_3ucgrnnl4f & cdwv54beu2vbzvh & bfp4chz8bvbs7e8m; 
  wire ptmaxvmkm2jpf6yl  = f_575odq4qxl04 & cdwv54beu2vbzvh & bfp4chz8bvbs7e8m; 

  wire tdceg4r4ocywxjcsuv     = wgqy37zae8oexwv & mg22fa39qkmi1381_;
  wire yyd3wantj           = wgqy37zae8oexwv & ft758uk96h0lere58vu;
  wire v_a3dq6           = wgqy37zae8oexwv & pw945i12_3q9tpbldo;

  wire d764kpemvglzpk9        = wgqy37zae8oexwv & t3skb9q5zbu_q_fb;
  wire jm6sitcu2sj        = wgqy37zae8oexwv & f9zuwwm5sc91jd4; 


  wire rqj6hf1k9f         = f9k8e7skb6cw2pkw3w & mg22fa39qkmi1381_;
  wire srcanpuv42e7t  = f9k8e7skb6cw2pkw3w & swilkhsvy0ciqh;
  wire e_qxxtaevvw          = 1'b0;
  wire mhz85qp           = f9k8e7skb6cw2pkw3w & ft758uk96h0lere58vu;
  wire br9ybmw_8qr_xw4ojzr = f9k8e7skb6cw2pkw3w & t3skb9q5zbu_q_fb;
  wire ta9huns52lhanjd      = f9k8e7skb6cw2pkw3w & lkhy22ju1fth_z;
  wire ei1me6y0            = f9k8e7skb6cw2pkw3w & atw4jjamnfmexzna29;
  wire tez8bez5l4r         = f9k8e7skb6cw2pkw3w & pw945i12_3q9tpbldo;
  wire zh62ppn61_4yw4         = f9k8e7skb6cw2pkw3w & f9zuwwm5sc91jd4;


  wire w5wv66al4ks3x         = mqwi5z31tkb1fz81y & mg22fa39qkmi1381_;
  wire mbzx7zhsly5         = mqwi5z31tkb1fz81y & ft758uk96h0lere58vu;
  wire lr08s8a1cosklchm4m  = mqwi5z31tkb1fz81y & lkhy22ju1fth_z;
  wire nh22c0jbg5o19         = mqwi5z31tkb1fz81y & pw945i12_3q9tpbldo;

  wire eiqmnomnjfe0      = mqwi5z31tkb1fz81y & t3skb9q5zbu_q_fb;
  wire qi_35cq273ym      = mqwi5z31tkb1fz81y & f9zuwwm5sc91jd4;


  wire sbyhjyyw1          = wgqy37zae8oexwv & swilkhsvy0ciqh;
  wire an_cjmmfv          = wgqy37zae8oexwv & atw4jjamnfmexzna29;
  wire iy0t317_b18b1        = mqwi5z31tkb1fz81y & swilkhsvy0ciqh;
  wire wf8o8lzblge        = mqwi5z31tkb1fz81y & atw4jjamnfmexzna29;

  wire gx2n0dmy9          = 1'b0;
  wire yxd3c1kl5vo15          = 1'b0;
  wire qdqvpvjvmba        = 1'b0;
  wire pfeg45fn01up        = 1'b0;






  wire t61y7hkwkrvm7s = (pq5pe3yehrqxr[6:0] == 7'b1111111);

  wire ww_v_rhq1pd2_fg    = mbzx7zhsly5 & zczkznydxqjksv;
  wire kjzbbod1qt47l8efz    = eiqmnomnjfe0 & zczkznydxqjksv;

  wire cqkv6i9dve          = rqj6hf1k9f  
                         & (~tm0dvbtguid67[12]) & (zczkznydxqjksv) & (y3zkr5mp7y4);

  wire h__4na2w1         = ta9huns52lhanjd  & (tm0dvbtguid67[11:10] == 2'b00);
  wire afnn1is_f9szbi         = ta9huns52lhanjd  & (tm0dvbtguid67[11:10] == 2'b01);
  wire bs3b85ifu         = ta9huns52lhanjd  & (tm0dvbtguid67[11:10] == 2'b10);
  wire pjq11l4lomf3lrph  = ta9huns52lhanjd  & (tm0dvbtguid67[12:10] == 3'b011);

  wire ai1ohlxb9k0vgo1d9      = ta9huns52lhanjd & (tm0dvbtguid67[12:10] == 3'b111) & (tm0dvbtguid67[6:5] == 2'b01); 
  wire cm7ij9pf198f0ifu      = ta9huns52lhanjd & (tm0dvbtguid67[12:10] == 3'b111) & (tm0dvbtguid67[6:5] == 2'b00);

  wire qzjna_8yrjwqibq75b9s = ta9huns52lhanjd & (~h__4na2w1) & (~afnn1is_f9szbi) & (~bs3b85ifu) & (~pjq11l4lomf3lrph) & (~ai1ohlxb9k0vgo1d9) & (~cm7ij9pf198f0ifu);

  wire iw15cor9fq56nb6q3w6   = (tm0dvbtguid67[12] == 1'b0);
  wire l7m0tpckww6nzxyn59cc5w13 = (tm0dvbtguid67[6:2] == 5'b0);

  wire sqhyu61nhtsicrqhpxcwc_4 = 
                 1'b1  
                 ;
  wire x9cbta8yo_b811qozvyp0tqoa =  (w5wv66al4ks3x | h__4na2w1 | afnn1is_f9szbi) & (~sqhyu61nhtsicrqhpxcwc_4);

  wire einxry70u73t166q     = br9ybmw_8qr_xw4ojzr & lrmd0wxme24;
  wire qvq4uyy0b          = br9ybmw_8qr_xw4ojzr & (~lrmd0wxme24);





  wire fy4_5ipo1it2p3xb7 = qvq4uyy0b & (l7m0tpckww6nzxyn59cc5w13 & iw15cor9fq56nb6q3w6);


  wire oa000fsbi9vz2933 = fy4_5ipo1it2p3xb7;

  wire epmy5pkue90oo6im57xozi = tdceg4r4ocywxjcsuv & (iw15cor9fq56nb6q3w6 & zczkznydxqjksv & w0s41titqc28jdt);
  wire kg80830otj0fcd2qp2u90 = einxry70u73t166q & iw15cor9fq56nb6q3w6 & l7m0tpckww6nzxyn59cc5w13; 

  wire tql5edti95od          = pjq11l4lomf3lrph & (tm0dvbtguid67[6:5] == 2'b00);
  wire doq55tb4z          = pjq11l4lomf3lrph & (tm0dvbtguid67[6:5] == 2'b01);
  wire itwlme_oz81a           = pjq11l4lomf3lrph & (tm0dvbtguid67[6:5] == 2'b10);
  wire gzjeu6o0tf4x          = pjq11l4lomf3lrph & (tm0dvbtguid67[6:5] == 2'b11);


  wire w72sj0ys3h3           = lr08s8a1cosklchm4m 
                         & (~tm0dvbtguid67[12]) & (~yv7txmfn9ad8dt) & (y3zkr5mp7y4);
  wire ekodeh8usegq           = lr08s8a1cosklchm4m 
                         & (~tm0dvbtguid67[12]) 

                         & (~y3zkr5mp7y4);
  wire uehd4657vxh53i9q       = lr08s8a1cosklchm4m 
                         & (tm0dvbtguid67[12]) & (zczkznydxqjksv) & (y3zkr5mp7y4);
  wire wgc_484cnth5         = lr08s8a1cosklchm4m 
                         & (tm0dvbtguid67[12]) & (~yv7txmfn9ad8dt) & (y3zkr5mp7y4);
  wire yu0d6pwfl6r          = lr08s8a1cosklchm4m 
                         & (tm0dvbtguid67[12]) 

                         & (~y3zkr5mp7y4);




  wire t6u2o2tra        = (glv8ztvxphxctm | kvnjxxg7anei8786qg | qwppxd4zz | wh7hmrmzlb | eueft5qh43m7e | jn7op2_63ozfv | aiuo7glh4vp0);
  wire i1q5w77apo6kh    = (pq5pe3yehrqxr[26:25] == 2'b00);
  wire l8rbj8208ycy    = (pq5pe3yehrqxr[26:25] == 2'b01);

  wire hschwo70vh36y        = glv8ztvxphxctm  & t8jc64yc1l6q8eclq_c;
  wire bx5js_t0gcoh8        = kvnjxxg7anei8786qg & t8jc64yc1l6q8eclq_c;
  wire gwoe477gldf8c9e    = qwppxd4zz  & i1q5w77apo6kh;
  wire my890tb6fuxn0ar    = wh7hmrmzlb  & i1q5w77apo6kh;
  wire i_43p0nivqch83l   = eueft5qh43m7e & i1q5w77apo6kh;
  wire lg8nys4yk9hgun1   = jn7op2_63ozfv & i1q5w77apo6kh;
  wire fz4uie4yxvn5     = lrptc0hyjyd7hdoypa0_g & aiuo7glh4vp0;
  wire snxdp3tvw7a     = mso_1l7nnv4ac14pv6qh & aiuo7glh4vp0;
  wire x0c94xeqpc8nzim7     = e9hn3j9k88f8miq238hz1 & aiuo7glh4vp0;
  wire kzyiyt0xi8d     = duf6qt_vm6jkmkv9xu9 & aiuo7glh4vp0;
  wire o4tc3g036bgoap    = gu_2fhfulrttqq4e_fiax & aiuo7glh4vp0;
  wire nlb5566a2kkzrak    = i6fh1oflvwwzfgicny1c & aiuo7glh4vp0 & ezupw6o2yfm5ojugrc3;
  wire t82iq62ywf1u_5   = i6fh1oflvwwzfgicny1c & aiuo7glh4vp0 & d24iqtxvb2trplxk2m;
  wire byqkkp26xdsszd   = i6fh1oflvwwzfgicny1c & aiuo7glh4vp0 & t8jc64yc1l6q8eclq_c;
  wire vzgrcege9g3qyat     = f6kcevztmpqpnc8xp3_r4 & aiuo7glh4vp0 & ezupw6o2yfm5ojugrc3;
  wire p0u65_oip3cn     = f6kcevztmpqpnc8xp3_r4 & aiuo7glh4vp0 & d24iqtxvb2trplxk2m;
  wire iz_sm_7y_ixfw1btmz  = l6zyb5b3_f8uuon8o3p & aiuo7glh4vp0 & y2hcqn22lsrsl;
  wire uz6maeeehzsn6uzwxk = l6zyb5b3_f8uuon8o3p & aiuo7glh4vp0 & e66cg2_0h2b4;
  wire gkj8ltdpe4tcqini4h   = k_h8qestuhin60n5ckxmkfx & aiuo7glh4vp0 & ezupw6o2yfm5ojugrc3;
  wire qfgkmomxjwhe      = c7npl5770szduubj6_grim & aiuo7glh4vp0 & t8jc64yc1l6q8eclq_c;
  wire v3he_44ycy65      = c7npl5770szduubj6_grim & aiuo7glh4vp0 & d24iqtxvb2trplxk2m;
  wire h5gjvo_bpoph5i      = c7npl5770szduubj6_grim & aiuo7glh4vp0 & ezupw6o2yfm5ojugrc3;
  wire l6qpfpq3ro_9gr   = k_h8qestuhin60n5ckxmkfx & aiuo7glh4vp0 & d24iqtxvb2trplxk2m;
  wire dywxta8oxdnj1q9i0d  = tx0e46vrruq3cgq9ghul4 & aiuo7glh4vp0 & y2hcqn22lsrsl;
  wire zqz28qv7052ajkf7 = tx0e46vrruq3cgq9ghul4 & aiuo7glh4vp0 & e66cg2_0h2b4;
  wire nxf52k3xp6im5o6p3   = v3hylq_n52mziras6qen & aiuo7glh4vp0;
  wire hx05sow34f5nxv  = l6zyb5b3_f8uuon8o3p & aiuo7glh4vp0 & k6belu_b9x2ayw;
  wire iboby_h0cqqucgnxw = l6zyb5b3_f8uuon8o3p & aiuo7glh4vp0 & qkb4tougtjjwxs;
  wire nu4l8_3i80k9r9huos  = tx0e46vrruq3cgq9ghul4 & aiuo7glh4vp0 & k6belu_b9x2ayw;
  wire wjhbw3uh3oljyutu2gel = tx0e46vrruq3cgq9ghul4 & aiuo7glh4vp0 & qkb4tougtjjwxs;

  wire hh5s1lrugs7        = 1'b0;
  wire wcsiqmn9v7po        = 1'b0;
  wire y1x6fpss6_6        = glv8ztvxphxctm  & w__ro7gwx6w331;
  wire hh5fb5xzanf14        = kvnjxxg7anei8786qg & w__ro7gwx6w331;
  wire j_tdnombv0p5jwn8    = qwppxd4zz  & l8rbj8208ycy;
  wire rog98nkwfh96pgah1    = wh7hmrmzlb  & l8rbj8208ycy;
  wire ryz5m33fgnp6ofcw   = eueft5qh43m7e & l8rbj8208ycy;
  wire ig6dxpy3sgfnd   = jn7op2_63ozfv & l8rbj8208ycy;
  wire knc4udhhcbv     = t6_6ypj94nny67ise0x9 & aiuo7glh4vp0;
  wire vou4ap3g4kukvz7a     = xfrai8f3331hb4z5ww5_ & aiuo7glh4vp0;
  wire ou19p6zx65a     = pvy429fepo5d_7j0eq5ky & aiuo7glh4vp0;
  wire lz1544702tkg0u     = cvhx1ne2we07dkbzbpwakl & aiuo7glh4vp0;
  wire cbru05_q5bm7    = k3sfqtpqynzqda4xtugl4 & aiuo7glh4vp0;
  wire vdmyb8x4qmwi7on2    = i0ahgxc7hvmvc1hsbq8 & aiuo7glh4vp0 & ezupw6o2yfm5ojugrc3;
  wire tfoxw8ia_xdt0   = i0ahgxc7hvmvc1hsbq8 & aiuo7glh4vp0 & d24iqtxvb2trplxk2m;
  wire f128ccj13txxdwpl   = i0ahgxc7hvmvc1hsbq8 & aiuo7glh4vp0 & t8jc64yc1l6q8eclq_c;
  wire hjq039vacscr     = toaowsb_5w3arwmyl2 & aiuo7glh4vp0 & ezupw6o2yfm5ojugrc3;
  wire n6f1xma1ku0cqc9     = toaowsb_5w3arwmyl2 & aiuo7glh4vp0 & d24iqtxvb2trplxk2m;
  wire tnkhekmenrbyvq  = bepkj4gbb77isq3_v9 & aiuo7glh4vp0 & e66cg2_0h2b4;
  wire gsqes4kpzyh7s4  = uncepq376ovruspfffvl5 & aiuo7glh4vp0 & y2hcqn22lsrsl;
  wire ns2ccb8p4kf3o      = whvtopzve8q_t001lyx & aiuo7glh4vp0 & t8jc64yc1l6q8eclq_c;
  wire wy5oiwkuovruvc      = whvtopzve8q_t001lyx & aiuo7glh4vp0 & d24iqtxvb2trplxk2m;
  wire mtnmu5bzb5z9      = whvtopzve8q_t001lyx & aiuo7glh4vp0 & ezupw6o2yfm5ojugrc3;
  wire u72qi7gmhj37d_h5c   = eu9j7rkhrocfjsewdf6mfvu & aiuo7glh4vp0 & y2hcqn22lsrsl & d24iqtxvb2trplxk2m;
  wire th_rx8vbgu0ydrx  = c9xaw73uh3hmihrn801brf & aiuo7glh4vp0 & y2hcqn22lsrsl;
  wire glahkq0rwcrj086j7k1j = c9xaw73uh3hmihrn801brf & aiuo7glh4vp0 & e66cg2_0h2b4;
  wire i_oja_fou8xg9_  = mnd8c7lvcdtsypyiygspg & aiuo7glh4vp0 & y2hcqn22lsrsl;
  wire jz2t1e591yva8m5 = mnd8c7lvcdtsypyiygspg & aiuo7glh4vp0 & e66cg2_0h2b4;
  wire knqkb_9b7915rg  = c9xaw73uh3hmihrn801brf & aiuo7glh4vp0 & k6belu_b9x2ayw;
  wire jlez7xntekztmffn06 = c9xaw73uh3hmihrn801brf & aiuo7glh4vp0 & qkb4tougtjjwxs;
  wire q1mnx00q446iezuqt  = mnd8c7lvcdtsypyiygspg & aiuo7glh4vp0 & k6belu_b9x2ayw;
  wire bvcgz8q5ffa32w7 = mnd8c7lvcdtsypyiygspg & aiuo7glh4vp0 & qkb4tougtjjwxs;
  wire va7j9_tx3li0xd   = eu9j7rkhrocfjsewdf6mfvu & aiuo7glh4vp0 & ezupw6o2yfm5ojugrc3 & ezupw6o2yfm5ojugrc3;
  wire tr03xi8fsjspsc   = rf284mrjg_bqa1hj60swyf & aiuo7glh4vp0 & ezupw6o2yfm5ojugrc3 & ezupw6o2yfm5ojugrc3;



  wire j19mr32tje7z      = cgfh21c1qcp & ezupw6o2yfm5ojugrc3;
  wire z_nqw2ea      = cgfh21c1qcp & d24iqtxvb2trplxk2m;
  wire i9jg2q2v0e9q      = cgfh21c1qcp & d0jauc9xnvhr53rq3;
  wire ofqth0x0_ej20      = cgfh21c1qcp & tcks0htkit9weu;
  wire mips8_vh9     = cgfh21c1qcp & o6hnybbrbqkztojg;
  wire ybsdpobpotarp     = cgfh21c1qcp & dwe8qnpoudm94xa;

  wire w15cfmvs_rdfsulo = cgfh21c1qcp & (
                     ~(j19mr32tje7z  |
                       z_nqw2ea  |
                       i9jg2q2v0e9q  |
                       ofqth0x0_ej20  |
                       mips8_vh9 |
                       ybsdpobpotarp )
                     );


  wire rlra2ebf_s      = 1'b0;
  wire j3wz5of15zrkr      = 1'b0;
  wire x47d8y9qh7l     = 1'b0;
  wire jq0ukfw42dsg0     = 1'b0;
  wire k0glq1z9c20ujfyc = 1'b0;
  wire [6:0] w4jk48u5zmn7 = 7'b0;
  wire [64-1:0] e2rml0d5xlemgdqf2a = 64'b0;



  wire cr12wtja7cvr    = sm_lqinid6ej & ezupw6o2yfm5ojugrc3 & (pq5pe3yehrqxr[31:20] == 12'b0000_0000_0000);
  wire obb913ycps11   = sm_lqinid6ej & ezupw6o2yfm5ojugrc3 & (pq5pe3yehrqxr[31:20] == 12'b0000_0000_0001);
  wire f5xtf96mnbjz     = sm_lqinid6ej & ezupw6o2yfm5ojugrc3 & (pq5pe3yehrqxr[31:20] == 12'b0011_0000_0010);
  wire h9l8g_opcyz48     = sm_lqinid6ej & ezupw6o2yfm5ojugrc3 & (pq5pe3yehrqxr[31:20] == 12'b0001_0000_0010);
  wire d4r5ikwsk     = sm_lqinid6ej & ezupw6o2yfm5ojugrc3 & (pq5pe3yehrqxr[31:20] == 12'b0111_1011_0010);
  wire rbt2ovi_6h      = sm_lqinid6ej & ezupw6o2yfm5ojugrc3 & (pq5pe3yehrqxr[31:20] == 12'b0001_0000_0101);


  wire zziyl6t8rs22kz2    = sm_lqinid6ej & d24iqtxvb2trplxk2m; 
  wire fb2hmea7xsh48i    = sm_lqinid6ej & t8jc64yc1l6q8eclq_c; 
  wire k7_rcb9pbl    = sm_lqinid6ej & w__ro7gwx6w331; 
  wire nt0rwqyh45801   = sm_lqinid6ej & tcks0htkit9weu; 
  wire ae9uh2qsyem1utk9   = sm_lqinid6ej & o6hnybbrbqkztojg; 
  wire vv6pnkge7dhr1ay_   = sm_lqinid6ej & dwe8qnpoudm94xa; 

  wire cicq2g9r_bh93 ;
  wire rb8rv_jwet5lap0p = sm_lqinid6ej  & (~
                         ( cr12wtja7cvr  |
                           obb913ycps11 |
                           f5xtf96mnbjz   |
                           d4r5ikwsk   |
                           h9l8g_opcyz48   |
                           cicq2g9r_bh93 |
                           rbt2ovi_6h    |
                           zziyl6t8rs22kz2  |
                           fb2hmea7xsh48i  |
                           k7_rcb9pbl  |
                           nt0rwqyh45801 |
                           ae9uh2qsyem1utk9 |
                           vv6pnkge7dhr1ay_ ));



  wire g0rwtpabeiisocfnwg = d4r5ikwsk & (~bktu0z1mk56);
  wire v91kaxeokzy6fv5 = f5xtf96mnbjz & (~u2k4dyp52s_m);
  wire r773brf2qafg123x   = h9l8g_opcyz48 & (~u2k4dyp52s_m) & (~djvj1e_ | (djvj1e_ & b0ry73kp6sc2)); 
  wire ebxkh3mj83gh00a86o_rb = cicq2g9r_bh93 & (~u2k4dyp52s_m) & (~djvj1e_ | (djvj1e_ & cz1hh6af7xp2)); 
  wire nh5pz0qwy9ffo2l1  = (pq5pe3yehrqxr[31:20] == 12'h180);
  wire r1pa5yctc1vd7e650n    = q1coyps2cz7xe & nh5pz0qwy9ffo2l1 & (~u2k4dyp52s_m) & (djvj1e_ & cz1hh6af7xp2);
  wire plr5quy6x6fvmq27ye    = rbt2ovi_6h & (~u2k4dyp52s_m) & (~djvj1e_ | (djvj1e_ & hr64e6c3gy));

  wire waejh__hl02blsw4eau2ir6332zz = sm_lqinid6ej & ezupw6o2yfm5ojugrc3
                                   & (~cicq2g9r_bh93)
                                   ;
  wire fpfh9sb3          = sm_lqinid6ej & (~ezupw6o2yfm5ojugrc3);





  assign o8rwk067     = h20g0j2jt    | e_qxxtaevvw  | ei1me6y0;
  assign r1on2k03r    = sa6649too5v5   | wgc_484cnth5 | w72sj0ys3h3;
  assign gw7452ctd577    = (h20g0j2jt & omz3uztjy6xo0_l) | e_qxxtaevvw
                     | (sa6649too5v5 & omz3uztjy6xo0_l & (~e_4dvc17j4r_lnf))
                     | (sa6649too5v5 & omz3uztjy6xo0_l & e_4dvc17j4r_lnf)
                     | wgc_484cnth5 
                     ;

  assign b1roq8tr9r     = (sa6649too5v5 & (~omz3uztjy6xo0_l) & e_4dvc17j4r_lnf)
                     | (sa6649too5v5 & omz3uztjy6xo0_l & e_4dvc17j4r_lnf &( adjmfzwj55ej != ga71__f5g1))
                     | (wgc_484cnth5 & m0ra34i4no544w2gpb)
                     | (w72sj0ys3h3 & m0ra34i4no544w2gpb)
                     ;

  assign j_ku88w81rg     = cgfh21c1qcp | tez8bez5l4r | zh62ppn61_4yw4
                     ;
  assign ld01d40_n3     = o8rwk067 | r1on2k03r | j_ku88w81rg;




  wire x0x8nq83jfrfkw14;
  wire zl2hdo5flk_x  ;
  wire l143yo227i5fe5s3;
  wire dw61vkalbiqitxbxy8n0;
  assign jw1vgacy_r0vr  = f5xtf96mnbjz | d4r5ikwsk
                     | x0x8nq83jfrfkw14 
                     | rbt2ovi_6h
                     | l143yo227i5fe5s3
                     | h9l8g_opcyz48
                     | cicq2g9r_bh93
                     ; 

  wire khaw8p = ld01d40_n3 | f5xtf96mnbjz | d4r5ikwsk  | dw61vkalbiqitxbxy8n0
              | h9l8g_opcyz48
              | cicq2g9r_bh93 
                ;

  wire [34-1:0] loymwnjzrl_cl;
  assign loymwnjzrl_cl[3:0    ]    = 4'd3;
  assign loymwnjzrl_cl[4:4   ]    = vlfahv69;
  assign loymwnjzrl_cl[5:5 ]  = o8rwk067;
  assign loymwnjzrl_cl[6:6]  = r1on2k03r;
  assign loymwnjzrl_cl[7:7]  = gw7452ctd577;
  assign loymwnjzrl_cl[8:8]   = b1roq8tr9r;
  assign loymwnjzrl_cl[9:9]  = qhyq467foflgyn5y;
  assign loymwnjzrl_cl[10:10  ]  = j19mr32tje7z | tez8bez5l4r;
  assign loymwnjzrl_cl[11:11  ]  = z_nqw2ea | zh62ppn61_4yw4;
  assign loymwnjzrl_cl[12:12  ]  = i9jg2q2v0e9q; 
  assign loymwnjzrl_cl[13:13  ]  = ofqth0x0_ej20 ;
  assign loymwnjzrl_cl[14:14 ]  = mips8_vh9;
  assign loymwnjzrl_cl[15:15 ]  = ybsdpobpotarp;
  assign loymwnjzrl_cl[16:16  ]  = j_ku88w81rg;
  assign loymwnjzrl_cl[17:17 ]  = f5xtf96mnbjz;
  assign loymwnjzrl_cl[19:19 ]  = d4r5ikwsk;
  assign loymwnjzrl_cl[20:20 ] = zl2hdo5flk_x;
  assign loymwnjzrl_cl[21:21] = l143yo227i5fe5s3;
  assign loymwnjzrl_cl[18:18 ]  = h9l8g_opcyz48;
  assign loymwnjzrl_cl[22:22] = cicq2g9r_bh93;
  assign loymwnjzrl_cl[23:23  ]  = rlra2ebf_s ;
  assign loymwnjzrl_cl[24:24  ]  = j3wz5of15zrkr ;
  assign loymwnjzrl_cl[25:25 ]  = x47d8y9qh7l;
  assign loymwnjzrl_cl[26:26 ]  = jq0ukfw42dsg0;
  assign loymwnjzrl_cl[33:27 ]  = w4jk48u5zmn7;




  wire u3oqktpp24ks4o     = (it3sb6rq7z2i67 & ezupw6o2yfm5ojugrc3)
                       ;
  wire kzy4s9z4ai2     = it3sb6rq7z2i67 & t8jc64yc1l6q8eclq_c;
  wire g5b6upa17uxdlc    = it3sb6rq7z2i67 & w__ro7gwx6w331;
  wire lu5f0x53z3m1     = it3sb6rq7z2i67 & d0jauc9xnvhr53rq3;
  wire y0wv1q1ravs4      = it3sb6rq7z2i67 & o6hnybbrbqkztojg;
  wire vh5zm21snh5hzb     = it3sb6rq7z2i67 & dwe8qnpoudm94xa;

  wire hx9u53hfqb     = it3sb6rq7z2i67 & d24iqtxvb2trplxk2m & (pq5pe3yehrqxr[31:26] == 6'b000000);
  wire pr4pv6nch2d     = it3sb6rq7z2i67 & tcks0htkit9weu & (pq5pe3yehrqxr[31:26] == 6'b000000);
  wire fgao9da88hto     = it3sb6rq7z2i67 & tcks0htkit9weu & (pq5pe3yehrqxr[31:26] == 6'b010000);

  wire piay0j_yijhago5y = it3sb6rq7z2i67 & ((tcks0htkit9weu & (~pr4pv6nch2d) & (~fgao9da88hto))
                                       | (d24iqtxvb2trplxk2m & (~hx9u53hfqb)) 
                                      );




  wire icw85efsw91jj    = h877ps0r0cih1_w_ & ezupw6o2yfm5ojugrc3;
  wire nk_7dsag_1qmj_    = h877ps0r0cih1_w_ & d24iqtxvb2trplxk2m & lrptc0hyjyd7hdoypa0_g;
  wire b4q7v3qyhprrukx    = h877ps0r0cih1_w_ & tcks0htkit9weu & lrptc0hyjyd7hdoypa0_g;
  wire ex08mtx1kg0    = h877ps0r0cih1_w_ & tcks0htkit9weu & bepkj4gbb77isq3_v9;

  wire coj7bezvnp6c5iibk0vvtu9 = h877ps0r0cih1_w_ & (~icw85efsw91jj) & (~nk_7dsag_1qmj_) & (~b4q7v3qyhprrukx) & (~ex08mtx1kg0);

  wire qu5h2fm8yi0cxb012s8_t9he = (pq5pe3yehrqxr[25] == 1'b0); 
  wire cyv0hhf3man9exnii4w2qrs = (nk_7dsag_1qmj_ | b4q7v3qyhprrukx | ex08mtx1kg0) & (~qu5h2fm8yi0cxb012s8_t9he);


  wire cwbhrq_h8      = v9zbczh8     & ezupw6o2yfm5ojugrc3 & lrptc0hyjyd7hdoypa0_g;
  wire e7e81dk96      = v9zbczh8     & ezupw6o2yfm5ojugrc3 & bepkj4gbb77isq3_v9;
  wire pwhj91c5h1ot4      = v9zbczh8     & d24iqtxvb2trplxk2m & lrptc0hyjyd7hdoypa0_g;
  wire schh4eesozj      = v9zbczh8     & t8jc64yc1l6q8eclq_c & lrptc0hyjyd7hdoypa0_g;
  wire m064pbifqkhsci     = v9zbczh8     & w__ro7gwx6w331 & lrptc0hyjyd7hdoypa0_g;
  wire ztgds1_2j1d      = v9zbczh8     & d0jauc9xnvhr53rq3 & lrptc0hyjyd7hdoypa0_g;
  wire dxwwmywt_      = v9zbczh8     & tcks0htkit9weu & lrptc0hyjyd7hdoypa0_g;
  wire jj4t0lhdb3l      = v9zbczh8     & tcks0htkit9weu & bepkj4gbb77isq3_v9;
  wire czthwvotcy1       = v9zbczh8     & o6hnybbrbqkztojg & lrptc0hyjyd7hdoypa0_g;
  wire pb3evqkebz      = v9zbczh8     & dwe8qnpoudm94xa & lrptc0hyjyd7hdoypa0_g;




  wire hdnmwh5v_     = aug3vtovlhu39z & ezupw6o2yfm5ojugrc3 & lrptc0hyjyd7hdoypa0_g;
  wire aa_ozibgfdhwo     = aug3vtovlhu39z & ezupw6o2yfm5ojugrc3 & bepkj4gbb77isq3_v9;

  wire ygydsp9lq5u5li     = aug3vtovlhu39z & d24iqtxvb2trplxk2m & lrptc0hyjyd7hdoypa0_g;
  wire qn4sshj3ct9     = aug3vtovlhu39z & tcks0htkit9weu & lrptc0hyjyd7hdoypa0_g;
  wire z05l25nz8     = aug3vtovlhu39z & tcks0htkit9weu & bepkj4gbb77isq3_v9;



  wire a6x0kl79q36      = v9zbczh8     & ezupw6o2yfm5ojugrc3 & t6_6ypj94nny67ise0x9;
  wire jgncnwo8lu01     = v9zbczh8     & d24iqtxvb2trplxk2m & t6_6ypj94nny67ise0x9;
  wire g_oka7qgfr5inx   = v9zbczh8     & t8jc64yc1l6q8eclq_c & t6_6ypj94nny67ise0x9;
  wire zswqi_bpr6dj    = v9zbczh8     & w__ro7gwx6w331 & t6_6ypj94nny67ise0x9;
  wire lpac9vygdosz      = v9zbczh8     & d0jauc9xnvhr53rq3 & t6_6ypj94nny67ise0x9;
  wire gu1ryj7evsze     = v9zbczh8     & tcks0htkit9weu & t6_6ypj94nny67ise0x9;
  wire ujvx9ip2      = v9zbczh8     & o6hnybbrbqkztojg & t6_6ypj94nny67ise0x9;
  wire ph174i8mt     = v9zbczh8     & dwe8qnpoudm94xa & t6_6ypj94nny67ise0x9;


  wire m_5r0ivgcn     = aug3vtovlhu39z  & ezupw6o2yfm5ojugrc3 & t6_6ypj94nny67ise0x9;
  wire vjyxyga4yc     = aug3vtovlhu39z  & d0jauc9xnvhr53rq3 & t6_6ypj94nny67ise0x9;
  wire veznwo9f7pzr    = aug3vtovlhu39z  & tcks0htkit9weu & t6_6ypj94nny67ise0x9;
  wire re57g9q8nl7bu     = aug3vtovlhu39z  & o6hnybbrbqkztojg & t6_6ypj94nny67ise0x9;
  wire cwupd7pgtwtjh    = aug3vtovlhu39z  & dwe8qnpoudm94xa & t6_6ypj94nny67ise0x9;


  wire elg6c3h_r04v5e71 = v9zbczh8 & (
                          ~(cwbhrq_h8   |
                            e7e81dk96   |
                            pwhj91c5h1ot4   |
                            schh4eesozj   |
                            m064pbifqkhsci  |
                            ztgds1_2j1d   |
                            dxwwmywt_   |
                            jj4t0lhdb3l   |
                            czthwvotcy1    |
                            pb3evqkebz   |

                            a6x0kl79q36   |
                            jgncnwo8lu01  |
                            g_oka7qgfr5inx|
                            zswqi_bpr6dj |
                            lpac9vygdosz   |
                            gu1ryj7evsze  |
                            ujvx9ip2   |
                            ph174i8mt  ));


  wire wa2rqb81bsgzs2g9adv = aug3vtovlhu39z & (
                                ~(hdnmwh5v_     |
                                  aa_ozibgfdhwo     |
                                  ygydsp9lq5u5li     |
                                  qn4sshj3ct9     |
                                  z05l25nz8     |

                                  m_5r0ivgcn     |
                                  vjyxyga4yc     |
                                  veznwo9f7pzr    |
                                  re57g9q8nl7bu     |
                                  cwupd7pgtwtjh    ));


  wire y4jtark0b_      = u3oqktpp24ks4o & jnhdayjoseb & adw7hffbin & (~(|pq5pe3yehrqxr[31:20])) 
                       ;

  assign x0x8nq83jfrfkw14 = cr12wtja7cvr | obb913ycps11 | uehd4657vxh53i9q;

  wire iokgk17mtvv7q9 = 1'b0;
  wire c_rxvcxopqt04e = 1'b0;
  wire [4:0] g0j_spv4odvr_ti_b = 5'b0;
  wire [4:0] peii_nky7f5_kkx3rj = 5'b0;

  wire jt89qnb7dg1f2yn   = 1'b0;
  wire h88nna043n7xx5claa8 = 1'b0;
  wire dwq5k2lv41hzl4uo = 1'b0;
  wire nqyi2a2r4nlo07ttm = 1'b0;
  wire rc60cnq6vhfqgj5     = 1'b0;
  wire p4c0hz04wynm2g_cm1r1 = 1'b0;
  wire u4z875qi66188zvw  = 1'b0;
  wire zu05kaer_n3ghc18wt  = 1'b0;

  wire ei82smlw45m = 
              ( it3sb6rq7z2i67
              | v9zbczh8 & (~t6_6ypj94nny67ise0x9) 
              | ccbtxbyh0qmcdfa
              | hwj750kj
              | tdceg4r4ocywxjcsuv
              | rqj6hf1k9f         
              | br9ybmw_8qr_xw4ojzr 
              | mhz85qp | ekodeh8usegq
              | w5wv66al4ks3x         
              | ta9huns52lhanjd  
              | yu0d6pwfl6r
              | cqkv6i9dve | y4jtark0b_
              | rbt2ovi_6h 
              | x0x8nq83jfrfkw14)
              | h877ps0r0cih1_w_
              | aug3vtovlhu39z & (~t6_6ypj94nny67ise0x9) 
              | srcanpuv42e7t
              | ai1ohlxb9k0vgo1d9
              ;

  wire hqkcyoh04f5d5j = ei82smlw45m & (~rbt2ovi_6h) & (~x0x8nq83jfrfkw14)
                        ;

  wire qt8cr87lzx1u;
  wire [47-1:0] deq9tleqxy3fq;
  assign deq9tleqxy3fq[3:0    ]    = 4'd1;
  assign deq9tleqxy3fq[4:4   ]    = vlfahv69;
  assign deq9tleqxy3fq[5:5]    = cwbhrq_h8  | u3oqktpp24ks4o | ccbtxbyh0qmcdfa |
                                                  tdceg4r4ocywxjcsuv | rqj6hf1k9f | einxry70u73t166q | yu0d6pwfl6r |


                                                  mhz85qp | ekodeh8usegq;
  assign deq9tleqxy3fq[6:6]    = e7e81dk96  | tql5edti95od ;      
  assign deq9tleqxy3fq[13:13]    = schh4eesozj  | kzy4s9z4ai2;     
  assign deq9tleqxy3fq[14:14]   = m064pbifqkhsci | g5b6upa17uxdlc;  
  assign deq9tleqxy3fq[7:7]    = ztgds1_2j1d  | lu5f0x53z3m1 | doq55tb4z;    
  assign deq9tleqxy3fq[8:8]    = pwhj91c5h1ot4  | hx9u53hfqb | w5wv66al4ks3x;   
  assign deq9tleqxy3fq[9:9]    = dxwwmywt_  | pr4pv6nch2d | h__4na2w1;
  assign deq9tleqxy3fq[10:10]    = jj4t0lhdb3l  | fgao9da88hto | afnn1is_f9szbi;   
  assign deq9tleqxy3fq[11:11 ]    = czthwvotcy1   | y0wv1q1ravs4  | itwlme_oz81a;     
  assign deq9tleqxy3fq[12:12]    = pb3evqkebz  | vh5zm21snh5hzb | bs3b85ifu | gzjeu6o0tf4x;
  assign deq9tleqxy3fq[15:15]    = hwj750kj  | qvq4uyy0b; 
  assign deq9tleqxy3fq[16:16] = qt8cr87lzx1u; 
  assign deq9tleqxy3fq[17:17 ] = ccbtxbyh0qmcdfa;
  assign deq9tleqxy3fq[18:18 ]   = cqkv6i9dve | y4jtark0b_;
  assign deq9tleqxy3fq[19:19 ]  = cr12wtja7cvr; 
  assign deq9tleqxy3fq[20:20 ]  = obb913ycps11 | uehd4657vxh53i9q;
  assign deq9tleqxy3fq[21:21  ]  = rbt2ovi_6h;
  assign deq9tleqxy3fq[22:22] = 1'b0;
  assign deq9tleqxy3fq[23:23  ] = iokgk17mtvv7q9;
  assign deq9tleqxy3fq[24:24  ] = c_rxvcxopqt04e;
  assign deq9tleqxy3fq[29:25 ] = g0j_spv4odvr_ti_b;
  assign deq9tleqxy3fq[34:30 ] = peii_nky7f5_kkx3rj;
  assign deq9tleqxy3fq[35:35 ] = h88nna043n7xx5claa8;
  assign deq9tleqxy3fq[36:36 ] = dwq5k2lv41hzl4uo;
  assign deq9tleqxy3fq[37:37 ] = nqyi2a2r4nlo07ttm;
  assign deq9tleqxy3fq[38:38     ] = rc60cnq6vhfqgj5    ;
  assign deq9tleqxy3fq[39:39 ] = p4c0hz04wynm2g_cm1r1;
  assign deq9tleqxy3fq[40:40  ] = u4z875qi66188zvw ;
  assign deq9tleqxy3fq[41:41  ] = zu05kaer_n3ghc18wt ;
  assign deq9tleqxy3fq[42:42 ]  = hdnmwh5v_ | icw85efsw91jj | ai1ohlxb9k0vgo1d9 | srcanpuv42e7t;
  assign deq9tleqxy3fq[43:43 ]  = aa_ozibgfdhwo | cm7ij9pf198f0ifu;
  assign deq9tleqxy3fq[44:44 ]  = ygydsp9lq5u5li | nk_7dsag_1qmj_;
  assign deq9tleqxy3fq[45:45 ]  = qn4sshj3ct9 | b4q7v3qyhprrukx;
  assign deq9tleqxy3fq[46:46 ]  = z05l25nz8 | ex08mtx1kg0;


  wire aw5pbsduwvhyhb3aka  = u2k4dyp52s_m & (nt0rwqyh45801) & (pq5pe3yehrqxr[31:20] == 12'h7EB);
  wire jbkjansoihuv2nv     = u2k4dyp52s_m & (nt0rwqyh45801) & (pq5pe3yehrqxr[31:20] == 12'h7EE);
  wire ql2xoldgv6si0j      = u2k4dyp52s_m & (nt0rwqyh45801) & (pq5pe3yehrqxr[31:20] == 12'h7EF);
  wire u_mgu2iomgss4kbb5q = (jbkjansoihuv2nv | ql2xoldgv6si0j | aw5pbsduwvhyhb3aka); 
  wire wqpng9lj3ibxslk       = (u2k4dyp52s_m | djvj1e_) & (nt0rwqyh45801) & (pq5pe3yehrqxr[31:20] == 12'h949);
  wire o2zokol469i9emxjt        = (u2k4dyp52s_m | djvj1e_) & (nt0rwqyh45801) & (pq5pe3yehrqxr[31:20] == 12'h94a);
  wire no5vijin9fx5kyxd3lop2wg4d = (wqpng9lj3ibxslk | o2zokol469i9emxjt); 

  wire a7bzgrh = fpfh9sb3 
                & (~u_mgu2iomgss4kbb5q)
                & (~no5vijin9fx5kyxd3lop2wg4d)
              ;
  assign rphjsg75001l2 = a7bzgrh & (  (pq5pe3yehrqxr[31:20] == 12'h001) 
                          || (pq5pe3yehrqxr[31:20] == 12'h002) 
                          || (pq5pe3yehrqxr[31:20] == 12'h003)
                          );

  assign hgvdw0qnels8 = a7bzgrh & (  (pq5pe3yehrqxr[31:20] == 12'h801));









  wire [27-1:0] krezi5k4lo8g;
  assign krezi5k4lo8g[3:0    ]    = 4'd4;
  assign krezi5k4lo8g[4:4   ]    = vlfahv69;
  assign krezi5k4lo8g[5:5 ] = zziyl6t8rs22kz2 | nt0rwqyh45801; 
  assign krezi5k4lo8g[6:6 ] = fb2hmea7xsh48i | ae9uh2qsyem1utk9;
  assign krezi5k4lo8g[7:7 ] = k7_rcb9pbl | vv6pnkge7dhr1ay_;
  assign krezi5k4lo8g[8:8] = nt0rwqyh45801 | ae9uh2qsyem1utk9 | vv6pnkge7dhr1ay_;
  assign krezi5k4lo8g[13:9 ] = ga71__f5g1;
  assign krezi5k4lo8g[14:14] = jnhdayjoseb;
  assign krezi5k4lo8g[26:15] = pq5pe3yehrqxr[31:20];




  assign zl2hdo5flk_x    = ifooo477tmr9ucsnr & ezupw6o2yfm5ojugrc3;
  assign l143yo227i5fe5s3  = ifooo477tmr9ucsnr & d24iqtxvb2trplxk2m;
  assign cicq2g9r_bh93    = sm_lqinid6ej & ezupw6o2yfm5ojugrc3 & pvy429fepo5d_7j0eq5ky;


  assign dw61vkalbiqitxbxy8n0  = zl2hdo5flk_x | l143yo227i5fe5s3;

  
  
  
  
  wire qfrdiaxh3i3k     = pq5pe3yehrqxr[24];
  wire x3m205i475_nt098cv   = (qfrdiaxh3i3k == 1'b0);
  wire km4hjrsbw2uxh2_qt   = (qfrdiaxh3i3k == 1'b1);
  
  wire [1:0] t2hwvtrrr2t1c53     = pq5pe3yehrqxr[24:23];
  wire r70hhozfmlgd3eqafzt  = (t2hwvtrrr2t1c53 == 2'b00);
  wire kis_u1bo6hhg_7rlffxs  = (t2hwvtrrr2t1c53 == 2'b01);
  wire cgtj86qjqc4whb8p2jo  = (t2hwvtrrr2t1c53 == 2'b10);
  
  wire [4:0] xfkngdj3jaifg = pq5pe3yehrqxr[24:20];

  wire asvcpbvzr7u9gfqr_hlh68 = (xfkngdj3jaifg == 5'b01000);           
  wire kre86u005m4jj77idkd170 = (xfkngdj3jaifg == 5'b01001);           
  wire h6jjzsxi8aw0us788h = (xfkngdj3jaifg == 5'b01010);           
  wire yswws2ff7bkbvaic3it7g = (xfkngdj3jaifg == 5'b01011);           
  wire yc8o21itzjuxfoo_32 = (xfkngdj3jaifg == 5'b10011);           
  wire z1_re9ax86eago99v6ic1ke = (xfkngdj3jaifg == 5'b01100);           
  wire yiprb7xpgx9hgyddnxoh = (xfkngdj3jaifg == 5'b01101);           
  wire hutky_0znezwi4oz7cs = (xfkngdj3jaifg == 5'b01110);           
  wire fe7237ktiiy1d5p48dam8 = (xfkngdj3jaifg == 5'b01111);           
  wire f9jz4kxv632mfmwjuwinhm = (xfkngdj3jaifg == 5'b10111);           
  wire qgge30ma6bacftkfuwr = (xfkngdj3jaifg == 5'b00000);           
  wire tv_mqy2vnetyki2mitz = (xfkngdj3jaifg == 5'b00001);
  wire iqlkuiiuioeb0zx_mespm = (xfkngdj3jaifg == 5'b00010);
  wire b2rqyt08n40btyec123 = (xfkngdj3jaifg == 5'b00011);
  wire nielo5a2gnsny_mbq2 = (xfkngdj3jaifg == 5'b00100);
  wire pnz7nx6huw6bc2xirgh = (xfkngdj3jaifg == 5'b00101);
  wire u1y9fqpjmgbvqp01zyup348 = (xfkngdj3jaifg == 5'b00110);
  wire mv0ortg5fw6xo5qko1gvm4 = (xfkngdj3jaifg == 5'b00111);



  wire qgai63fi1e6hqmwnsi7t = (xfkngdj3jaifg == 5'b11000);           
  wire yzqtbppdh3mlkyfzf0g6at = (xfkngdj3jaifg == 5'b11001);           
  wire nf2wc7g6poblu9r9_r = (xfkngdj3jaifg == 5'b11011);           

  wire auauwu7otyuaf2eindwrip = (xfkngdj3jaifg == 5'b10001);           
  wire jzb70ho_u3wii0cb_zw = (xfkngdj3jaifg == 5'b10000);           
  wire c6svrw070n8tv5npikqj18 = (xfkngdj3jaifg == 5'b10100);           
  wire pk4bj6ne4riq5l_gqv9maw_ = (xfkngdj3jaifg == 5'b10010);           





  wire osr23kerkrxjqbsvthv5n5 = (uk0ahn6nnbba7 == 7'b0111100);
  wire wambasxikyrgwdud7610fe = (uk0ahn6nnbba7 == 7'b0110100);


  wire g1qw0ijt6cz4o1fnmqoyhd = (uk0ahn6nnbba7 == 7'b0111101);
  wire bja_lg9vofv9y0s4oddhrjc = (uk0ahn6nnbba7 == 7'b0110101);
  wire flv_cd606fxf7i739917y8 = (uk0ahn6nnbba7 == 7'b0100100);
  wire rc04_8vnldazobtsw8nkr8 = (uk0ahn6nnbba7 == 7'b0100101);

  wire xxejssnpnxt8oi1caja = (uk0ahn6nnbba7 == 7'b0101110);
  wire rywrk93gumczcc8csvqrzq = (uk0ahn6nnbba7 == 7'b0111110);
  wire jysojps4nkgwbif943 = (uk0ahn6nnbba7 == 7'b0100110);
  wire rh5f36cuohtogtfizd = (uk0ahn6nnbba7 == 7'b0100111);
  wire n9p62t8e0cj6fl5zrn5 = (uk0ahn6nnbba7 == 7'b1100100);
  wire yurptvixnwx0aqsvdhdz = (uk0ahn6nnbba7 == 7'b1100110);
  wire of66mj2r_fom_q_y69j = (uk0ahn6nnbba7 == 7'b1100101);
  wire kwpxw02f_f6zyvb3it4sg4 = (uk0ahn6nnbba7 == 7'b0110110);

  wire as0og67e31vm7n6eodm = (uk0ahn6nnbba7 == 7'b1101110); 
  wire eong280dut8vgr73a14ab = (uk0ahn6nnbba7 == 7'b1110110);
  wire fn4lp09r_3zy48ytjb88 = (uk0ahn6nnbba7 == 7'b1101101);
  wire yukkytmyqpym19_1wwu_wg = (uk0ahn6nnbba7 == 7'b1110101);
  wire g4rhn7qi8xjp3mjyfl14ar3 = (uk0ahn6nnbba7 == 7'b1110100);
  wire d_7ca9przr4vewb9fcojf6l = (uk0ahn6nnbba7 == 7'b1101100);
  wire gr5b6bl6ypmzx3z57tmi = (uk0ahn6nnbba7 == 7'b0101111);
  wire vubg64i36fbtxkcl4s776lk = (uk0ahn6nnbba7 == 7'b1000100);
  wire gankodz2wzpdwh5hez = (uk0ahn6nnbba7 == 7'b1001100);
  wire opprr4u0rfe_9t1ilq = (uk0ahn6nnbba7 == 7'b0110111);
  wire ra742uamumnh7ulbty15 = (uk0ahn6nnbba7 == 7'b0101000);           



  wire xalf55zxhxx021sqlvd9_9 = (uk0ahn6nnbba7 == 7'b0101001);
  wire hfkmqai7ufo0_uc36i = (uk0ahn6nnbba7 == 7'b0111001);
  wire bwbrcnczkn_1flyk41tn5q8 = (uk0ahn6nnbba7 == 7'b0110001);

  wire mw5b0jbgrdfc4zozpy333k = (uk0ahn6nnbba7 == 7'b0101010);
  wire xvbpjhbrdw506s4r5je_v = (uk0ahn6nnbba7 == 7'b0100010);
  wire i_npu8b57pt8jq9y8wi6 = (uk0ahn6nnbba7 == 7'b0111010);
  wire ot56pcza1qpiqzjwuib4ioq = (uk0ahn6nnbba7 == 7'b0110010);

  wire umom31fkh4dmsle8dt = (uk0ahn6nnbba7 == 7'b0100011);
  wire ew4asffkh_z5lao1cnzk9g = (uk0ahn6nnbba7 == 7'b0101011);
  wire q4yuw6wl9o929gj8k2ovt = (uk0ahn6nnbba7 == 7'b0110011);
  wire zieb2_ok0e3farrv89q = (uk0ahn6nnbba7 == 7'b0111011);

  wire e9kyqn6z0nnxcqwggfu2c = (uk0ahn6nnbba7[6:1] == 6'b110101);       

  wire qr23_2sadkfk2963qo = (uk0ahn6nnbba7 == 7'b0111111);

  wire fr9vuzzy67toa8_rpz_ = (uk0ahn6nnbba7 == 7'b0011011);
  wire t33zd67g1c1fzxs_g27e34r = (uk0ahn6nnbba7 == 7'b1000110);           
  wire n0cr2bdx84qfgao3_gy8g9 = (uk0ahn6nnbba7 == 7'b1001110);
  wire crhfv2tcnpzr02ktjbc = (uk0ahn6nnbba7 == 7'b1000101);
  wire hmrtc229uz_sqjxkb8myxe = (uk0ahn6nnbba7 == 7'b1001101);
  wire pq_m0zj_hjvfii9out1 = (uk0ahn6nnbba7 == 7'b1000010);           
  wire brnnngwkv59w2kz9usv3k8 = (uk0ahn6nnbba7 == 7'b1110010);           
  wire sketktuyfh2vxjbshrr = (uk0ahn6nnbba7 == 7'b1111010);
  wire styktg7w7fi36jw0e5n4h93 = (uk0ahn6nnbba7 == 7'b1010110);           

  wire b12f43e4j_bhgigw_xvwmqe = (uk0ahn6nnbba7 == 7'b0001111);
  wire i_nd_auanr4nliiv9ru_mjy = (uk0ahn6nnbba7 == 7'b0010111);
  wire ha7x94wp2o8bpzvtiq_d = (uk0ahn6nnbba7 == 7'b0011111);
  wire tfcuen58mdto351cstsry5 = (uk0ahn6nnbba7 == 7'b1010111);           
  wire gp1add95ubo7akpuxefg1 = (uk0ahn6nnbba7 == 7'b1011111);
  wire wp2e1icm345eqoi7xse0mo = (uk0ahn6nnbba7 == 7'b1110011);           
  wire i37i_iou1kvjw2svv8 = (uk0ahn6nnbba7[6:1] == 6'b111010);       
  wire ny5cwervdr0wq805l6q = (uk0ahn6nnbba7 == 7'b1100111);           
  wire cbgxogbpgug3v8_faeo3 = (uk0ahn6nnbba7 == 7'b1101111);
  wire ij_r_y_kd47mgo6xio4viq = (uk0ahn6nnbba7 == 7'b1110111);
  wire lxbdxce1h6f_1nvn8vmkz = (uk0ahn6nnbba7 == 7'b1011110);
  wire w8iyjc4aw5thgv1c4vqr9vl = (uk0ahn6nnbba7[6:5] == 2'b11);           
  wire x99kg2smyvi6ahhq46x = (uk0ahn6nnbba7[1:0] == 2'b00);           


  
  
  
  

  
  
  
  wire pmmtjgnf20j2o_r     = t61y7hkwkrvm7s & c7npl5770szduubj6_grim & ezupw6o2yfm5ojugrc3;						
  wire wgjot58w1__ndyr81f    = t61y7hkwkrvm7s & whvtopzve8q_t001lyx & ezupw6o2yfm5ojugrc3;
  wire py50qt89qihhrq6frt60     = t61y7hkwkrvm7s & d9gmx9ccvp0rgcy7n_ii & ezupw6o2yfm5ojugrc3;						
  wire uxmg0dt8ik73agsf    = t61y7hkwkrvm7s & vrn4ssw1i97fztoyaq5kq & ezupw6o2yfm5ojugrc3;
  wire x9o36wx2sxi_96riv      = t61y7hkwkrvm7s & q8xucja6w9gzw4ujn6f7 & ezupw6o2yfm5ojugrc3;
  wire l2mrfrrlbbj8wb25j     = t61y7hkwkrvm7s & gv_izfe7yqh4gkvf76e93ct & ezupw6o2yfm5ojugrc3;
  wire sx2u7wkkrnzxotilhg      = t61y7hkwkrvm7s & wbsrjrrr8rt_27m9rwnm_ & ezupw6o2yfm5ojugrc3;
  wire jjudyrfeov9o45jiy     = t61y7hkwkrvm7s & l9_rbvynoe7x8o0_n_27icr & ezupw6o2yfm5ojugrc3;
  wire peoqulwt1lrkwd      = t61y7hkwkrvm7s & puc5pybv0exsbi1jenrc & ezupw6o2yfm5ojugrc3;
  wire tgghwgdy9ilyjs3vanp8     = t61y7hkwkrvm7s & uzvf9tjdfep6fv53xc6uakt & ezupw6o2yfm5ojugrc3;
  wire y5g_0z60_kaqxvn1       = t61y7hkwkrvm7s & iye23utobc0hah06xcesc14 & ezupw6o2yfm5ojugrc3;
  wire xdg0xfnp9f4p17fux      = t61y7hkwkrvm7s & tqsbmvgi1q8l40_d8_5 & ezupw6o2yfm5ojugrc3;
  wire stw6xp6m1y7hi5xy      = t61y7hkwkrvm7s & bepkj4gbb77isq3_v9 & d24iqtxvb2trplxk2m;
  wire sganc4k2sd9qhhyt     = t61y7hkwkrvm7s & ra742uamumnh7ulbty15 & d24iqtxvb2trplxk2m;
  wire m668z5d_2pgvlzqtt0r      = t61y7hkwkrvm7s & i3yg5uqgsrfhxxu1pt4o3 & d24iqtxvb2trplxk2m;
  wire f5obla9jfvqtwy50zglh     = t61y7hkwkrvm7s & po6ddes535c20_mmy_2u85p & d24iqtxvb2trplxk2m;
  wire yxhb2hnxchdqcag9u9      = t61y7hkwkrvm7s & uncepq376ovruspfffvl5 & d24iqtxvb2trplxk2m;
  wire af7cl38e7futiwz7m5     = t61y7hkwkrvm7s & xalf55zxhxx021sqlvd9_9 & d24iqtxvb2trplxk2m;
  wire xh3sniad_mq0m5j2ilk     = t61y7hkwkrvm7s & bwbrcnczkn_1flyk41tn5q8 & d24iqtxvb2trplxk2m;
  wire qcbi1__w_lbxar86    = t61y7hkwkrvm7s & hfkmqai7ufo0_uc36i & d24iqtxvb2trplxk2m;
  wire ngyb9j0p18mjlul4      = t61y7hkwkrvm7s & xvbpjhbrdw506s4r5je_v & d24iqtxvb2trplxk2m;
  wire zuhncrmyvsvqe31yah     = t61y7hkwkrvm7s & mw5b0jbgrdfc4zozpy333k & d24iqtxvb2trplxk2m;
  wire q7cxn6cfqixhf1j5c      = t61y7hkwkrvm7s & ot56pcza1qpiqzjwuib4ioq & d24iqtxvb2trplxk2m;
  wire as106js7z_6a17kl     = t61y7hkwkrvm7s & i_npu8b57pt8jq9y8wi6 & d24iqtxvb2trplxk2m;
  wire z1u9mb0is61kapi     = t61y7hkwkrvm7s & umom31fkh4dmsle8dt & d24iqtxvb2trplxk2m;
  wire hjj29yefty1oa5g1    = t61y7hkwkrvm7s & ew4asffkh_z5lao1cnzk9g & d24iqtxvb2trplxk2m;
  wire dgoqvucxrbc7u23zbh1     = t61y7hkwkrvm7s & q4yuw6wl9o929gj8k2ovt & d24iqtxvb2trplxk2m;
  wire k7u3ztuoje2dfwlb    = t61y7hkwkrvm7s & zieb2_ok0e3farrv89q & d24iqtxvb2trplxk2m;
  wire no41cqtslidyozjc3b4     = t61y7hkwkrvm7s & iye23utobc0hah06xcesc14 & d24iqtxvb2trplxk2m;
  wire yo4avylbzg3xikezi    = t61y7hkwkrvm7s & tqsbmvgi1q8l40_d8_5 & d24iqtxvb2trplxk2m;
  wire ytpvnxr5ldhrfhe     = t61y7hkwkrvm7s & tfcuen58mdto351cstsry5 & d24iqtxvb2trplxk2m;
  wire wyzwj_3yh41jvmcgv    = t61y7hkwkrvm7s & gp1add95ubo7akpuxefg1 & d24iqtxvb2trplxk2m;
  wire fgg6hxc67s_zufvn    = t61y7hkwkrvm7s & ny5cwervdr0wq805l6q & d24iqtxvb2trplxk2m;
  wire bx8ta8ntqmkd296igjj5cm   = t61y7hkwkrvm7s & cbgxogbpgug3v8_faeo3 & d24iqtxvb2trplxk2m;
  wire x7i6k3jtvgugfgwm    = t61y7hkwkrvm7s & ij_r_y_kd47mgo6xio4viq & d24iqtxvb2trplxk2m;
  wire cmayk4nyxf2fgdyrgbdm   = t61y7hkwkrvm7s & yf083xcjpnohrzqky4 & d24iqtxvb2trplxk2m;
  wire mtjkl28_lqkguy1g96p4     = t61y7hkwkrvm7s & styktg7w7fi36jw0e5n4h93 & d24iqtxvb2trplxk2m;
  wire d_rtbt5u2waj29pq38aw    = t61y7hkwkrvm7s & lxbdxce1h6f_1nvn8vmkz & d24iqtxvb2trplxk2m;
  wire n61z5eg85z3qt6ym     = t61y7hkwkrvm7s & mso_1l7nnv4ac14pv6qh & d24iqtxvb2trplxk2m;
  wire tpxnwqn02te7dxkfod1c     = t61y7hkwkrvm7s & duf6qt_vm6jkmkv9xu9 & d24iqtxvb2trplxk2m;
  wire zociru6_rc45yinp5k     = t61y7hkwkrvm7s & f6kcevztmpqpnc8xp3_r4 & d24iqtxvb2trplxk2m;
  wire pp7lw68tzorrt1ry       = t61y7hkwkrvm7s & m33lelq8_5u26vfl7hl6z & d24iqtxvb2trplxk2m;
  wire qwszvnfbt4kifn      = t61y7hkwkrvm7s & amf97jdmi0f4r4z2kmw & d24iqtxvb2trplxk2m;
  wire l8skguypzoiw9k       = t61y7hkwkrvm7s & gu_2fhfulrttqq4e_fiax & d24iqtxvb2trplxk2m;
  wire bqonmn9o0yi3pta98ja      = t61y7hkwkrvm7s & wambasxikyrgwdud7610fe & d24iqtxvb2trplxk2m;
  wire zse6ubdm7b85h4fv      = t61y7hkwkrvm7s & osr23kerkrxjqbsvthv5n5 & d24iqtxvb2trplxk2m;
  wire w6ojhbqk3lmsoe464      = t61y7hkwkrvm7s & k3sfqtpqynzqda4xtugl4 & d24iqtxvb2trplxk2m;
  wire l47a5b8y1b7jw87t      = t61y7hkwkrvm7s & bja_lg9vofv9y0s4oddhrjc & d24iqtxvb2trplxk2m;
  wire f3zsw2wieuvu92v24b      = t61y7hkwkrvm7s & g1qw0ijt6cz4o1fnmqoyhd & d24iqtxvb2trplxk2m;
  wire ata32ab_8ia7entoq1d      = t61y7hkwkrvm7s & flv_cd606fxf7i739917y8 & d24iqtxvb2trplxk2m;
  wire wxfxhstnh27mwfsba43x     = t61y7hkwkrvm7s & rc04_8vnldazobtsw8nkr8 & d24iqtxvb2trplxk2m;
  wire g1bqvr3iwplkb20wpvq      = t61y7hkwkrvm7s & xxejssnpnxt8oi1caja & d24iqtxvb2trplxk2m;
  wire cflo9l4odlq3l0so     = t61y7hkwkrvm7s & kwpxw02f_f6zyvb3it4sg4 & d24iqtxvb2trplxk2m;
  wire aw1b57cswb2mmub     = t61y7hkwkrvm7s & rywrk93gumczcc8csvqrzq & d24iqtxvb2trplxk2m;
  wire jv62xshm61xc3633g      = t61y7hkwkrvm7s & jysojps4nkgwbif943 & d24iqtxvb2trplxk2m;
  wire casdl4x6djchiuqej     = t61y7hkwkrvm7s & rh5f36cuohtogtfizd & d24iqtxvb2trplxk2m;
  wire os5cdj3yxqxq58sz      = t61y7hkwkrvm7s & n9p62t8e0cj6fl5zrn5 & ezupw6o2yfm5ojugrc3;
  wire neja7y5h1cux76u7ru      = t61y7hkwkrvm7s & yurptvixnwx0aqsvdhdz & ezupw6o2yfm5ojugrc3;
  wire uxstixgq52wcp394s2bq    = t61y7hkwkrvm7s & of66mj2r_fom_q_y69j & ezupw6o2yfm5ojugrc3;
  wire g_k_2hcsq4fllbhbyvp      = t61y7hkwkrvm7s & fcpfa9hp28k7bapl82 & d24iqtxvb2trplxk2m;
  wire fy_5mx58b8k0rbva      = t61y7hkwkrvm7s & hx3wrp4j8s1ov27syy & d24iqtxvb2trplxk2m;
  wire mbbkhwc6igem3g      = t61y7hkwkrvm7s & naged_b50dbpmu745zp & d24iqtxvb2trplxk2m;
  wire w8kkipg2caprcl38r      = t61y7hkwkrvm7s & xfrai8f3331hb4z5ww5_ & d24iqtxvb2trplxk2m;
  wire b4z_up9nkirbcj3jl      = t61y7hkwkrvm7s & cvhx1ne2we07dkbzbpwakl & d24iqtxvb2trplxk2m;
  wire xpa9jhun_nud6epww      = t61y7hkwkrvm7s & toaowsb_5w3arwmyl2 & d24iqtxvb2trplxk2m;
  wire sv78kz_4osrj8ymh53m     = t61y7hkwkrvm7s & mnd8c7lvcdtsypyiygspg & d24iqtxvb2trplxk2m;
  wire zdwvt5v7m2azz1zncqlz     = t61y7hkwkrvm7s & eu9j7rkhrocfjsewdf6mfvu & d24iqtxvb2trplxk2m;
  wire l_5fge2sjzcghz15     = t61y7hkwkrvm7s & rf284mrjg_bqa1hj60swyf & d24iqtxvb2trplxk2m;
  wire ikrh3ggnb20z70nz    = t61y7hkwkrvm7s & rgjf1vrs4iai2hif_09x & d24iqtxvb2trplxk2m;
  wire gh34i2cii_rlj2      = t61y7hkwkrvm7s & ng7__qxmefe1xunqibay7zg & ezupw6o2yfm5ojugrc3;
  wire jhx20z5y9lr18q       = t61y7hkwkrvm7s & rf284mrjg_bqa1hj60swyf & ezupw6o2yfm5ojugrc3;
  wire obzhb904qzxr8b3       = t61y7hkwkrvm7s & v3hylq_n52mziras6qen & ezupw6o2yfm5ojugrc3;
  wire drexvwdx10vfyckm2w    = t61y7hkwkrvm7s & qcpti7i25_4w_aexyk1 & d24iqtxvb2trplxk2m;
  wire emfepzk_i3iart3w     = t61y7hkwkrvm7s & v3hylq_n52mziras6qen & d24iqtxvb2trplxk2m;
  wire bpctswvy4clemt9h    = t61y7hkwkrvm7s & k_h8qestuhin60n5ckxmkfx & d24iqtxvb2trplxk2m;
  wire w9tkyl3th_cayu_wvi      = t61y7hkwkrvm7s & ei5le5r3u2ub_qlszr3u6lq & ezupw6o2yfm5ojugrc3;
  wire gkfxs8wvvzhw35g2w       = t61y7hkwkrvm7s & gr5b6bl6ypmzx3z57tmi & d24iqtxvb2trplxk2m;
  wire qo4hl0cqzct4xyimucu     = t61y7hkwkrvm7s & vubg64i36fbtxkcl4s776lk & d24iqtxvb2trplxk2m;
  wire jqc0fopjngrnmrha1ca9     = t61y7hkwkrvm7s & gankodz2wzpdwh5hez & d24iqtxvb2trplxk2m;
  wire nris9imni2zozl_9adll     = t61y7hkwkrvm7s & wbsrjrrr8rt_27m9rwnm_ & d24iqtxvb2trplxk2m;
  wire gp2roes6p_wvpktfh     = t61y7hkwkrvm7s & t33zd67g1c1fzxs_g27e34r & d24iqtxvb2trplxk2m;
  wire rhpud0ssrcsrol8rx8nu4    = t61y7hkwkrvm7s & n0cr2bdx84qfgao3_gy8g9 & d24iqtxvb2trplxk2m;
  wire p57xv2ht1u5oz2jyd9m     = t61y7hkwkrvm7s & crhfv2tcnpzr02ktjbc & d24iqtxvb2trplxk2m;
  wire yikkze0bi4xdf5kgp    = t61y7hkwkrvm7s & hmrtc229uz_sqjxkb8myxe & d24iqtxvb2trplxk2m;
  wire ewo2z4ywjzk3rqw0c9di    = t61y7hkwkrvm7s & l9_rbvynoe7x8o0_n_27icr & d24iqtxvb2trplxk2m;
  wire g9bfl499lfhirrrjln     = t61y7hkwkrvm7s & pq_m0zj_hjvfii9out1 & d24iqtxvb2trplxk2m;
  wire g2esflomposu_jm     = t61y7hkwkrvm7s & q8xucja6w9gzw4ujn6f7 & d24iqtxvb2trplxk2m;
  wire d1knhe17l7248qdlx3d    = t61y7hkwkrvm7s & zpue29q3_sghsyln86mp & d24iqtxvb2trplxk2m;
  wire tdtkoiumk_q1_zlrgx1n_    = t61y7hkwkrvm7s & ef0qt3ctq84209xo8ti63mv & d24iqtxvb2trplxk2m;
  wire nn04ut84g694dyj3ngt     = t61y7hkwkrvm7s & gv_izfe7yqh4gkvf76e93ct & d24iqtxvb2trplxk2m;
  wire fx8tfw6ht51x591xovf     = t61y7hkwkrvm7s & hobxt8_ayp1au2dt6zmqdcc & d24iqtxvb2trplxk2m;
  wire m06_keb0crbj3pkd_     = t61y7hkwkrvm7s & bju5h0qfjwac44bgx65qbdh & d24iqtxvb2trplxk2m;
  wire yo0gy1w6lzj_sxzxb0a     = t61y7hkwkrvm7s & hhf4if064tv59lxifk & d24iqtxvb2trplxk2m;
  wire aquf29t5dbq4elt      = t61y7hkwkrvm7s & o5frxem9qrhhps9sw7n & ezupw6o2yfm5ojugrc3;
  wire eaqgia_mu1yu9vo2nszk     = t61y7hkwkrvm7s & yf083xcjpnohrzqky4 & ezupw6o2yfm5ojugrc3;

  wire i92ohq_11aclejsw9    = t61y7hkwkrvm7s & as0og67e31vm7n6eodm & d24iqtxvb2trplxk2m; 
  wire lihv1jjl5cbn0k8m1    = t61y7hkwkrvm7s & eong280dut8vgr73a14ab & d24iqtxvb2trplxk2m; 
  wire ogxv3q5tyb1genv51czg    = t61y7hkwkrvm7s & o5frxem9qrhhps9sw7n & d24iqtxvb2trplxk2m; 
  wire d_t7c_en995wivae5jc6g    = t61y7hkwkrvm7s & fn4lp09r_3zy48ytjb88 & d24iqtxvb2trplxk2m; 
  wire r0oo_zmre7ja5s9h    = t61y7hkwkrvm7s & yukkytmyqpym19_1wwu_wg & d24iqtxvb2trplxk2m; 
  wire o63p86lpcfcy7xuj55    = t61y7hkwkrvm7s & ng7__qxmefe1xunqibay7zg & d24iqtxvb2trplxk2m; 
  wire x43fhodherbcf_w4w   = t61y7hkwkrvm7s & d_7ca9przr4vewb9fcojf6l & d24iqtxvb2trplxk2m; 
  wire hc6mrm8abcf82sqypnsn   = t61y7hkwkrvm7s & g4rhn7qi8xjp3mjyfl14ar3 & d24iqtxvb2trplxk2m; 
  wire tsfbnnx02_rdxvvpvk5a   = t61y7hkwkrvm7s & ei5le5r3u2ub_qlszr3u6lq & d24iqtxvb2trplxk2m; 

  wire htdih4lhmspfu8_     = bpctswvy4clemt9h;
  wire dserv0gb0p2c2yof     = t61y7hkwkrvm7s & duf6qt_vm6jkmkv9xu9 & t8jc64yc1l6q8eclq_c; 
  wire g2625iw5_kvvco4hf     = t61y7hkwkrvm7s & f6kcevztmpqpnc8xp3_r4 & t8jc64yc1l6q8eclq_c; 

  wire nhxdacdf6m8xlgp0gi    = t61y7hkwkrvm7s & k3sfqtpqynzqda4xtugl4 & t8jc64yc1l6q8eclq_c; 
  wire xdtf0ycp133xtiom9    = t61y7hkwkrvm7s & bja_lg9vofv9y0s4oddhrjc & t8jc64yc1l6q8eclq_c; 
  wire fimif9coi4wgjje86n652    = t61y7hkwkrvm7s & g1qw0ijt6cz4o1fnmqoyhd & t8jc64yc1l6q8eclq_c; 

  wire g690wip_77275ygun     = t61y7hkwkrvm7s & m33lelq8_5u26vfl7hl6z & t8jc64yc1l6q8eclq_c; 
  wire eo1ocops3gp9phz4jc3    = t61y7hkwkrvm7s & amf97jdmi0f4r4z2kmw & t8jc64yc1l6q8eclq_c; 
  wire akky00pxrb96le0sige5g    = fx8tfw6ht51x591xovf;
  wire s94qy2bqkpnqqumbxck   = t61y7hkwkrvm7s & rc04_8vnldazobtsw8nkr8 & t8jc64yc1l6q8eclq_c; 
  wire ds6le0delcgakxcymi    = t61y7hkwkrvm7s & xxejssnpnxt8oi1caja & t8jc64yc1l6q8eclq_c; 
  wire kjwyayvk_cqc5s0li40i   = t61y7hkwkrvm7s & kwpxw02f_f6zyvb3it4sg4 & t8jc64yc1l6q8eclq_c; 
  wire l45fdj1kcz0x06i9k   = t61y7hkwkrvm7s & rywrk93gumczcc8csvqrzq & t8jc64yc1l6q8eclq_c; 
  wire e65i99f2zhb74wze9lg    = t61y7hkwkrvm7s & jysojps4nkgwbif943 & t8jc64yc1l6q8eclq_c; 
  wire sqy4k5rpyr8won7x_a3h   = t61y7hkwkrvm7s & rh5f36cuohtogtfizd & t8jc64yc1l6q8eclq_c; 
  wire dogjt36yta_opjg     = t61y7hkwkrvm7s & gu_2fhfulrttqq4e_fiax & t8jc64yc1l6q8eclq_c; 
  wire k8wg766owq6fcetyyuo    = t61y7hkwkrvm7s & wambasxikyrgwdud7610fe & t8jc64yc1l6q8eclq_c; 
  wire m5fgnytsm5kbh2sbrzf    = t61y7hkwkrvm7s & osr23kerkrxjqbsvthv5n5 & t8jc64yc1l6q8eclq_c; 

  wire a24tfk9zcc_2qh6mtd_1dsw = 
                                 y5g_0z60_kaqxvn1
                               | xdg0xfnp9f4p17fux
                               | sx2u7wkkrnzxotilhg
                               | jjudyrfeov9o45jiy
                               | peoqulwt1lrkwd
                               | tgghwgdy9ilyjs3vanp8
                               | x9o36wx2sxi_96riv
                               | l2mrfrrlbbj8wb25j
                               | pmmtjgnf20j2o_r
                               | wgjot58w1__ndyr81f
                               | py50qt89qihhrq6frt60
                               | uxmg0dt8ik73agsf
                               ;

  wire niiot38ff0zsxxncd0u_5fljm__dl  = 
                              | g_k_2hcsq4fllbhbyvp
                              | fy_5mx58b8k0rbva
                              | mbbkhwc6igem3g
                              | w8kkipg2caprcl38r
                              | b4z_up9nkirbcj3jl
                              | xpa9jhun_nud6epww
                              ;
  wire bsjfhtce07tsob5_b486_ou_y_h6cae = 
                                ngyb9j0p18mjlul4
                              | q7cxn6cfqixhf1j5c
                              | n61z5eg85z3qt6ym
                              | tpxnwqn02te7dxkfod1c
                              | zociru6_rc45yinp5k
                              | no41cqtslidyozjc3b4
                              | ytpvnxr5ldhrfhe
                              | xh3sniad_mq0m5j2ilk
                              | stw6xp6m1y7hi5xy
                              | emfepzk_i3iart3w
                              | bpctswvy4clemt9h
                              | i92ohq_11aclejsw9
                              | lihv1jjl5cbn0k8m1
                              | ogxv3q5tyb1genv51czg
                              | d_t7c_en995wivae5jc6g
                              | r0oo_zmre7ja5s9h
                              | o63p86lpcfcy7xuj55
                              | htdih4lhmspfu8_
                              | dserv0gb0p2c2yof
                              | g2625iw5_kvvco4hf
                              ;

  wire hxv8akm9tnbagx = a24tfk9zcc_2qh6mtd_1dsw | niiot38ff0zsxxncd0u_5fljm__dl;

  wire ucwkku1t4g36u3iukgb = 
                      x9o36wx2sxi_96riv  | l2mrfrrlbbj8wb25j | pmmtjgnf20j2o_r | wgjot58w1__ndyr81f | py50qt89qihhrq6frt60 | uxmg0dt8ik73agsf
                    | pp7lw68tzorrt1ry | qwszvnfbt4kifn | l8skguypzoiw9k | bqonmn9o0yi3pta98ja | zse6ubdm7b85h4fv | ata32ab_8ia7entoq1d | wxfxhstnh27mwfsba43x
                    | g1bqvr3iwplkb20wpvq | cflo9l4odlq3l0so | aw1b57cswb2mmub | jv62xshm61xc3633g | casdl4x6djchiuqej | mtjkl28_lqkguy1g96p4
                    | d_rtbt5u2waj29pq38aw | gp2roes6p_wvpktfh | rhpud0ssrcsrol8rx8nu4 | p57xv2ht1u5oz2jyd9m | yikkze0bi4xdf5kgp | ewo2z4ywjzk3rqw0c9di
                    ;

  wire avjo592wbov8cr5i = y5g_0z60_kaqxvn1  | xdg0xfnp9f4p17fux | sx2u7wkkrnzxotilhg | jjudyrfeov9o45jiy | peoqulwt1lrkwd
                      | tgghwgdy9ilyjs3vanp8 | os5cdj3yxqxq58sz | neja7y5h1cux76u7ru | uxstixgq52wcp394s2bq
                      ;
  wire kp1fyknoq74q3vs   = avjo592wbov8cr5i | ucwkku1t4g36u3iukgb;

  wire yunpydbojvbs7t1vv3n9ir = y5g_0z60_kaqxvn1 | xdg0xfnp9f4p17fux 
                        ;
  wire rh93dqz7x7e76_rwvdq_gv = yunpydbojvbs7t1vv3n9ir;
  wire wewa0sb6nm_e_8n25xoi = g_k_2hcsq4fllbhbyvp |fy_5mx58b8k0rbva |mbbkhwc6igem3g |x9o36wx2sxi_96riv |l2mrfrrlbbj8wb25j 
                          ;
  wire dwf3ct8epliykbwg6fpvn1d = wewa0sb6nm_e_8n25xoi; 

  wire f_l92j9mkhdmknnhn2 = w8kkipg2caprcl38r |b4z_up9nkirbcj3jl |xpa9jhun_nud6epww 
                          
                          | d_t7c_en995wivae5jc6g | r0oo_zmre7ja5s9h | o63p86lpcfcy7xuj55
                          
                          ; 
  wire syyd9204a47y6qq9cyxvn7s = 
                            d_t7c_en995wivae5jc6g | r0oo_zmre7ja5s9h | o63p86lpcfcy7xuj55
                          
                          ;
  wire woiza4felzgpik5ue3hx8 = yunpydbojvbs7t1vv3n9ir | wewa0sb6nm_e_8n25xoi | f_l92j9mkhdmknnhn2; 
  wire x4zc788yz37xi4o6fcfpux = rh93dqz7x7e76_rwvdq_gv | dwf3ct8epliykbwg6fpvn1d | syyd9204a47y6qq9cyxvn7s; 
 
 
 
 
 

  wire n4dlb4x1wzqqyr98jl7v8t_apmfb = xdg0xfnp9f4p17fux | jjudyrfeov9o45jiy | tgghwgdy9ilyjs3vanp8 | l2mrfrrlbbj8wb25j | wgjot58w1__ndyr81f | uxmg0dt8ik73agsf
                                | tpxnwqn02te7dxkfod1c | qwszvnfbt4kifn | zse6ubdm7b85h4fv | wxfxhstnh27mwfsba43x | aw1b57cswb2mmub | casdl4x6djchiuqej
                                | d_rtbt5u2waj29pq38aw | rhpud0ssrcsrol8rx8nu4 | ewo2z4ywjzk3rqw0c9di
                                
                                
                                
                                ;


  wire pm3poaltg6mtmffm_87yhorfj9eort_ = qo4hl0cqzct4xyimucu
                               | jqc0fopjngrnmrha1ca9
                               | nris9imni2zozl_9adll
                               | w6ojhbqk3lmsoe464
                               | l47a5b8y1b7jw87t
                               | f3zsw2wieuvu92v24b
                               | sv78kz_4osrj8ymh53m
                               | zdwvt5v7m2azz1zncqlz
                               | l_5fge2sjzcghz15
                               | gkfxs8wvvzhw35g2w
                               | sganc4k2sd9qhhyt
                               | qcbi1__w_lbxar86
                               | wyzwj_3yh41jvmcgv
                               | yo4avylbzg3xikezi
                               | as106js7z_6a17kl
                               | zuhncrmyvsvqe31yah
                               | ikrh3ggnb20z70nz
                               | drexvwdx10vfyckm2w
                               | hjj29yefty1oa5g1
                               | dgoqvucxrbc7u23zbh1
                               | k7u3ztuoje2dfwlb
                               | fgg6hxc67s_zufvn
                               | bx8ta8ntqmkd296igjj5cm
                               | x7i6k3jtvgugfgwm
                               | cmayk4nyxf2fgdyrgbdm
                               | z1u9mb0is61kapi
                               | m668z5d_2pgvlzqtt0r
                               | f5obla9jfvqtwy50zglh
                               | yxhb2hnxchdqcag9u9
                               | af7cl38e7futiwz7m5
                               | g9bfl499lfhirrrjln
                               | g2esflomposu_jm
                               | nn04ut84g694dyj3ngt
                               | fx8tfw6ht51x591xovf
                               | d1knhe17l7248qdlx3d
                               | tdtkoiumk_q1_zlrgx1n_
                               | m06_keb0crbj3pkd_
                               | yo0gy1w6lzj_sxzxb0a
                               | bsjfhtce07tsob5_b486_ou_y_h6cae
                               | nhxdacdf6m8xlgp0gi
                               | xdtf0ycp133xtiom9
                               | fimif9coi4wgjje86n652
                               | akky00pxrb96le0sige5g
                               | s94qy2bqkpnqqumbxck
                               | g690wip_77275ygun
                               | eo1ocops3gp9phz4jc3
                               | ds6le0delcgakxcymi
                               | kjwyayvk_cqc5s0li40i
                               | l45fdj1kcz0x06i9k
                               | e65i99f2zhb74wze9lg
                               | sqy4k5rpyr8won7x_a3h
                               | dogjt36yta_opjg
                               | k8wg766owq6fcetyyuo
                               | m5fgnytsm5kbh2sbrzf
                               | x43fhodherbcf_w4w
                               | hc6mrm8abcf82sqypnsn
                               | tsfbnnx02_rdxvvpvk5a
                               ;

  wire hf3_u19xhtm47jygm346ih5592f =  niiot38ff0zsxxncd0u_5fljm__dl | pm3poaltg6mtmffm_87yhorfj9eort_;                               

  wire upbbycb5makv3xss7d_ueoxns88bj;


  wire ccb88tt72pm4kk3aiztl_ = 
                             gkfxs8wvvzhw35g2w
                           | sganc4k2sd9qhhyt
                           | qcbi1__w_lbxar86
                           | wyzwj_3yh41jvmcgv
                           | yo4avylbzg3xikezi
                           | as106js7z_6a17kl
                           | zuhncrmyvsvqe31yah
                           | pp7lw68tzorrt1ry
                           | qwszvnfbt4kifn
                           | l8skguypzoiw9k
                           | bqonmn9o0yi3pta98ja
                           | zse6ubdm7b85h4fv
                           | g690wip_77275ygun
                           | eo1ocops3gp9phz4jc3
                           | dogjt36yta_opjg
                           | k8wg766owq6fcetyyuo
                           | m5fgnytsm5kbh2sbrzf
                           | bsjfhtce07tsob5_b486_ou_y_h6cae
                           ;

  wire y1fgyae1uzj7ujuxqi3znyfnbb19hjsl = ngyb9j0p18mjlul4 | q7cxn6cfqixhf1j5c | no41cqtslidyozjc3b4 | ytpvnxr5ldhrfhe | xh3sniad_mq0m5j2ilk | stw6xp6m1y7hi5xy
                            | sganc4k2sd9qhhyt | qcbi1__w_lbxar86 | wyzwj_3yh41jvmcgv | yo4avylbzg3xikezi
                            | as106js7z_6a17kl | zuhncrmyvsvqe31yah | ikrh3ggnb20z70nz | drexvwdx10vfyckm2w | hjj29yefty1oa5g1 | dgoqvucxrbc7u23zbh1
                            | k7u3ztuoje2dfwlb | fgg6hxc67s_zufvn | bx8ta8ntqmkd296igjj5cm | x7i6k3jtvgugfgwm | cmayk4nyxf2fgdyrgbdm | z1u9mb0is61kapi
                            | m668z5d_2pgvlzqtt0r | f5obla9jfvqtwy50zglh | yxhb2hnxchdqcag9u9 | af7cl38e7futiwz7m5 | g9bfl499lfhirrrjln | g2esflomposu_jm
                            | nn04ut84g694dyj3ngt | fx8tfw6ht51x591xovf | d1knhe17l7248qdlx3d | tdtkoiumk_q1_zlrgx1n_ | m06_keb0crbj3pkd_ | yo0gy1w6lzj_sxzxb0a
                            | emfepzk_i3iart3w | bpctswvy4clemt9h
                            | htdih4lhmspfu8_ | nhxdacdf6m8xlgp0gi | g690wip_77275ygun | akky00pxrb96le0sige5g | ds6le0delcgakxcymi | kjwyayvk_cqc5s0li40i | e65i99f2zhb74wze9lg
                            | dogjt36yta_opjg | k8wg766owq6fcetyyuo 
                            ;

  wire sfwi4o77fiwv1s1kb4mmixcewjetb_1 = n61z5eg85z3qt6ym | tpxnwqn02te7dxkfod1c | fy_5mx58b8k0rbva | g_k_2hcsq4fllbhbyvp | qo4hl0cqzct4xyimucu | jqc0fopjngrnmrha1ca9
                                    | w6ojhbqk3lmsoe464 | l47a5b8y1b7jw87t | sv78kz_4osrj8ymh53m | zdwvt5v7m2azz1zncqlz | w8kkipg2caprcl38r  | b4z_up9nkirbcj3jl
                                    | d_t7c_en995wivae5jc6g | r0oo_zmre7ja5s9h
                                    | i92ohq_11aclejsw9 | lihv1jjl5cbn0k8m1
                                    | x43fhodherbcf_w4w | hc6mrm8abcf82sqypnsn
                                    ;

  wire oboq9ew68wxfv1zbbzbw6ovxumvp4ms = zociru6_rc45yinp5k | mbbkhwc6igem3g | xpa9jhun_nud6epww | nris9imni2zozl_9adll | f3zsw2wieuvu92v24b | l_5fge2sjzcghz15
                                       | ogxv3q5tyb1genv51czg |  o63p86lpcfcy7xuj55 | tsfbnnx02_rdxvvpvk5a
                                       ;

  wire ozipqe_4brzi2opcs5pi232jtqiu7_m6kuv = gkfxs8wvvzhw35g2w; 
  wire imwjfayr9ztr86owxp26dtq0onjtd6dp = eo1ocops3gp9phz4jc3 | s94qy2bqkpnqqumbxck | l45fdj1kcz0x06i9k | sqy4k5rpyr8won7x_a3h | m5fgnytsm5kbh2sbrzf; 

  wire n38usa0n35mgmntamkuxh2l5pd2gcwghz = xh3sniad_mq0m5j2ilk | stw6xp6m1y7hi5xy | sganc4k2sd9qhhyt | qcbi1__w_lbxar86
                                     | ikrh3ggnb20z70nz | drexvwdx10vfyckm2w | m668z5d_2pgvlzqtt0r | f5obla9jfvqtwy50zglh | yxhb2hnxchdqcag9u9 | af7cl38e7futiwz7m5   
                                     | g9bfl499lfhirrrjln | g2esflomposu_jm | nn04ut84g694dyj3ngt | fx8tfw6ht51x591xovf
                                     | emfepzk_i3iart3w | bpctswvy4clemt9h | d1knhe17l7248qdlx3d | tdtkoiumk_q1_zlrgx1n_ | m06_keb0crbj3pkd_ | yo0gy1w6lzj_sxzxb0a
                                     | htdih4lhmspfu8_ | nhxdacdf6m8xlgp0gi | g690wip_77275ygun | eo1ocops3gp9phz4jc3 | akky00pxrb96le0sige5g | s94qy2bqkpnqqumbxck
                                     | ds6le0delcgakxcymi | kjwyayvk_cqc5s0li40i | l45fdj1kcz0x06i9k | e65i99f2zhb74wze9lg | sqy4k5rpyr8won7x_a3h
                                     | dogjt36yta_opjg | k8wg766owq6fcetyyuo  | m5fgnytsm5kbh2sbrzf
                                     ;

  wire gm3156cuu5w0z0iabqd970k351i652n1u =  n61z5eg85z3qt6ym | g_k_2hcsq4fllbhbyvp | w8kkipg2caprcl38r | qo4hl0cqzct4xyimucu | w6ojhbqk3lmsoe464 
                                        | ngyb9j0p18mjlul4  | no41cqtslidyozjc3b4| yo4avylbzg3xikezi | zuhncrmyvsvqe31yah | z1u9mb0is61kapi| hjj29yefty1oa5g1 
                                        | fgg6hxc67s_zufvn | bx8ta8ntqmkd296igjj5cm
                                         | i92ohq_11aclejsw9
                                        ;

  wire n93vkxau7xxglljhnhsxg_4jddx13kcy =  tpxnwqn02te7dxkfod1c | fy_5mx58b8k0rbva | b4z_up9nkirbcj3jl | jqc0fopjngrnmrha1ca9 | l47a5b8y1b7jw87t
                                        | zociru6_rc45yinp5k | mbbkhwc6igem3g | xpa9jhun_nud6epww | nris9imni2zozl_9adll | f3zsw2wieuvu92v24b 
                                        | q7cxn6cfqixhf1j5c  | ytpvnxr5ldhrfhe| wyzwj_3yh41jvmcgv | as106js7z_6a17kl | dgoqvucxrbc7u23zbh1| k7u3ztuoje2dfwlb 
                                        | x7i6k3jtvgugfgwm | cmayk4nyxf2fgdyrgbdm | gkfxs8wvvzhw35g2w
                                        | lihv1jjl5cbn0k8m1 | ogxv3q5tyb1genv51czg
                                        ;
  wire t88i3logg39o9_7fi_4qgfve8slrofj4j = sv78kz_4osrj8ymh53m
                                        | d_t7c_en995wivae5jc6g | x43fhodherbcf_w4w
                                        ;
  wire e7ilxivhp9g8urh1klgvakcpqfmwjd5tw = zdwvt5v7m2azz1zncqlz  | l_5fge2sjzcghz15
                                       | r0oo_zmre7ja5s9h  | o63p86lpcfcy7xuj55
                                       | hc6mrm8abcf82sqypnsn  | tsfbnnx02_rdxvvpvk5a
                                       ;
  wire hhf5vk7i4v5m5s0diu0q2m6pmxzvm7zeyiv7r = ngyb9j0p18mjlul4 | q7cxn6cfqixhf1j5c | no41cqtslidyozjc3b4 | ytpvnxr5ldhrfhe | xh3sniad_mq0m5j2ilk | stw6xp6m1y7hi5xy
                            | sganc4k2sd9qhhyt | qcbi1__w_lbxar86 | wyzwj_3yh41jvmcgv | yo4avylbzg3xikezi
                            | as106js7z_6a17kl | zuhncrmyvsvqe31yah | hjj29yefty1oa5g1 | dgoqvucxrbc7u23zbh1
                            | k7u3ztuoje2dfwlb | fgg6hxc67s_zufvn | bx8ta8ntqmkd296igjj5cm | x7i6k3jtvgugfgwm | cmayk4nyxf2fgdyrgbdm | z1u9mb0is61kapi
                            | m668z5d_2pgvlzqtt0r | f5obla9jfvqtwy50zglh | yxhb2hnxchdqcag9u9 | af7cl38e7futiwz7m5 | g9bfl499lfhirrrjln | g2esflomposu_jm
                            | nn04ut84g694dyj3ngt | fx8tfw6ht51x591xovf | d1knhe17l7248qdlx3d | tdtkoiumk_q1_zlrgx1n_ | m06_keb0crbj3pkd_ | yo0gy1w6lzj_sxzxb0a
                            | g2625iw5_kvvco4hf | fimif9coi4wgjje86n652
                            | g690wip_77275ygun | akky00pxrb96le0sige5g | ds6le0delcgakxcymi | kjwyayvk_cqc5s0li40i | e65i99f2zhb74wze9lg
                            | dogjt36yta_opjg | k8wg766owq6fcetyyuo 
                            ;
  wire e9gctcgx_15frdmbcrevvtf_2lldmasrmr9gp = n61z5eg85z3qt6ym | tpxnwqn02te7dxkfod1c 
                                    | w6ojhbqk3lmsoe464 | l47a5b8y1b7jw87t  
                                    | d_t7c_en995wivae5jc6g | r0oo_zmre7ja5s9h
                                    | i92ohq_11aclejsw9 | lihv1jjl5cbn0k8m1
                                    | x43fhodherbcf_w4w | hc6mrm8abcf82sqypnsn 
                                    | qo4hl0cqzct4xyimucu | jqc0fopjngrnmrha1ca9
                                    ;

  wire wj4suc8dinc_9d5409y_to9toxtea5b3afqoc = zociru6_rc45yinp5k | f3zsw2wieuvu92v24b | l_5fge2sjzcghz15 
                                          | o63p86lpcfcy7xuj55 | tsfbnnx02_rdxvvpvk5a  | ogxv3q5tyb1genv51czg | nris9imni2zozl_9adll;

  wire o44zcer7fjl2e666o3w3zxacak78idnwavnn = gkfxs8wvvzhw35g2w; 

  wire iue4b0u82l97gr25u35a4wkzrr64s8kyxgwm = dserv0gb0p2c2yof | xdtf0ycp133xtiom9 |  eo1ocops3gp9phz4jc3 
                                           | s94qy2bqkpnqqumbxck | l45fdj1kcz0x06i9k | sqy4k5rpyr8won7x_a3h | m5fgnytsm5kbh2sbrzf; 

  wire mr9h2nuumis0_vx1kbbu849xvlx89du725kw = xh3sniad_mq0m5j2ilk | stw6xp6m1y7hi5xy | sganc4k2sd9qhhyt | qcbi1__w_lbxar86
                                     | m668z5d_2pgvlzqtt0r | f5obla9jfvqtwy50zglh | yxhb2hnxchdqcag9u9 | af7cl38e7futiwz7m5   
                                     | g9bfl499lfhirrrjln | g2esflomposu_jm | nn04ut84g694dyj3ngt | fx8tfw6ht51x591xovf
                                     | d1knhe17l7248qdlx3d | tdtkoiumk_q1_zlrgx1n_ | m06_keb0crbj3pkd_ | yo0gy1w6lzj_sxzxb0a
                                     | dserv0gb0p2c2yof | g2625iw5_kvvco4hf | xdtf0ycp133xtiom9 | fimif9coi4wgjje86n652
                                     | g690wip_77275ygun | eo1ocops3gp9phz4jc3 | akky00pxrb96le0sige5g | s94qy2bqkpnqqumbxck 
                                     | ds6le0delcgakxcymi | kjwyayvk_cqc5s0li40i | l45fdj1kcz0x06i9k | m5fgnytsm5kbh2sbrzf
                                     | dogjt36yta_opjg | k8wg766owq6fcetyyuo 
                                     | e65i99f2zhb74wze9lg | sqy4k5rpyr8won7x_a3h
                                     ;

  wire k0ly3yt_k96klqrmoe2jg2fjd6qz2edc5j87l =  n61z5eg85z3qt6ym | w6ojhbqk3lmsoe464 
                                        | ngyb9j0p18mjlul4  | no41cqtslidyozjc3b4| yo4avylbzg3xikezi | zuhncrmyvsvqe31yah | z1u9mb0is61kapi| hjj29yefty1oa5g1 
                                        | fgg6hxc67s_zufvn | bx8ta8ntqmkd296igjj5cm | qo4hl0cqzct4xyimucu | i92ohq_11aclejsw9
                                        ;

  wire tivrapwmioo0momgw9hmmlzhrcqyoa8a6wdu2yh =  tpxnwqn02te7dxkfod1c | l47a5b8y1b7jw87t
                                        | zociru6_rc45yinp5k | f3zsw2wieuvu92v24b | q7cxn6cfqixhf1j5c  | ytpvnxr5ldhrfhe
                                        | wyzwj_3yh41jvmcgv | as106js7z_6a17kl | dgoqvucxrbc7u23zbh1| k7u3ztuoje2dfwlb 
                                        | x7i6k3jtvgugfgwm | cmayk4nyxf2fgdyrgbdm | gkfxs8wvvzhw35g2w | lihv1jjl5cbn0k8m1 
                                        | ogxv3q5tyb1genv51czg | jqc0fopjngrnmrha1ca9 | nris9imni2zozl_9adll
                                        ;
  wire s89z9cptleb2csl1iyj0lg_altgx5k1f6316m1h = x43fhodherbcf_w4w | d_t7c_en995wivae5jc6g 
                                           ;
  wire oy_6emad9374dtcw5eu89i4o6o5kuiqu26hsgcb = hc6mrm8abcf82sqypnsn | tsfbnnx02_rdxvvpvk5a
                                           | r0oo_zmre7ja5s9h  | o63p86lpcfcy7xuj55
                                           ;
  wire isxv0tqhyam =
                    | qo4hl0cqzct4xyimucu | jqc0fopjngrnmrha1ca9 | nris9imni2zozl_9adll | g9bfl499lfhirrrjln | g2esflomposu_jm | nn04ut84g694dyj3ngt | fx8tfw6ht51x591xovf
                    | d1knhe17l7248qdlx3d | tdtkoiumk_q1_zlrgx1n_ | m06_keb0crbj3pkd_ | yo0gy1w6lzj_sxzxb0a | mtjkl28_lqkguy1g96p4 | d_rtbt5u2waj29pq38aw | gp2roes6p_wvpktfh
                    | rhpud0ssrcsrol8rx8nu4 | p57xv2ht1u5oz2jyd9m | yikkze0bi4xdf5kgp | ewo2z4ywjzk3rqw0c9di | w6ojhbqk3lmsoe464 | l47a5b8y1b7jw87t | f3zsw2wieuvu92v24b
                    | sv78kz_4osrj8ymh53m | zdwvt5v7m2azz1zncqlz | l_5fge2sjzcghz15 | ikrh3ggnb20z70nz | drexvwdx10vfyckm2w | hjj29yefty1oa5g1 | dgoqvucxrbc7u23zbh1
                    | k7u3ztuoje2dfwlb | fgg6hxc67s_zufvn | bx8ta8ntqmkd296igjj5cm | x7i6k3jtvgugfgwm | cmayk4nyxf2fgdyrgbdm | z1u9mb0is61kapi | m668z5d_2pgvlzqtt0r
                    | f5obla9jfvqtwy50zglh | yxhb2hnxchdqcag9u9 | af7cl38e7futiwz7m5 | os5cdj3yxqxq58sz | neja7y5h1cux76u7ru | uxstixgq52wcp394s2bq | ata32ab_8ia7entoq1d | wxfxhstnh27mwfsba43x
                    | g1bqvr3iwplkb20wpvq | cflo9l4odlq3l0so | aw1b57cswb2mmub | jv62xshm61xc3633g | casdl4x6djchiuqej | eaqgia_mu1yu9vo2nszk
                    
                    | x43fhodherbcf_w4w |  hc6mrm8abcf82sqypnsn |  tsfbnnx02_rdxvvpvk5a
                    | nhxdacdf6m8xlgp0gi | xdtf0ycp133xtiom9 | fimif9coi4wgjje86n652
                    | akky00pxrb96le0sige5g | s94qy2bqkpnqqumbxck | ds6le0delcgakxcymi | kjwyayvk_cqc5s0li40i 
                    | l45fdj1kcz0x06i9k | e65i99f2zhb74wze9lg | sqy4k5rpyr8won7x_a3h
                    ;

  wire qhmdzlcppcq8 = isxv0tqhyam | ccb88tt72pm4kk3aiztl_ | aquf29t5dbq4elt;
  wire pcdpwbqiqrxvx76lbm7p0 =
                             neja7y5h1cux76u7ru  | peoqulwt1lrkwd | tgghwgdy9ilyjs3vanp8 | py50qt89qihhrq6frt60
                           | uxmg0dt8ik73agsf | emfepzk_i3iart3w | d1knhe17l7248qdlx3d | tdtkoiumk_q1_zlrgx1n_ 
                           | m06_keb0crbj3pkd_  | yo0gy1w6lzj_sxzxb0a  
                           ;
 wire gdebc5b6o6bv57ax1bw = (~pcdpwbqiqrxvx76lbm7p0); 

  wire [23-1:0] nhqiwwnz4lmleg;
  assign  nhqiwwnz4lmleg[3:0]           = 4'd10;
  assign  nhqiwwnz4lmleg[4:4]          = vlfahv69;
  assign  nhqiwwnz4lmleg[5]    = pmmtjgnf20j2o_r;
  assign  nhqiwwnz4lmleg[6]   = wgjot58w1__ndyr81f;
  assign  nhqiwwnz4lmleg[7]    = py50qt89qihhrq6frt60;
  assign  nhqiwwnz4lmleg[8]   = uxmg0dt8ik73agsf;
  assign  nhqiwwnz4lmleg[9]     = x9o36wx2sxi_96riv;
  assign  nhqiwwnz4lmleg[10]    = l2mrfrrlbbj8wb25j;
  assign  nhqiwwnz4lmleg[11]     = sx2u7wkkrnzxotilhg;
  assign  nhqiwwnz4lmleg[12]    = jjudyrfeov9o45jiy;
  assign  nhqiwwnz4lmleg[13]     = peoqulwt1lrkwd;
  assign  nhqiwwnz4lmleg[14]    = tgghwgdy9ilyjs3vanp8;
  assign  nhqiwwnz4lmleg[15]      = y5g_0z60_kaqxvn1;
  assign  nhqiwwnz4lmleg[16]     = xdg0xfnp9f4p17fux;
  assign  nhqiwwnz4lmleg[17]     = g_k_2hcsq4fllbhbyvp;
  assign  nhqiwwnz4lmleg[18]     = fy_5mx58b8k0rbva;
  assign  nhqiwwnz4lmleg[19]     = mbbkhwc6igem3g;
  assign  nhqiwwnz4lmleg[20]     = w8kkipg2caprcl38r;
  assign  nhqiwwnz4lmleg[21]     = b4z_up9nkirbcj3jl;
  assign  nhqiwwnz4lmleg[22]     = xpa9jhun_nud6epww;

  wire [105-1:0] w98a0gvni829u3;
  assign w98a0gvni829u3[48]     = n61z5eg85z3qt6ym;
  assign w98a0gvni829u3[49]     = tpxnwqn02te7dxkfod1c;
  assign w98a0gvni829u3[50]     = zociru6_rc45yinp5k;
  assign w98a0gvni829u3[68]    = d_t7c_en995wivae5jc6g;
  assign w98a0gvni829u3[69]    = r0oo_zmre7ja5s9h;
  assign w98a0gvni829u3[70]    = o63p86lpcfcy7xuj55;
  assign w98a0gvni829u3[71]    = i92ohq_11aclejsw9;
  assign w98a0gvni829u3[72]    = lihv1jjl5cbn0k8m1;
  assign w98a0gvni829u3[73]    = ogxv3q5tyb1genv51czg;
  assign w98a0gvni829u3[74 ]    = htdih4lhmspfu8_ ;
  assign w98a0gvni829u3[75 ]    = dserv0gb0p2c2yof ;
  assign w98a0gvni829u3[76 ]    = g2625iw5_kvvco4hf ;
  assign  w98a0gvni829u3[3:0]           = 4'd11;
  assign  w98a0gvni829u3[4:4]          = vlfahv69;
  assign  w98a0gvni829u3[7]    = sganc4k2sd9qhhyt;
  assign  w98a0gvni829u3[6]     = m668z5d_2pgvlzqtt0r;
  assign  w98a0gvni829u3[5]    = f5obla9jfvqtwy50zglh;
  assign  w98a0gvni829u3[8]     = yxhb2hnxchdqcag9u9;
  assign  w98a0gvni829u3[9]    = af7cl38e7futiwz7m5;
  assign  w98a0gvni829u3[10]   = qcbi1__w_lbxar86;
  assign  w98a0gvni829u3[11]    = zuhncrmyvsvqe31yah;
  assign  w98a0gvni829u3[12]    = as106js7z_6a17kl;
  assign  w98a0gvni829u3[13]    = z1u9mb0is61kapi;
  assign  w98a0gvni829u3[14]   = hjj29yefty1oa5g1;
  assign  w98a0gvni829u3[15]    = dgoqvucxrbc7u23zbh1;
  assign  w98a0gvni829u3[16]   = k7u3ztuoje2dfwlb;
  assign  w98a0gvni829u3[17]   = yo4avylbzg3xikezi;
  assign  w98a0gvni829u3[18]   = wyzwj_3yh41jvmcgv;
  assign  w98a0gvni829u3[19]   = fgg6hxc67s_zufvn;
  assign  w98a0gvni829u3[20]  = bx8ta8ntqmkd296igjj5cm;
  assign  w98a0gvni829u3[21]   = x7i6k3jtvgugfgwm;
  assign  w98a0gvni829u3[22]  = cmayk4nyxf2fgdyrgbdm;
  assign  w98a0gvni829u3[25]      = pp7lw68tzorrt1ry;
  assign  w98a0gvni829u3[26]     = qwszvnfbt4kifn;
  assign  w98a0gvni829u3[27]      = l8skguypzoiw9k;
  assign  w98a0gvni829u3[28]     = bqonmn9o0yi3pta98ja;
  assign  w98a0gvni829u3[29]     = zse6ubdm7b85h4fv;
  assign  w98a0gvni829u3[30]     = w6ojhbqk3lmsoe464;
  assign  w98a0gvni829u3[31]     = l47a5b8y1b7jw87t;
  assign  w98a0gvni829u3[32]     = f3zsw2wieuvu92v24b;
  assign  w98a0gvni829u3[33]     = ata32ab_8ia7entoq1d;
  assign  w98a0gvni829u3[34]    = wxfxhstnh27mwfsba43x;
  assign  w98a0gvni829u3[35]     = g1bqvr3iwplkb20wpvq;
  assign  w98a0gvni829u3[36]    = cflo9l4odlq3l0so;
  assign  w98a0gvni829u3[37]    = aw1b57cswb2mmub;
  assign  w98a0gvni829u3[38]     = jv62xshm61xc3633g;
  assign  w98a0gvni829u3[39]    = casdl4x6djchiuqej;
  assign  w98a0gvni829u3[40]     = os5cdj3yxqxq58sz;
  assign  w98a0gvni829u3[41]     = neja7y5h1cux76u7ru;
  assign  w98a0gvni829u3[42]   = uxstixgq52wcp394s2bq;
  assign  w98a0gvni829u3[43]    = sv78kz_4osrj8ymh53m;
  assign  w98a0gvni829u3[44]    = zdwvt5v7m2azz1zncqlz;
  assign  w98a0gvni829u3[45]    = l_5fge2sjzcghz15;
  assign  w98a0gvni829u3[46]   = ikrh3ggnb20z70nz;
  assign  w98a0gvni829u3[47]   = drexvwdx10vfyckm2w;
  assign  w98a0gvni829u3[51]      = gkfxs8wvvzhw35g2w;
  assign  w98a0gvni829u3[52]    = qo4hl0cqzct4xyimucu;
  assign  w98a0gvni829u3[53]    = jqc0fopjngrnmrha1ca9;
  assign  w98a0gvni829u3[54]    = nris9imni2zozl_9adll;
  assign  w98a0gvni829u3[60]    = g9bfl499lfhirrrjln;
  assign  w98a0gvni829u3[61]    = g2esflomposu_jm;
  assign  w98a0gvni829u3[62]    = nn04ut84g694dyj3ngt;
  assign  w98a0gvni829u3[63]    = fx8tfw6ht51x591xovf;
  assign  w98a0gvni829u3[64]   = d1knhe17l7248qdlx3d;
  assign  w98a0gvni829u3[65]   = tdtkoiumk_q1_zlrgx1n_;
  assign  w98a0gvni829u3[66]    = m06_keb0crbj3pkd_;
  assign  w98a0gvni829u3[67]    = yo0gy1w6lzj_sxzxb0a;
  assign  w98a0gvni829u3[95]     = aquf29t5dbq4elt    ;
  assign  w98a0gvni829u3[96]    = eaqgia_mu1yu9vo2nszk   ;
  assign  w98a0gvni829u3[23]    = mtjkl28_lqkguy1g96p4;
  assign  w98a0gvni829u3[24]   = d_rtbt5u2waj29pq38aw;
  assign  w98a0gvni829u3[57]   = ewo2z4ywjzk3rqw0c9di;
  assign  w98a0gvni829u3[55]    = gp2roes6p_wvpktfh;
  assign  w98a0gvni829u3[56]   = rhpud0ssrcsrol8rx8nu4;
  assign  w98a0gvni829u3[58]    = p57xv2ht1u5oz2jyd9m;
  assign  w98a0gvni829u3[59]   = yikkze0bi4xdf5kgp;
  assign  w98a0gvni829u3[97]     = stw6xp6m1y7hi5xy;
  assign  w98a0gvni829u3[98]    = xh3sniad_mq0m5j2ilk;
  assign  w98a0gvni829u3[99]     = ngyb9j0p18mjlul4;
  assign  w98a0gvni829u3[100]     = q7cxn6cfqixhf1j5c;
  assign  w98a0gvni829u3[101]    = no41cqtslidyozjc3b4;
  assign  w98a0gvni829u3[102]    = ytpvnxr5ldhrfhe;
  assign  w98a0gvni829u3[103]    = emfepzk_i3iart3w;
  assign  w98a0gvni829u3[104]   = bpctswvy4clemt9h;
  assign  w98a0gvni829u3[77]  = x43fhodherbcf_w4w;
  assign  w98a0gvni829u3[78]  = hc6mrm8abcf82sqypnsn;
  assign  w98a0gvni829u3[79]  = tsfbnnx02_rdxvvpvk5a;
  assign  w98a0gvni829u3[80 ]  = nhxdacdf6m8xlgp0gi;
  assign  w98a0gvni829u3[81 ]  = xdtf0ycp133xtiom9;
  assign  w98a0gvni829u3[82 ]  = fimif9coi4wgjje86n652;
  assign  w98a0gvni829u3[83 ]  = akky00pxrb96le0sige5g;
  assign  w98a0gvni829u3[84]  = s94qy2bqkpnqqumbxck;
  assign  w98a0gvni829u3[85  ]  = g690wip_77275ygun;
  assign  w98a0gvni829u3[86 ]  = eo1ocops3gp9phz4jc3;
  assign  w98a0gvni829u3[87 ]  = ds6le0delcgakxcymi;
  assign  w98a0gvni829u3[88]  = kjwyayvk_cqc5s0li40i;
  assign  w98a0gvni829u3[89]  = l45fdj1kcz0x06i9k;
  assign  w98a0gvni829u3[90 ]  = e65i99f2zhb74wze9lg;
  assign  w98a0gvni829u3[91]  = sqy4k5rpyr8won7x_a3h;
  assign  w98a0gvni829u3[92  ]  = dogjt36yta_opjg;
  assign  w98a0gvni829u3[93 ]  = k8wg766owq6fcetyyuo;
  assign  w98a0gvni829u3[94 ]  = m5fgnytsm5kbh2sbrzf;

  


  wire zwwawd7qp5fytirkxl7jq9 = uk0ahn6nnbba7 == 7'b0011001;
  wire x_c94bnppi8ngabfz2iw = uk0ahn6nnbba7 == 7'b0011010;    
  wire wnw9q4wbzz7l6o9hrj4mh0 = uk0ahn6nnbba7 == 7'b0011110;    
  wire oezo_lnpso_pe9xd5gp = uk0ahn6nnbba7 == 7'b1000001;   
  wire xx5u6vajn90lcpxcfi_d26 = uk0ahn6nnbba7 == 7'b1000000;   
  wire mvw4y_tgvq9mm6qumk = uk0ahn6nnbba7 == 7'b1001001;   
  wire tibdvktu29n8xskpw3bmj = uk0ahn6nnbba7 == 7'b1001000;   
  wire i36pvh6w3hnu_emqkln = uk0ahn6nnbba7 == 7'b0000010;   
  wire n32bsi8b7sx1l4j93oy = uk0ahn6nnbba7 == 7'b0001010;   
  wire pwap35izr3ob3wmq64wu7 = uk0ahn6nnbba7 == 7'b0000011;   
  wire aaqwysz6l35fjqvf53x2w_7 = uk0ahn6nnbba7 == 7'b0001011;   
  wire ir_e6u4eazbj13c944p = uk0ahn6nnbba7 == 7'b0011000;

  wire mae_6a_pxmep9hv     = flv_cd606fxf7i739917y8 & ezupw6o2yfm5ojugrc3 & t61y7hkwkrvm7s ;
  wire vjw25i19dpz3    = mso_1l7nnv4ac14pv6qh & ezupw6o2yfm5ojugrc3 & t61y7hkwkrvm7s ;
  wire k9vvweo5_a_q_ip2l   = f6kcevztmpqpnc8xp3_r4 & ezupw6o2yfm5ojugrc3 & t61y7hkwkrvm7s ;
  wire w3njc277ysi3uz1    = duf6qt_vm6jkmkv9xu9 & ezupw6o2yfm5ojugrc3 & t61y7hkwkrvm7s ;
  wire g8wclh3x6xlwa3ncq   = m33lelq8_5u26vfl7hl6z & ezupw6o2yfm5ojugrc3 & t61y7hkwkrvm7s ;
  wire go4w_xvuj1m     = rc04_8vnldazobtsw8nkr8 & ezupw6o2yfm5ojugrc3 & t61y7hkwkrvm7s ;
  wire swvisnb87cxn83z    = xfrai8f3331hb4z5ww5_ & ezupw6o2yfm5ojugrc3 & t61y7hkwkrvm7s ;
  wire hp66bsfn_5mnw7gw6   = toaowsb_5w3arwmyl2 & ezupw6o2yfm5ojugrc3 & t61y7hkwkrvm7s ;
  wire szsij0guhgpj    = cvhx1ne2we07dkbzbpwakl & ezupw6o2yfm5ojugrc3 & t61y7hkwkrvm7s ;
  wire hugyxq6gvlbt7tp   = amf97jdmi0f4r4z2kmw & ezupw6o2yfm5ojugrc3 & t61y7hkwkrvm7s ;
  wire tpv9dscg_ntzh_rhh4   = rh5f36cuohtogtfizd & ezupw6o2yfm5ojugrc3 & t61y7hkwkrvm7s ;
  wire b0wowenfcyq_6_e  = jhbiy5xf0ygws7apfg03 & ezupw6o2yfm5ojugrc3 & t61y7hkwkrvm7s ;
  wire c784pnrp9fe0jg6ne39  = b12f43e4j_bhgigw_xvwmqe & ezupw6o2yfm5ojugrc3 & t61y7hkwkrvm7s ;
  wire kc_yoe3swf_o07x7p  = i_nd_auanr4nliiv9ru_mjy & ezupw6o2yfm5ojugrc3 & t61y7hkwkrvm7s ;
  wire ugiayevhrf3oqht9  = ha7x94wp2o8bpzvtiq_d & ezupw6o2yfm5ojugrc3 & t61y7hkwkrvm7s ;
  wire higk3ii9e9i_f    = crhfv2tcnpzr02ktjbc & ezupw6o2yfm5ojugrc3 & t61y7hkwkrvm7s ;
  wire g6_j6lr4ti9yu    = vubg64i36fbtxkcl4s776lk & ezupw6o2yfm5ojugrc3 & t61y7hkwkrvm7s ;
  wire jr97br_y15cmo2ku    = hmrtc229uz_sqjxkb8myxe & ezupw6o2yfm5ojugrc3 & t61y7hkwkrvm7s ;
  wire k0tmdbnsotlk    = gankodz2wzpdwh5hez & ezupw6o2yfm5ojugrc3 & t61y7hkwkrvm7s ;
  wire hfqcy171lm219z2    = styktg7w7fi36jw0e5n4h93 & jzb70ho_u3wii0cb_zw & ezupw6o2yfm5ojugrc3 & t61y7hkwkrvm7s;
  wire gjhl0yua7khqyyj7    = bepkj4gbb77isq3_v9 & ezupw6o2yfm5ojugrc3 & t61y7hkwkrvm7s ;
  wire n7z6su9ff17vc26hu   = lrptc0hyjyd7hdoypa0_g & ezupw6o2yfm5ojugrc3 & t61y7hkwkrvm7s ;
  wire rp86b05b7wi0gsy7np  = i6fh1oflvwwzfgicny1c & ezupw6o2yfm5ojugrc3 & t61y7hkwkrvm7s ;
  wire jt75suen_okjf02   = e9hn3j9k88f8miq238hz1 & ezupw6o2yfm5ojugrc3 & t61y7hkwkrvm7s ;
  wire uoy8pb4b3_q04van  = ir_e6u4eazbj13c944p & ezupw6o2yfm5ojugrc3 & t61y7hkwkrvm7s ;
  wire esnmi_yufd7l1af    = uncepq376ovruspfffvl5 & ezupw6o2yfm5ojugrc3 & t61y7hkwkrvm7s ;
  wire hp3zdh34mwyu_   = t6_6ypj94nny67ise0x9 & ezupw6o2yfm5ojugrc3 & t61y7hkwkrvm7s ;
  wire quh0wjpu8_60_00  = i0ahgxc7hvmvc1hsbq8 & ezupw6o2yfm5ojugrc3 & t61y7hkwkrvm7s ;
  wire yyq89zr8ntwjgvv9dh   = pvy429fepo5d_7j0eq5ky & ezupw6o2yfm5ojugrc3 & t61y7hkwkrvm7s ;
  wire blezqucpbhjpa4v9  = zwwawd7qp5fytirkxl7jq9 & ezupw6o2yfm5ojugrc3 & t61y7hkwkrvm7s ;
  wire o5obw4mzrir4f2ofd   = xvbpjhbrdw506s4r5je_v & ezupw6o2yfm5ojugrc3 & t61y7hkwkrvm7s ;    
  wire osn82rwdapvn3cunh  = i36pvh6w3hnu_emqkln & ezupw6o2yfm5ojugrc3 & t61y7hkwkrvm7s ;    
  wire jto_jycd4wmbzar = lipdgvrqr439y_cnsv & ezupw6o2yfm5ojugrc3 & t61y7hkwkrvm7s ;    
  wire d4roaqpdp0v1368y  = n32bsi8b7sx1l4j93oy & ezupw6o2yfm5ojugrc3 & t61y7hkwkrvm7s ;    
  wire owqgxd_mnoeuh58 = x_c94bnppi8ngabfz2iw & ezupw6o2yfm5ojugrc3 & t61y7hkwkrvm7s ;    
  wire vq0ayiqnvwy2exgn   = umom31fkh4dmsle8dt & ezupw6o2yfm5ojugrc3 & t61y7hkwkrvm7s ;    
  wire yrp4tnx0z0vr9if  = pwap35izr3ob3wmq64wu7 & ezupw6o2yfm5ojugrc3 & t61y7hkwkrvm7s ;    
  wire bha_2ihvu1x5vf6 = veb9c0lxewgh_4qiy5 & ezupw6o2yfm5ojugrc3 & t61y7hkwkrvm7s ;    
  wire rrlsg7zpsrnhfxb  = aaqwysz6l35fjqvf53x2w_7 & ezupw6o2yfm5ojugrc3 & t61y7hkwkrvm7s ;    
  wire krefblqj6lij3t4p = fr9vuzzy67toa8_rpz_ & ezupw6o2yfm5ojugrc3 & t61y7hkwkrvm7s ;    
  wire k06e5l0uw9wzwp2it   = sketktuyfh2vxjbshrr & t8jc64yc1l6q8eclq_c & t61y7hkwkrvm7s ;    
  wire ha32lltdxd7x19  = ef0qt3ctq84209xo8ti63mv & t8jc64yc1l6q8eclq_c & t61y7hkwkrvm7s ;    
  wire itt7e1z4g56bjpzdcq = q1g4g81fl48iq3ndywfle3 & t8jc64yc1l6q8eclq_c & t61y7hkwkrvm7s ;    
  wire m52a83vna7cr18mdn  = rgjf1vrs4iai2hif_09x & t8jc64yc1l6q8eclq_c & t61y7hkwkrvm7s ;    
  wire c80ogd8uqs8qta9l1ev = brnnngwkv59w2kz9usv3k8 & t8jc64yc1l6q8eclq_c & t61y7hkwkrvm7s ;    
  wire z53vzzym9v5v6   = a70w9nx14ytij6ok0iq & t8jc64yc1l6q8eclq_c & t61y7hkwkrvm7s ;    
  wire ns6x4s_o3pi6ax2n  = zpue29q3_sghsyln86mp & t8jc64yc1l6q8eclq_c & t61y7hkwkrvm7s ;    
  wire nb0wrp9_4ugc6qkjx7 = tgij_tz20n4mlmn8gc & t8jc64yc1l6q8eclq_c & t61y7hkwkrvm7s ;    
  wire z5bi2emm96esv_geki  = qcpti7i25_4w_aexyk1 & t8jc64yc1l6q8eclq_c & t61y7hkwkrvm7s ;    
  wire jmbuhj5mdexw1m3uqq = wp2e1icm345eqoi7xse0mo & t8jc64yc1l6q8eclq_c & t61y7hkwkrvm7s ;
  wire lnchd6wpif2lsuic_  = jysojps4nkgwbif943 & ezupw6o2yfm5ojugrc3 & t61y7hkwkrvm7s ;    
  wire v2k3hrn_5xg64b7aocn = fcpfa9hp28k7bapl82 & ezupw6o2yfm5ojugrc3 & t61y7hkwkrvm7s ;    
  wire akr76mirt0394rwypu = hx3wrp4j8s1ov27syy & ezupw6o2yfm5ojugrc3 & t61y7hkwkrvm7s ;    
  wire mckx1mltgmxacp_ = naged_b50dbpmu745zp & ezupw6o2yfm5ojugrc3 & t61y7hkwkrvm7s ;    
  wire typ6wj08ixws3lsuso = wnw9q4wbzz7l6o9hrj4mh0 & ezupw6o2yfm5ojugrc3 & t61y7hkwkrvm7s ;    
  wire ijvh48b4xaa54zh   = oezo_lnpso_pe9xd5gp & ezupw6o2yfm5ojugrc3 & t61y7hkwkrvm7s ;   
  wire qawzrnnnqu9zw8   = xx5u6vajn90lcpxcfi_d26 & ezupw6o2yfm5ojugrc3 & t61y7hkwkrvm7s ;   
  wire k4x3xpwe9_94trje   = mvw4y_tgvq9mm6qumk & ezupw6o2yfm5ojugrc3 & t61y7hkwkrvm7s ;   
  wire eytzcjin8i_o7qgg2g   = tibdvktu29n8xskpw3bmj & ezupw6o2yfm5ojugrc3 & t61y7hkwkrvm7s ;   
  wire ecccb2oy3kp6vbt   = styktg7w7fi36jw0e5n4h93 & auauwu7otyuaf2eindwrip & ezupw6o2yfm5ojugrc3 & t61y7hkwkrvm7s;
  wire xnb761cg1sb1d    = i36pvh6w3hnu_emqkln & d24iqtxvb2trplxk2m & t61y7hkwkrvm7s ;   
  wire e02lkx_fya1ouym7h   = n32bsi8b7sx1l4j93oy & d24iqtxvb2trplxk2m & t61y7hkwkrvm7s ;   
  wire elcvhpi2hcg0    = pwap35izr3ob3wmq64wu7 & d24iqtxvb2trplxk2m & t61y7hkwkrvm7s ;   
  wire n8r0676nkk3s04b7   = aaqwysz6l35fjqvf53x2w_7 & d24iqtxvb2trplxk2m & t61y7hkwkrvm7s ;   
  wire m3fice1xap_p463s    = lrptc0hyjyd7hdoypa0_g & d24iqtxvb2trplxk2m & t61y7hkwkrvm7s ; 
  wire et2vvn5b9hs2dsxc   = e9hn3j9k88f8miq238hz1 & d24iqtxvb2trplxk2m & t61y7hkwkrvm7s ; 
  wire q92dtkdebjot0e    = i6fh1oflvwwzfgicny1c & d24iqtxvb2trplxk2m & t61y7hkwkrvm7s ;
  wire dpm72l5g2io4k   = ir_e6u4eazbj13c944p & d24iqtxvb2trplxk2m & t61y7hkwkrvm7s ;
  wire lf8nodmhavxf    = t6_6ypj94nny67ise0x9 & d24iqtxvb2trplxk2m & t61y7hkwkrvm7s ;
  wire ta99gbty1xpqs6_ahm   = pvy429fepo5d_7j0eq5ky & d24iqtxvb2trplxk2m & t61y7hkwkrvm7s ;   
  wire blk15yrqxkt8zs2br    = i0ahgxc7hvmvc1hsbq8 & d24iqtxvb2trplxk2m & t61y7hkwkrvm7s ;  
  wire phiws9b8v856wgd   = zwwawd7qp5fytirkxl7jq9 & d24iqtxvb2trplxk2m & t61y7hkwkrvm7s ;  
  wire fj50cc2xxbpn     = rf284mrjg_bqa1hj60swyf & ezupw6o2yfm5ojugrc3 & t61y7hkwkrvm7s ; 
  wire uavbu3i6ubzz     = v3hylq_n52mziras6qen & ezupw6o2yfm5ojugrc3 & t61y7hkwkrvm7s ; 
  wire dsp656i_shm9fbrjf    = styktg7w7fi36jw0e5n4h93 & c6svrw070n8tv5npikqj18 & ezupw6o2yfm5ojugrc3 & t61y7hkwkrvm7s;
  wire fklgk6eyb2vd8    = l6zyb5b3_f8uuon8o3p	& d24iqtxvb2trplxk2m & t61y7hkwkrvm7s ;
  wire zfotdct2of6_kc   = xx5u6vajn90lcpxcfi_d26	& d24iqtxvb2trplxk2m & t61y7hkwkrvm7s ;
  wire k1oqlvc677n04h94z31  = c7npl5770szduubj6_grim	& d24iqtxvb2trplxk2m & t61y7hkwkrvm7s ;
  wire wean5xmif_myv   = tibdvktu29n8xskpw3bmj	& d24iqtxvb2trplxk2m & t61y7hkwkrvm7s ;
  wire qzptr55gc1d815k  = d9gmx9ccvp0rgcy7n_ii	& d24iqtxvb2trplxk2m & t61y7hkwkrvm7s ;
  wire fouln9y77frzodomf    = c9xaw73uh3hmihrn801brf	& d24iqtxvb2trplxk2m & t61y7hkwkrvm7s ;
  wire ot7hpozxj594mxo0o8   = oezo_lnpso_pe9xd5gp	& d24iqtxvb2trplxk2m & t61y7hkwkrvm7s ;
  wire q9uit_5jup8pgp6l  = whvtopzve8q_t001lyx	& d24iqtxvb2trplxk2m & t61y7hkwkrvm7s ;
  wire hked2y47eglmii   = mvw4y_tgvq9mm6qumk	& d24iqtxvb2trplxk2m & t61y7hkwkrvm7s ;
  wire utvej5knrsiltp5b  = vrn4ssw1i97fztoyaq5kq	& d24iqtxvb2trplxk2m & t61y7hkwkrvm7s ;
  wire r2icw20xk206b      = k_h8qestuhin60n5ckxmkfx & ezupw6o2yfm5ojugrc3 & t61y7hkwkrvm7s ;
  wire tv4hqiny5afky9w   = 1'b0; 
  wire vwmbmpalhwfnoi_0g  = 1'b0; 
  wire we6wj_afzuesr1zwnl   = 1'b0; 
  wire jzbjl5cnc_hb5hixv  = 1'b0; 
  wire qusz_xa0ku_toij493   = 1'b0; 
  wire bi0wblozr4jb8yf4  = 1'b0; 
                       
  wire olzyli2shf6m0eu    = bepkj4gbb77isq3_v9 & t8jc64yc1l6q8eclq_c & t61y7hkwkrvm7s ;
  wire r7cnjrtmoa4z3wzm   = lrptc0hyjyd7hdoypa0_g & t8jc64yc1l6q8eclq_c & t61y7hkwkrvm7s ;
  wire xs9gkwo3sk9927f  = i6fh1oflvwwzfgicny1c & t8jc64yc1l6q8eclq_c & t61y7hkwkrvm7s ;
  wire t622z2sipa9amny   = e9hn3j9k88f8miq238hz1 & t8jc64yc1l6q8eclq_c & t61y7hkwkrvm7s ;
  wire gplqhxgap4qxw2585n  = ir_e6u4eazbj13c944p & t8jc64yc1l6q8eclq_c & t61y7hkwkrvm7s ;
  wire hd73e7ysgqar7d82    = uncepq376ovruspfffvl5 & t8jc64yc1l6q8eclq_c & t61y7hkwkrvm7s ;
  wire ouz2qqdkqv42w   = t6_6ypj94nny67ise0x9 & t8jc64yc1l6q8eclq_c & t61y7hkwkrvm7s ;
  wire i9k7gr9f1m5x4z9m7sw  = i0ahgxc7hvmvc1hsbq8 & t8jc64yc1l6q8eclq_c & t61y7hkwkrvm7s ;
  wire w1064psfmbve8hpe   = pvy429fepo5d_7j0eq5ky & t8jc64yc1l6q8eclq_c & t61y7hkwkrvm7s ;
  wire gisgif8kbt3puleu  = zwwawd7qp5fytirkxl7jq9 & t8jc64yc1l6q8eclq_c & t61y7hkwkrvm7s ;
  wire rnblmzik1pew6va2h   = xvbpjhbrdw506s4r5je_v & t8jc64yc1l6q8eclq_c & t61y7hkwkrvm7s ;    
  wire dimrfoq94vmw2xn1t  = i36pvh6w3hnu_emqkln & t8jc64yc1l6q8eclq_c & t61y7hkwkrvm7s ;    
  wire xppjwy_axpkzto1n_hs = lipdgvrqr439y_cnsv & t8jc64yc1l6q8eclq_c & t61y7hkwkrvm7s ;    
  wire ev_fa6s12jdsf7  = n32bsi8b7sx1l4j93oy & t8jc64yc1l6q8eclq_c & t61y7hkwkrvm7s ;    
  wire da7q3cxfn4d3s1k50 = x_c94bnppi8ngabfz2iw & t8jc64yc1l6q8eclq_c & t61y7hkwkrvm7s ;    
  wire dmzs8qjfkowxd   = umom31fkh4dmsle8dt & t8jc64yc1l6q8eclq_c & t61y7hkwkrvm7s ;    
  wire xq79ouq18ya2qxjmwx  = pwap35izr3ob3wmq64wu7 & t8jc64yc1l6q8eclq_c & t61y7hkwkrvm7s ;    
  wire xm5w1y9xnpmzt7_fp2aq = veb9c0lxewgh_4qiy5 & t8jc64yc1l6q8eclq_c & t61y7hkwkrvm7s ;    
  wire elkxwjgl9ny2u6k3dg  = aaqwysz6l35fjqvf53x2w_7 & t8jc64yc1l6q8eclq_c & t61y7hkwkrvm7s ;    
  wire g73i4v_qd7tqi0fc = fr9vuzzy67toa8_rpz_ & t8jc64yc1l6q8eclq_c & t61y7hkwkrvm7s ;    
  wire j_jcm4qgb9x62   = v3hylq_n52mziras6qen & t8jc64yc1l6q8eclq_c & t61y7hkwkrvm7s ;    
  wire cf2ndyjmh3psm0oe2  = d9gmx9ccvp0rgcy7n_ii & t8jc64yc1l6q8eclq_c & t61y7hkwkrvm7s ;    
  wire pcx1a0uxtq0mr8gyc = tx0e46vrruq3cgq9ghul4 & t8jc64yc1l6q8eclq_c & t61y7hkwkrvm7s ;    
  wire hu6futh2tv8zrpvuhbq  = l6zyb5b3_f8uuon8o3p & t8jc64yc1l6q8eclq_c & t61y7hkwkrvm7s ;    
  wire r7_qpw537yx2nx2tbsj = k_h8qestuhin60n5ckxmkfx & t8jc64yc1l6q8eclq_c & t61y7hkwkrvm7s ;    
  wire uxzv2w6nerfya6b   = rf284mrjg_bqa1hj60swyf & t8jc64yc1l6q8eclq_c & t61y7hkwkrvm7s ;    
  wire ky8_zvpu3hzcuwzma  = vrn4ssw1i97fztoyaq5kq & t8jc64yc1l6q8eclq_c & t61y7hkwkrvm7s ;    
  wire fffc565224sv9zh5bt9 = mnd8c7lvcdtsypyiygspg & t8jc64yc1l6q8eclq_c & t61y7hkwkrvm7s ;    
  wire q5kg_hwy37mzu95q  = c9xaw73uh3hmihrn801brf & t8jc64yc1l6q8eclq_c & t61y7hkwkrvm7s ;    
  wire kv6sfx3a9qhkrx75k = eu9j7rkhrocfjsewdf6mfvu & t8jc64yc1l6q8eclq_c & t61y7hkwkrvm7s ;    
  wire nwvvvndgm3k0n   = mvw4y_tgvq9mm6qumk & t8jc64yc1l6q8eclq_c & t61y7hkwkrvm7s ;   
  wire e_giw7b4ut0jmmpy9a   = tibdvktu29n8xskpw3bmj & t8jc64yc1l6q8eclq_c & t61y7hkwkrvm7s ;   
  wire z79y6w0q_w4smuqg   = whvtopzve8q_t001lyx & t8jc64yc1l6q8eclq_c & t61y7hkwkrvm7s ;   
  wire buou043vqauc4   = c7npl5770szduubj6_grim & t8jc64yc1l6q8eclq_c & t61y7hkwkrvm7s ;   
  wire v_b574hro993x   = styktg7w7fi36jw0e5n4h93 & pk4bj6ne4riq5l_gqv9maw_ & ezupw6o2yfm5ojugrc3 & t61y7hkwkrvm7s;

  assign upbbycb5makv3xss7d_ueoxns88bj =                           
                         | aquf29t5dbq4elt    
                         | eaqgia_mu1yu9vo2nszk   
                         ;

  wire qm17qduoi54r_53z; 
  wire vu8cn0tjzmmmjqj_9; 

  wire [54-1:0] wazt073vrvkujb_lpjze6;
  assign wazt073vrvkujb_lpjze6[3:0]           = 4'd8;
  assign wazt073vrvkujb_lpjze6[4:4]          = vlfahv69;
  assign wazt073vrvkujb_lpjze6[5     ] = mae_6a_pxmep9hv     ;
  assign wazt073vrvkujb_lpjze6[6    ] = vjw25i19dpz3    ;
  assign wazt073vrvkujb_lpjze6[7   ] = k9vvweo5_a_q_ip2l   ;
  assign wazt073vrvkujb_lpjze6[8    ] = w3njc277ysi3uz1    ;
  assign wazt073vrvkujb_lpjze6[10   ] = g8wclh3x6xlwa3ncq   ;
  assign wazt073vrvkujb_lpjze6[11     ] = go4w_xvuj1m     ;
  assign wazt073vrvkujb_lpjze6[12    ] = swvisnb87cxn83z    ;
  assign wazt073vrvkujb_lpjze6[13   ] = hp66bsfn_5mnw7gw6   ;
  assign wazt073vrvkujb_lpjze6[14    ] = szsij0guhgpj    ;
  assign wazt073vrvkujb_lpjze6[16   ] = hugyxq6gvlbt7tp   ;
  assign wazt073vrvkujb_lpjze6[17   ] = tpv9dscg_ntzh_rhh4   ;
  assign wazt073vrvkujb_lpjze6[18  ] = b0wowenfcyq_6_e  ;
  assign wazt073vrvkujb_lpjze6[19  ] = c784pnrp9fe0jg6ne39  ;
  assign wazt073vrvkujb_lpjze6[20  ] = kc_yoe3swf_o07x7p  ;
  assign wazt073vrvkujb_lpjze6[21  ] = ugiayevhrf3oqht9  ;
  assign wazt073vrvkujb_lpjze6[22    ] = higk3ii9e9i_f    ;
  assign wazt073vrvkujb_lpjze6[23    ] = g6_j6lr4ti9yu    ;
  assign wazt073vrvkujb_lpjze6[24    ] = jr97br_y15cmo2ku    ;
  assign wazt073vrvkujb_lpjze6[25    ] = k0tmdbnsotlk    ;
  assign wazt073vrvkujb_lpjze6[26    ] = hfqcy171lm219z2    ;
  assign wazt073vrvkujb_lpjze6[27   ] = tv4hqiny5afky9w   ;   
  assign wazt073vrvkujb_lpjze6[9   ] = we6wj_afzuesr1zwnl   ;
  assign wazt073vrvkujb_lpjze6[15   ] = qusz_xa0ku_toij493   ;
  assign wazt073vrvkujb_lpjze6[28    ] = xnb761cg1sb1d    ;   
  assign wazt073vrvkujb_lpjze6[29   ] = e02lkx_fya1ouym7h   ;   
  assign wazt073vrvkujb_lpjze6[30    ] = elcvhpi2hcg0    ;   
  assign wazt073vrvkujb_lpjze6[31   ] = n8r0676nkk3s04b7   ;   
  assign wazt073vrvkujb_lpjze6[32    ] = m3fice1xap_p463s    ; 
  assign wazt073vrvkujb_lpjze6[33   ] = et2vvn5b9hs2dsxc   ; 
  assign wazt073vrvkujb_lpjze6[34    ] = q92dtkdebjot0e    ;
  assign wazt073vrvkujb_lpjze6[35   ] = dpm72l5g2io4k   ;
  assign wazt073vrvkujb_lpjze6[36    ] = lf8nodmhavxf    ;
  assign wazt073vrvkujb_lpjze6[37   ] = ta99gbty1xpqs6_ahm   ;   
  assign wazt073vrvkujb_lpjze6[38    ] = blk15yrqxkt8zs2br    ;  
  assign wazt073vrvkujb_lpjze6[39   ] = phiws9b8v856wgd   ;  
  assign wazt073vrvkujb_lpjze6[40     ] = fj50cc2xxbpn     ; 
  assign wazt073vrvkujb_lpjze6[41     ] = uavbu3i6ubzz     ; 
  assign wazt073vrvkujb_lpjze6[42    ] = dsp656i_shm9fbrjf    ; 
  assign wazt073vrvkujb_lpjze6[43    ] = fklgk6eyb2vd8    ;
  assign wazt073vrvkujb_lpjze6[44   ] = zfotdct2of6_kc   ;   
  assign wazt073vrvkujb_lpjze6[45  ] = k1oqlvc677n04h94z31  ;  
  assign wazt073vrvkujb_lpjze6[46   ] = wean5xmif_myv   ;  
  assign wazt073vrvkujb_lpjze6[47  ] = qzptr55gc1d815k  ; 
  assign wazt073vrvkujb_lpjze6[48    ] = fouln9y77frzodomf    ; 
  assign wazt073vrvkujb_lpjze6[49   ] = ot7hpozxj594mxo0o8   ; 
  assign wazt073vrvkujb_lpjze6[50  ] = q9uit_5jup8pgp6l  ;
  assign wazt073vrvkujb_lpjze6[51   ] = hked2y47eglmii   ;
  assign wazt073vrvkujb_lpjze6[52  ] = utvej5knrsiltp5b  ;
  assign wazt073vrvkujb_lpjze6[53      ] = r2icw20xk206b      ;

  wire [48-1:0] azvwipii1valwcdp80j3_oq;
  assign azvwipii1valwcdp80j3_oq[3:0]           = 4'd9;
  assign azvwipii1valwcdp80j3_oq[4:4]          = vlfahv69;
  assign azvwipii1valwcdp80j3_oq[5    ] = gjhl0yua7khqyyj7    ;
  assign azvwipii1valwcdp80j3_oq[6   ] = n7z6su9ff17vc26hu   ;
  assign azvwipii1valwcdp80j3_oq[7  ] = rp86b05b7wi0gsy7np  ;
  assign azvwipii1valwcdp80j3_oq[8   ] = jt75suen_okjf02   ;
  assign azvwipii1valwcdp80j3_oq[10  ] = uoy8pb4b3_q04van  ;
  assign azvwipii1valwcdp80j3_oq[11    ] = esnmi_yufd7l1af    ;
  assign azvwipii1valwcdp80j3_oq[12   ] = hp3zdh34mwyu_   ;
  assign azvwipii1valwcdp80j3_oq[13  ] = quh0wjpu8_60_00  ;
  assign azvwipii1valwcdp80j3_oq[14   ] = yyq89zr8ntwjgvv9dh   ;
  assign azvwipii1valwcdp80j3_oq[16  ] = blezqucpbhjpa4v9  ;
  assign azvwipii1valwcdp80j3_oq[17   ] = o5obw4mzrir4f2ofd   ;    
  assign azvwipii1valwcdp80j3_oq[18  ] = osn82rwdapvn3cunh  ;    
  assign azvwipii1valwcdp80j3_oq[19 ] = jto_jycd4wmbzar ;    
  assign azvwipii1valwcdp80j3_oq[20  ] = d4roaqpdp0v1368y  ;    
  assign azvwipii1valwcdp80j3_oq[21 ] = owqgxd_mnoeuh58 ;    
  assign azvwipii1valwcdp80j3_oq[22   ] = vq0ayiqnvwy2exgn   ;    
  assign azvwipii1valwcdp80j3_oq[23  ] = yrp4tnx0z0vr9if  ;    
  assign azvwipii1valwcdp80j3_oq[24 ] = bha_2ihvu1x5vf6 ;    
  assign azvwipii1valwcdp80j3_oq[25  ] = rrlsg7zpsrnhfxb  ;    
  assign azvwipii1valwcdp80j3_oq[26 ] = krefblqj6lij3t4p ;    
  assign azvwipii1valwcdp80j3_oq[27   ] = k06e5l0uw9wzwp2it   ;    
  assign azvwipii1valwcdp80j3_oq[28  ] = ha32lltdxd7x19  ;    
  assign azvwipii1valwcdp80j3_oq[29 ] = itt7e1z4g56bjpzdcq ;    
  assign azvwipii1valwcdp80j3_oq[30  ] = m52a83vna7cr18mdn  ;    
  assign azvwipii1valwcdp80j3_oq[31 ] = c80ogd8uqs8qta9l1ev ;    
  assign azvwipii1valwcdp80j3_oq[32   ] = z53vzzym9v5v6   ;    
  assign azvwipii1valwcdp80j3_oq[33  ] = ns6x4s_o3pi6ax2n  ;    
  assign azvwipii1valwcdp80j3_oq[34 ] = nb0wrp9_4ugc6qkjx7 ;    
  assign azvwipii1valwcdp80j3_oq[35  ] = z5bi2emm96esv_geki  ;    
  assign azvwipii1valwcdp80j3_oq[36 ] = jmbuhj5mdexw1m3uqq ;    
  assign azvwipii1valwcdp80j3_oq[37  ] = lnchd6wpif2lsuic_  ;    
  assign azvwipii1valwcdp80j3_oq[38 ] = v2k3hrn_5xg64b7aocn ;    
  assign azvwipii1valwcdp80j3_oq[39 ] = akr76mirt0394rwypu ;    
  assign azvwipii1valwcdp80j3_oq[40 ] = mckx1mltgmxacp_ ;    
  assign azvwipii1valwcdp80j3_oq[41 ] = typ6wj08ixws3lsuso ;    
  assign azvwipii1valwcdp80j3_oq[42   ] = ijvh48b4xaa54zh   ;   
  assign azvwipii1valwcdp80j3_oq[43   ] = qawzrnnnqu9zw8   ;   
  assign azvwipii1valwcdp80j3_oq[44   ] = k4x3xpwe9_94trje   ;   
  assign azvwipii1valwcdp80j3_oq[45   ] = eytzcjin8i_o7qgg2g   ;   
  assign azvwipii1valwcdp80j3_oq[46   ] = ecccb2oy3kp6vbt   ;   
  assign azvwipii1valwcdp80j3_oq[9  ] = jzbjl5cnc_hb5hixv  ;
  assign azvwipii1valwcdp80j3_oq[47  ] = vwmbmpalhwfnoi_0g  ;   
  assign azvwipii1valwcdp80j3_oq[15  ] = bi0wblozr4jb8yf4  ;


  wire [40-1:0] no56h0p6kag9edi57joc3m;
  assign no56h0p6kag9edi57joc3m[3:0]           = 4'd9;
  assign no56h0p6kag9edi57joc3m[4:4]          = vlfahv69; 
  assign no56h0p6kag9edi57joc3m[5    ] = olzyli2shf6m0eu    ;
  assign no56h0p6kag9edi57joc3m[6   ] = r7cnjrtmoa4z3wzm   ;
  assign no56h0p6kag9edi57joc3m[7  ] = xs9gkwo3sk9927f  ;
  assign no56h0p6kag9edi57joc3m[8   ] = t622z2sipa9amny   ;
  assign no56h0p6kag9edi57joc3m[9  ] = gplqhxgap4qxw2585n  ;
  assign no56h0p6kag9edi57joc3m[10    ] = hd73e7ysgqar7d82    ;
  assign no56h0p6kag9edi57joc3m[11   ] = ouz2qqdkqv42w   ;
  assign no56h0p6kag9edi57joc3m[12  ] = i9k7gr9f1m5x4z9m7sw  ;
  assign no56h0p6kag9edi57joc3m[13   ] = w1064psfmbve8hpe   ;
  assign no56h0p6kag9edi57joc3m[14  ] = gisgif8kbt3puleu  ;
  assign no56h0p6kag9edi57joc3m[15   ] = rnblmzik1pew6va2h   ;    
  assign no56h0p6kag9edi57joc3m[16  ] = dimrfoq94vmw2xn1t  ;    
  assign no56h0p6kag9edi57joc3m[17 ] = xppjwy_axpkzto1n_hs ;    
  assign no56h0p6kag9edi57joc3m[18  ] = ev_fa6s12jdsf7  ;    
  assign no56h0p6kag9edi57joc3m[19 ] = da7q3cxfn4d3s1k50 ;    
  assign no56h0p6kag9edi57joc3m[20   ] = dmzs8qjfkowxd   ;    
  assign no56h0p6kag9edi57joc3m[21  ] = xq79ouq18ya2qxjmwx  ;    
  assign no56h0p6kag9edi57joc3m[22 ] = xm5w1y9xnpmzt7_fp2aq ;    
  assign no56h0p6kag9edi57joc3m[23  ] = elkxwjgl9ny2u6k3dg  ;    
  assign no56h0p6kag9edi57joc3m[24 ] = g73i4v_qd7tqi0fc ;    
  assign no56h0p6kag9edi57joc3m[25   ] = j_jcm4qgb9x62   ;    
  assign no56h0p6kag9edi57joc3m[26  ] = cf2ndyjmh3psm0oe2  ;    
  assign no56h0p6kag9edi57joc3m[27 ] = pcx1a0uxtq0mr8gyc ;    
  assign no56h0p6kag9edi57joc3m[28  ] = hu6futh2tv8zrpvuhbq  ;    
  assign no56h0p6kag9edi57joc3m[29 ] = r7_qpw537yx2nx2tbsj ;    
  assign no56h0p6kag9edi57joc3m[30   ] = uxzv2w6nerfya6b   ;    
  assign no56h0p6kag9edi57joc3m[31  ] = ky8_zvpu3hzcuwzma  ;    
  assign no56h0p6kag9edi57joc3m[32 ] = fffc565224sv9zh5bt9 ;    
  assign no56h0p6kag9edi57joc3m[33  ] = q5kg_hwy37mzu95q  ;    
  assign no56h0p6kag9edi57joc3m[34 ] = kv6sfx3a9qhkrx75k ;    
  assign no56h0p6kag9edi57joc3m[35   ] = nwvvvndgm3k0n   ;   
  assign no56h0p6kag9edi57joc3m[36   ] = e_giw7b4ut0jmmpy9a   ;   
  assign no56h0p6kag9edi57joc3m[37   ] = z79y6w0q_w4smuqg   ;   
  assign no56h0p6kag9edi57joc3m[38   ] = buou043vqauc4   ;   
  assign no56h0p6kag9edi57joc3m[39   ] = v_b574hro993x   ;   


  assign qm17qduoi54r_53z =
                            tv4hqiny5afky9w   
                          | we6wj_afzuesr1zwnl   
                          | qusz_xa0ku_toij493    
                          | jzbjl5cnc_hb5hixv   
                          | vwmbmpalhwfnoi_0g   
                          | bi0wblozr4jb8yf4    
                          ;


  wire fkdm70orcrtvcpzq7ojzw4s = mae_6a_pxmep9hv     
                         | vjw25i19dpz3    
                         | k9vvweo5_a_q_ip2l   
                         | w3njc277ysi3uz1    
                         | g8wclh3x6xlwa3ncq   
                         | go4w_xvuj1m     
                         | swvisnb87cxn83z    
                         | hp66bsfn_5mnw7gw6   
                         | szsij0guhgpj    
                         | hugyxq6gvlbt7tp   
                         | tpv9dscg_ntzh_rhh4   
                         | b0wowenfcyq_6_e  
                         | c784pnrp9fe0jg6ne39  
                         | kc_yoe3swf_o07x7p  
                         | ugiayevhrf3oqht9  
                         | higk3ii9e9i_f    
                         | g6_j6lr4ti9yu    
                         | jr97br_y15cmo2ku    
                         | k0tmdbnsotlk    
                         | hfqcy171lm219z2    
                         | tv4hqiny5afky9w   
                         | we6wj_afzuesr1zwnl   
                         | qusz_xa0ku_toij493    
                         | xnb761cg1sb1d    
                         | e02lkx_fya1ouym7h   
                         | elcvhpi2hcg0    
                         | n8r0676nkk3s04b7   
                         | m3fice1xap_p463s    
                         | et2vvn5b9hs2dsxc   
                         | q92dtkdebjot0e    
                         | dpm72l5g2io4k   
                         | lf8nodmhavxf    
                         | ta99gbty1xpqs6_ahm   
                         | blk15yrqxkt8zs2br    
                         | phiws9b8v856wgd   
                         | fj50cc2xxbpn     
                         | uavbu3i6ubzz     
                         | dsp656i_shm9fbrjf    
                         | fklgk6eyb2vd8    
                         | zfotdct2of6_kc   
                         | k1oqlvc677n04h94z31  
                         | wean5xmif_myv   
                         | qzptr55gc1d815k  
                         | fouln9y77frzodomf    
                         | ot7hpozxj594mxo0o8   
                         | q9uit_5jup8pgp6l  
                         | hked2y47eglmii   
                         | utvej5knrsiltp5b  
                         | r2icw20xk206b  
                         ;
  wire jvifik1nc718375n_1ge =                         
                           gjhl0yua7khqyyj7    
                         | n7z6su9ff17vc26hu   
                         | rp86b05b7wi0gsy7np  
                         | jt75suen_okjf02   
                         | uoy8pb4b3_q04van  
                         | esnmi_yufd7l1af    
                         | hp3zdh34mwyu_   
                         | quh0wjpu8_60_00  
                         | yyq89zr8ntwjgvv9dh   
                         | blezqucpbhjpa4v9  
                         | o5obw4mzrir4f2ofd    
                         | osn82rwdapvn3cunh   
                         | jto_jycd4wmbzar  
                         | d4roaqpdp0v1368y   
                         | owqgxd_mnoeuh58 
                         | vq0ayiqnvwy2exgn   
                         | yrp4tnx0z0vr9if  
                         | bha_2ihvu1x5vf6 
                         | rrlsg7zpsrnhfxb  
                         | krefblqj6lij3t4p 
                         | k06e5l0uw9wzwp2it   
                         | ha32lltdxd7x19  
                         | itt7e1z4g56bjpzdcq 
                         | m52a83vna7cr18mdn  
                         | c80ogd8uqs8qta9l1ev 
                         | z53vzzym9v5v6   
                         | ns6x4s_o3pi6ax2n  
                         | nb0wrp9_4ugc6qkjx7 
                         | z5bi2emm96esv_geki  
                         | jmbuhj5mdexw1m3uqq 
                         | lnchd6wpif2lsuic_  
                         | v2k3hrn_5xg64b7aocn 
                         | akr76mirt0394rwypu 
                         | mckx1mltgmxacp_ 
                         | typ6wj08ixws3lsuso 
                         | ijvh48b4xaa54zh   
                         | qawzrnnnqu9zw8   
                         | k4x3xpwe9_94trje   
                         | eytzcjin8i_o7qgg2g   
                         | ecccb2oy3kp6vbt   
                         | jzbjl5cnc_hb5hixv   
                         | vwmbmpalhwfnoi_0g   
                         | bi0wblozr4jb8yf4    
                         ;

  wire v6xqyug4ri5kzkcv8gkoa3z =                         
                           olzyli2shf6m0eu    
                         | r7cnjrtmoa4z3wzm   
                         | xs9gkwo3sk9927f  
                         | t622z2sipa9amny   
                         | gplqhxgap4qxw2585n  
                         | hd73e7ysgqar7d82    
                         | ouz2qqdkqv42w   
                         | i9k7gr9f1m5x4z9m7sw  
                         | w1064psfmbve8hpe   
                         | gisgif8kbt3puleu  
                         | rnblmzik1pew6va2h    
                         | dimrfoq94vmw2xn1t   
                         | xppjwy_axpkzto1n_hs  
                         | ev_fa6s12jdsf7   
                         | da7q3cxfn4d3s1k50 
                         | dmzs8qjfkowxd   
                         | xq79ouq18ya2qxjmwx  
                         | xm5w1y9xnpmzt7_fp2aq 
                         | elkxwjgl9ny2u6k3dg  
                         | g73i4v_qd7tqi0fc 
                         | j_jcm4qgb9x62   
                         | cf2ndyjmh3psm0oe2  
                         | pcx1a0uxtq0mr8gyc 
                         | hu6futh2tv8zrpvuhbq  
                         | r7_qpw537yx2nx2tbsj 
                         | uxzv2w6nerfya6b   
                         | ky8_zvpu3hzcuwzma  
                         | fffc565224sv9zh5bt9 
                         | q5kg_hwy37mzu95q  
                         | kv6sfx3a9qhkrx75k 
                         | nwvvvndgm3k0n   
                         | e_giw7b4ut0jmmpy9a   
                         | z79y6w0q_w4smuqg   
                         | buou043vqauc4   
                         | v_b574hro993x   
                         ;

  assign vu8cn0tjzmmmjqj_9   = 
                           fkdm70orcrtvcpzq7ojzw4s
                         | jvifik1nc718375n_1ge
                         | v6xqyug4ri5kzkcv8gkoa3z
                           ;



  
  

  
  
  
  
  
  wire w56r8eynob2o6o2f      = t61y7hkwkrvm7s & ezupw6o2yfm5ojugrc3 & gu_2fhfulrttqq4e_fiax;
  wire rr2t_274mgggv4l     = t61y7hkwkrvm7s & ezupw6o2yfm5ojugrc3 & osr23kerkrxjqbsvthv5n5 & r70hhozfmlgd3eqafzt;    
  wire ohirsq2vr6upw1     = t61y7hkwkrvm7s & ezupw6o2yfm5ojugrc3 & wambasxikyrgwdud7610fe;
  wire dd2765se3n92h_4qm    = t61y7hkwkrvm7s & ezupw6o2yfm5ojugrc3 & osr23kerkrxjqbsvthv5n5 & kis_u1bo6hhg_7rlffxs;    
  wire mvahzj2wotaon8k5      = t61y7hkwkrvm7s & ezupw6o2yfm5ojugrc3 & k3sfqtpqynzqda4xtugl4;
  wire ze2pvt1ckieqvubdc     = t61y7hkwkrvm7s & ezupw6o2yfm5ojugrc3 & g1qw0ijt6cz4o1fnmqoyhd & r70hhozfmlgd3eqafzt;    
  wire cec0fhw3i5d0d     = t61y7hkwkrvm7s & ezupw6o2yfm5ojugrc3 & bja_lg9vofv9y0s4oddhrjc;
  wire us8ffe1ajwplzv    = t61y7hkwkrvm7s & ezupw6o2yfm5ojugrc3 & g1qw0ijt6cz4o1fnmqoyhd & kis_u1bo6hhg_7rlffxs;    
  wire s5punsx6wlx69cp5      = t61y7hkwkrvm7s & ezupw6o2yfm5ojugrc3 & xxejssnpnxt8oi1caja;
  wire e0i6g36mshur     = t61y7hkwkrvm7s & ezupw6o2yfm5ojugrc3 & rywrk93gumczcc8csvqrzq & r70hhozfmlgd3eqafzt;    
  wire hi18wnm3p8d8     = t61y7hkwkrvm7s & ezupw6o2yfm5ojugrc3 & kwpxw02f_f6zyvb3it4sg4;
  wire k1t9wj3kakgh8lgi    = t61y7hkwkrvm7s & ezupw6o2yfm5ojugrc3 & rywrk93gumczcc8csvqrzq & kis_u1bo6hhg_7rlffxs;    
  wire h2g7hojc13xd1o    = t61y7hkwkrvm7s & ezupw6o2yfm5ojugrc3 & gr5b6bl6ypmzx3z57tmi;
  wire a5mk33koimh2hpws5um   = t61y7hkwkrvm7s & ezupw6o2yfm5ojugrc3 & opprr4u0rfe_9t1ilq;
  wire r4ql1yhsypyd     = t61y7hkwkrvm7s & ezupw6o2yfm5ojugrc3 & ra742uamumnh7ulbty15;
  wire wp21v56lwrh7tyhwwg    = t61y7hkwkrvm7s & ezupw6o2yfm5ojugrc3 & po6ddes535c20_mmy_2u85p & x3m205i475_nt098cv;     
  wire cheq4_h7001nganzk4    = t61y7hkwkrvm7s & ezupw6o2yfm5ojugrc3 & i3yg5uqgsrfhxxu1pt4o3;
  wire wlt11ejucxvlshgz   = t61y7hkwkrvm7s & ezupw6o2yfm5ojugrc3 & po6ddes535c20_mmy_2u85p & km4hjrsbw2uxh2_qt;     
  wire ayuau69afu1g     = t61y7hkwkrvm7s & ezupw6o2yfm5ojugrc3 & xalf55zxhxx021sqlvd9_9;
  wire nb683t6oih_ek14    = t61y7hkwkrvm7s & ezupw6o2yfm5ojugrc3 & hfkmqai7ufo0_uc36i & x3m205i475_nt098cv;     
  wire frhfg7rk6sjyfnw5z3    = t61y7hkwkrvm7s & ezupw6o2yfm5ojugrc3 & bwbrcnczkn_1flyk41tn5q8;
  wire y5khcw8jpof6ude5   = t61y7hkwkrvm7s & ezupw6o2yfm5ojugrc3 & hfkmqai7ufo0_uc36i & km4hjrsbw2uxh2_qt;     
  wire kpp0vn2f3g0x     = t61y7hkwkrvm7s & ezupw6o2yfm5ojugrc3 & mw5b0jbgrdfc4zozpy333k;
  wire cuf6ntg4j_lumj4pox    = t61y7hkwkrvm7s & ezupw6o2yfm5ojugrc3 & i_npu8b57pt8jq9y8wi6 & x3m205i475_nt098cv;     
  wire f4rqm494l0jjw7use    = t61y7hkwkrvm7s & ezupw6o2yfm5ojugrc3 & ot56pcza1qpiqzjwuib4ioq;
  wire yy2boizah9n6vll94z   = t61y7hkwkrvm7s & ezupw6o2yfm5ojugrc3 & i_npu8b57pt8jq9y8wi6 & km4hjrsbw2uxh2_qt;     
  wire y10yq62t_2h9f_i_d1   = t61y7hkwkrvm7s & ezupw6o2yfm5ojugrc3 & ew4asffkh_z5lao1cnzk9g;
  wire qbj_bpx859fqfk9sd  = t61y7hkwkrvm7s & ezupw6o2yfm5ojugrc3 & q4yuw6wl9o929gj8k2ovt;
  wire yny8lgx5s6i7mpr     = t61y7hkwkrvm7s & t8jc64yc1l6q8eclq_c & ra742uamumnh7ulbty15;
  wire l1zwxuvb407cnts    = t61y7hkwkrvm7s & t8jc64yc1l6q8eclq_c & po6ddes535c20_mmy_2u85p;     
  wire tnkhbxhqbrvp13vu    = t61y7hkwkrvm7s & t8jc64yc1l6q8eclq_c & i3yg5uqgsrfhxxu1pt4o3;
  wire ivse5_zisiibgf8oum   = t61y7hkwkrvm7s & t8jc64yc1l6q8eclq_c & xx5u6vajn90lcpxcfi_d26;     
  wire ig66294d77dyx_izt     = t61y7hkwkrvm7s & t8jc64yc1l6q8eclq_c & xalf55zxhxx021sqlvd9_9;
  wire oizf0jkb_iwlm68mrw    = t61y7hkwkrvm7s & t8jc64yc1l6q8eclq_c & hfkmqai7ufo0_uc36i;     
  wire uf77s2stj_9j6ex    = t61y7hkwkrvm7s & t8jc64yc1l6q8eclq_c & bwbrcnczkn_1flyk41tn5q8;
  wire wyit9nrrvctc4ii9rb   = t61y7hkwkrvm7s & t8jc64yc1l6q8eclq_c & oezo_lnpso_pe9xd5gp;     
  wire vlgbdo21_xc2k     = t61y7hkwkrvm7s & t8jc64yc1l6q8eclq_c & mw5b0jbgrdfc4zozpy333k;
  wire dqmsf6gtvzuqhis21l    = t61y7hkwkrvm7s & t8jc64yc1l6q8eclq_c & i_npu8b57pt8jq9y8wi6;     
  wire dvn60wqlpj1v67en3    = t61y7hkwkrvm7s & t8jc64yc1l6q8eclq_c & ot56pcza1qpiqzjwuib4ioq;
  wire i6q7_tpl_4f61n   = t61y7hkwkrvm7s & t8jc64yc1l6q8eclq_c & pq_m0zj_hjvfii9out1;     
  wire samkfqmeumr_fpwz43   = t61y7hkwkrvm7s & t8jc64yc1l6q8eclq_c & ew4asffkh_z5lao1cnzk9g;
  wire hdf0loxgf2t36h7izpqs  = t61y7hkwkrvm7s & t8jc64yc1l6q8eclq_c & q4yuw6wl9o929gj8k2ovt;
  wire vz7mnovu_m51dq1    = t61y7hkwkrvm7s & d24iqtxvb2trplxk2m & x_c94bnppi8ngabfz2iw;  
  wire jr9hao6bk8d      = t61y7hkwkrvm7s & d24iqtxvb2trplxk2m & lipdgvrqr439y_cnsv;
  wire jicp1hi2zypaj     = t61y7hkwkrvm7s & d24iqtxvb2trplxk2m & e9kyqn6z0nnxcqwggfu2c;                      
  wire wtsb9emi6nj0dzl_0b    = t61y7hkwkrvm7s & d24iqtxvb2trplxk2m & opprr4u0rfe_9t1ilq;
  wire mishqln22ifbrftv47c   = t61y7hkwkrvm7s & d24iqtxvb2trplxk2m & qr23_2sadkfk2963qo;
  wire uya11_4faw_3bxv5     = t61y7hkwkrvm7s & d24iqtxvb2trplxk2m & veb9c0lxewgh_4qiy5;
  wire rkx2z9tuldgd39zp    = t61y7hkwkrvm7s & d24iqtxvb2trplxk2m & fr9vuzzy67toa8_rpz_;
  
  wire s_6vyiuywqqrd9say   = 1'b0;
  wire k7c8gfhghnfklxr2  = 1'b0;


  

  
  wire [62-1:0] ykn2abyw7s2voefu;
  assign ykn2abyw7s2voefu[3:0]           = 4'd13;
  assign ykn2abyw7s2voefu[4:4]          = vlfahv69;
  assign ykn2abyw7s2voefu[10:5      ] = pq5pe3yehrqxr[25:20];
  assign ykn2abyw7s2voefu[11:11     ] = w56r8eynob2o6o2f    ; 
  assign ykn2abyw7s2voefu[12:12    ] = rr2t_274mgggv4l   ;
  assign ykn2abyw7s2voefu[13:13    ] = ohirsq2vr6upw1   ;
  assign ykn2abyw7s2voefu[14:14   ] = dd2765se3n92h_4qm  ;
  assign ykn2abyw7s2voefu[15:15     ] = mvahzj2wotaon8k5    ;
  assign ykn2abyw7s2voefu[16:16    ] = ze2pvt1ckieqvubdc   ;
  assign ykn2abyw7s2voefu[17:17    ] = cec0fhw3i5d0d   ;
  assign ykn2abyw7s2voefu[18:18   ] = us8ffe1ajwplzv  ;
  assign ykn2abyw7s2voefu[19:19     ] = s5punsx6wlx69cp5    ;
  assign ykn2abyw7s2voefu[20:20    ] = e0i6g36mshur   ;
  assign ykn2abyw7s2voefu[21:21    ] = hi18wnm3p8d8   ;
  assign ykn2abyw7s2voefu[22:22   ] = k1t9wj3kakgh8lgi  ;
  assign ykn2abyw7s2voefu[23:23   ] = h2g7hojc13xd1o  ;
  assign ykn2abyw7s2voefu[25:25  ] = a5mk33koimh2hpws5um ;
  assign ykn2abyw7s2voefu[26:26    ] = r4ql1yhsypyd   ;
  assign ykn2abyw7s2voefu[27:27   ] = wp21v56lwrh7tyhwwg  ;
  assign ykn2abyw7s2voefu[28:28   ] = cheq4_h7001nganzk4  ;
  assign ykn2abyw7s2voefu[29:29  ] = wlt11ejucxvlshgz ;
  assign ykn2abyw7s2voefu[30:30    ] = ayuau69afu1g   ;
  assign ykn2abyw7s2voefu[31:31   ] = nb683t6oih_ek14  ;
  assign ykn2abyw7s2voefu[32:32   ] = frhfg7rk6sjyfnw5z3  ;
  assign ykn2abyw7s2voefu[33:33  ] = y5khcw8jpof6ude5 ;
  assign ykn2abyw7s2voefu[34:34   ] = kpp0vn2f3g0x   ;
  assign ykn2abyw7s2voefu[35:35  ] = cuf6ntg4j_lumj4pox  ;
  assign ykn2abyw7s2voefu[36:36   ] = f4rqm494l0jjw7use  ;
  assign ykn2abyw7s2voefu[37:37  ] = yy2boizah9n6vll94z ;
  assign ykn2abyw7s2voefu[38:38  ] = y10yq62t_2h9f_i_d1 ;
  assign ykn2abyw7s2voefu[40:40 ] = qbj_bpx859fqfk9sd;
  assign ykn2abyw7s2voefu[41:41     ] = jr9hao6bk8d    ;
  assign ykn2abyw7s2voefu[42:42    ] = jicp1hi2zypaj   ;
  assign ykn2abyw7s2voefu[43:43   ] = wtsb9emi6nj0dzl_0b  ;
  assign ykn2abyw7s2voefu[44:44  ] = mishqln22ifbrftv47c ;
  assign ykn2abyw7s2voefu[45:45    ] = uya11_4faw_3bxv5   ;
  assign ykn2abyw7s2voefu[46:46   ] = rkx2z9tuldgd39zp  ;
  assign ykn2abyw7s2voefu[39 ] = k7c8gfhghnfklxr2 ;
  assign ykn2abyw7s2voefu[24  ] = s_6vyiuywqqrd9say  ;
  assign ykn2abyw7s2voefu[47:47    ] = yny8lgx5s6i7mpr   ;   
  assign ykn2abyw7s2voefu[48:48   ] = l1zwxuvb407cnts  ;   
  assign ykn2abyw7s2voefu[49:49   ] = tnkhbxhqbrvp13vu  ;   
  assign ykn2abyw7s2voefu[50:50  ] = ivse5_zisiibgf8oum ;   
  assign ykn2abyw7s2voefu[51:51    ] = ig66294d77dyx_izt   ;   
  assign ykn2abyw7s2voefu[52:52   ] = oizf0jkb_iwlm68mrw  ;   
  assign ykn2abyw7s2voefu[53:53   ] = uf77s2stj_9j6ex  ;   
  assign ykn2abyw7s2voefu[54:54  ] = wyit9nrrvctc4ii9rb ;   
  assign ykn2abyw7s2voefu[55:55    ] = vlgbdo21_xc2k   ;   
  assign ykn2abyw7s2voefu[56:56   ] = dqmsf6gtvzuqhis21l  ;   
  assign ykn2abyw7s2voefu[57:57   ] = dvn60wqlpj1v67en3  ;   
  assign ykn2abyw7s2voefu[58:58  ] = i6q7_tpl_4f61n ;   
  assign ykn2abyw7s2voefu[59:59  ] = samkfqmeumr_fpwz43 ;   
  assign ykn2abyw7s2voefu[60:60 ] = hdf0loxgf2t36h7izpqs;   
  assign ykn2abyw7s2voefu[61:61   ] = vz7mnovu_m51dq1  ;   

  
  wire yg_3i0cfu6iwmj = 
                      | w56r8eynob2o6o2f    
                      | rr2t_274mgggv4l   
                      | ohirsq2vr6upw1   
                      | dd2765se3n92h_4qm  
                      | mvahzj2wotaon8k5    
                      | ze2pvt1ckieqvubdc   
                      | cec0fhw3i5d0d   
                      | us8ffe1ajwplzv  
                      | s5punsx6wlx69cp5    
                      | e0i6g36mshur   
                      | hi18wnm3p8d8   
                      | k1t9wj3kakgh8lgi  
                      | h2g7hojc13xd1o  
                      | a5mk33koimh2hpws5um 
                      | r4ql1yhsypyd   
                      | wp21v56lwrh7tyhwwg  
                      | cheq4_h7001nganzk4  
                      | wlt11ejucxvlshgz 
                      | ayuau69afu1g   
                      | nb683t6oih_ek14  
                      | frhfg7rk6sjyfnw5z3  
                      | y5khcw8jpof6ude5 
                      | kpp0vn2f3g0x   
                      | cuf6ntg4j_lumj4pox  
                      | f4rqm494l0jjw7use  
                      | yy2boizah9n6vll94z 
                      | y10yq62t_2h9f_i_d1 
                      | qbj_bpx859fqfk9sd
                      | yny8lgx5s6i7mpr   
                      | l1zwxuvb407cnts  
                      | tnkhbxhqbrvp13vu  
                      | ivse5_zisiibgf8oum 
                      | ig66294d77dyx_izt   
                      | oizf0jkb_iwlm68mrw  
                      | uf77s2stj_9j6ex  
                      | wyit9nrrvctc4ii9rb 
                      | vlgbdo21_xc2k   
                      | dqmsf6gtvzuqhis21l  
                      | dvn60wqlpj1v67en3  
                      | i6q7_tpl_4f61n 
                      | samkfqmeumr_fpwz43 
                      | hdf0loxgf2t36h7izpqs
                      | vz7mnovu_m51dq1
                      | jr9hao6bk8d    
                      | jicp1hi2zypaj   
                      | wtsb9emi6nj0dzl_0b  
                      | mishqln22ifbrftv47c 
                      | uya11_4faw_3bxv5   
                      | rkx2z9tuldgd39zp  
                      | s_6vyiuywqqrd9say  
                      | k7c8gfhghnfklxr2  
                      ;
                      
  
  wire podz_mnetypiu7    = t61y7hkwkrvm7s & ezupw6o2yfm5ojugrc3 & t33zd67g1c1fzxs_g27e34r & r70hhozfmlgd3eqafzt;    
  wire fkaztmo9sputf    = t61y7hkwkrvm7s & ezupw6o2yfm5ojugrc3 & t33zd67g1c1fzxs_g27e34r & cgtj86qjqc4whb8p2jo;    
  wire dl4pq4785d2evg   = t61y7hkwkrvm7s & ezupw6o2yfm5ojugrc3 & pq_m0zj_hjvfii9out1 & x3m205i475_nt098cv;     
  wire a90cuq3gcnfvujvq4t   = t61y7hkwkrvm7s & ezupw6o2yfm5ojugrc3 & pq_m0zj_hjvfii9out1 & km4hjrsbw2uxh2_qt;     
  wire a7bnvi_up37cgwlgo   = t61y7hkwkrvm7s & ezupw6o2yfm5ojugrc3 & brnnngwkv59w2kz9usv3k8;						
  wire p0wx5tkzaf886os   = t61y7hkwkrvm7s & ezupw6o2yfm5ojugrc3 & sketktuyfh2vxjbshrr;
  wire qe8meo02o4s562hq = t61y7hkwkrvm7s & ezupw6o2yfm5ojugrc3 & styktg7w7fi36jw0e5n4h93 & asvcpbvzr7u9gfqr_hlh68; 
  wire yxwrh57b5d5hqw19s7waz = t61y7hkwkrvm7s & ezupw6o2yfm5ojugrc3 & styktg7w7fi36jw0e5n4h93 & kre86u005m4jj77idkd170; 
  wire pos61lm9pwmw50y3ycsi = t61y7hkwkrvm7s & ezupw6o2yfm5ojugrc3 & styktg7w7fi36jw0e5n4h93 & h6jjzsxi8aw0us788h; 
  wire p27yz0zu7tm7s9fjd6r = t61y7hkwkrvm7s & ezupw6o2yfm5ojugrc3 & styktg7w7fi36jw0e5n4h93 & yswws2ff7bkbvaic3it7g; 
  wire yflkcdpfbgtf0_au_ = t61y7hkwkrvm7s & ezupw6o2yfm5ojugrc3 & styktg7w7fi36jw0e5n4h93 & yc8o21itzjuxfoo_32; 
  wire q7enr9cewlaqzs11e = t61y7hkwkrvm7s & ezupw6o2yfm5ojugrc3 & styktg7w7fi36jw0e5n4h93 & z1_re9ax86eago99v6ic1ke; 
  wire w2ht8y0gz2gav1oxv_x = t61y7hkwkrvm7s & ezupw6o2yfm5ojugrc3 & styktg7w7fi36jw0e5n4h93 & yiprb7xpgx9hgyddnxoh; 
  wire k_dh889fnsknt8gtnr = t61y7hkwkrvm7s & ezupw6o2yfm5ojugrc3 & styktg7w7fi36jw0e5n4h93 & hutky_0znezwi4oz7cs; 
  wire p9ke7v3lz3w4tjmp7 = t61y7hkwkrvm7s & ezupw6o2yfm5ojugrc3 & styktg7w7fi36jw0e5n4h93 & fe7237ktiiy1d5p48dam8; 
  wire xe7xs7at6t0eaa288 = t61y7hkwkrvm7s & ezupw6o2yfm5ojugrc3 & styktg7w7fi36jw0e5n4h93 & f9jz4kxv632mfmwjuwinhm; 
  wire ai0h133sxmklw2sh  = t61y7hkwkrvm7s & d24iqtxvb2trplxk2m & jhbiy5xf0ygws7apfg03;
  wire z2wowpcfaid11_i2  = t61y7hkwkrvm7s & d24iqtxvb2trplxk2m & b12f43e4j_bhgigw_xvwmqe;
  wire h53qoytt_1mtyfcas464  = t61y7hkwkrvm7s & d24iqtxvb2trplxk2m & ha7x94wp2o8bpzvtiq_d;
  wire uhcjsl31yez759e  = t61y7hkwkrvm7s & d24iqtxvb2trplxk2m & i_nd_auanr4nliiv9ru_mjy;
  wire ey6lu8os16zzfpjn  = t61y7hkwkrvm7s & t8jc64yc1l6q8eclq_c & jhbiy5xf0ygws7apfg03;
  wire zjlc5cdmk3h_py1d37_o  = t61y7hkwkrvm7s & t8jc64yc1l6q8eclq_c & b12f43e4j_bhgigw_xvwmqe;
  wire wkjozhj8gkzn17m  = t61y7hkwkrvm7s & t8jc64yc1l6q8eclq_c & ha7x94wp2o8bpzvtiq_d;
  wire hbc1edn1_8f285is51x  = t61y7hkwkrvm7s & t8jc64yc1l6q8eclq_c & i_nd_auanr4nliiv9ru_mjy;
  wire rf_x1axtwqsgz14s    = t61y7hkwkrvm7s & dwe8qnpoudm94xa & lipdgvrqr439y_cnsv & qgge30ma6bacftkfuwr;
  wire h193fufzl9k9j8_bi    = t61y7hkwkrvm7s & dwe8qnpoudm94xa & lipdgvrqr439y_cnsv & tv_mqy2vnetyki2mitz;
  wire vhzlyir7ae3m3dx_o    = t61y7hkwkrvm7s & dwe8qnpoudm94xa & lipdgvrqr439y_cnsv & iqlkuiiuioeb0zx_mespm;
  wire brwqtymgz1q318trw    = t61y7hkwkrvm7s & dwe8qnpoudm94xa & lipdgvrqr439y_cnsv & b2rqyt08n40btyec123;
  wire g3eepk0cdmakl1u    = t61y7hkwkrvm7s & dwe8qnpoudm94xa & lipdgvrqr439y_cnsv & nielo5a2gnsny_mbq2;
  wire nybn83l8h8rmm5tk    = t61y7hkwkrvm7s & dwe8qnpoudm94xa & lipdgvrqr439y_cnsv & pnz7nx6huw6bc2xirgh;
  wire ss1_hx3eo4rnxdbn6    = t61y7hkwkrvm7s & dwe8qnpoudm94xa & lipdgvrqr439y_cnsv & u1y9fqpjmgbvqp01zyup348;
  wire i679vkh0e1766qyk    = t61y7hkwkrvm7s & dwe8qnpoudm94xa & lipdgvrqr439y_cnsv & mv0ortg5fw6xo5qko1gvm4;
  wire yjv8gea4klbna3j3p     = t61y7hkwkrvm7s & ezupw6o2yfm5ojugrc3 & tfcuen58mdto351cstsry5 & qgge30ma6bacftkfuwr; 
  wire kqdvzyoypaurb      = t61y7hkwkrvm7s & ezupw6o2yfm5ojugrc3 & tfcuen58mdto351cstsry5 & tv_mqy2vnetyki2mitz; 
  wire slq7c7rnln8nm776      = t61y7hkwkrvm7s & ezupw6o2yfm5ojugrc3 & tfcuen58mdto351cstsry5 & b2rqyt08n40btyec123; 
  wire wwcr_z51mt1s8b13e    = t61y7hkwkrvm7s & ezupw6o2yfm5ojugrc3 & tfcuen58mdto351cstsry5 & asvcpbvzr7u9gfqr_hlh68; 
  wire xehsykkcziznmy0     = t61y7hkwkrvm7s & ezupw6o2yfm5ojugrc3 & tfcuen58mdto351cstsry5 & kre86u005m4jj77idkd170; 
  wire o1bf95sjlu96k0md     = t61y7hkwkrvm7s & ezupw6o2yfm5ojugrc3 & tfcuen58mdto351cstsry5 & yswws2ff7bkbvaic3it7g; 
  wire h10rn5j_pjeeh_gi    = t61y7hkwkrvm7s & ezupw6o2yfm5ojugrc3 & tfcuen58mdto351cstsry5 & qgai63fi1e6hqmwnsi7t; 
  wire u41dwwpt95uk     = t61y7hkwkrvm7s & ezupw6o2yfm5ojugrc3 & tfcuen58mdto351cstsry5 & yzqtbppdh3mlkyfzf0g6at; 
  wire xen0hyummyuh     = t61y7hkwkrvm7s & ezupw6o2yfm5ojugrc3 & tfcuen58mdto351cstsry5 & nf2wc7g6poblu9r9_r; 
  wire vkh3wnxoirfr15dtj    = t61y7hkwkrvm7s & ezupw6o2yfm5ojugrc3 & wp2e1icm345eqoi7xse0mo;
  wire lhx06f20_s0toyo1q7   = t61y7hkwkrvm7s & ezupw6o2yfm5ojugrc3 & i37i_iou1kvjw2svv8;                      
  wire o0rfcptm6iob1mej      = t61y7hkwkrvm7s & ezupw6o2yfm5ojugrc3 & ny5cwervdr0wq805l6q;
  wire z3kk91ocqzu25     = t61y7hkwkrvm7s & ezupw6o2yfm5ojugrc3 & cbgxogbpgug3v8_faeo3;
  wire tx04m_rvbl9sow     = t61y7hkwkrvm7s & w__ro7gwx6w331 & x99kg2smyvi6ahhq46x;
  wire r5qet1mocbtcig      = t61y7hkwkrvm7s & ezupw6o2yfm5ojugrc3 & styktg7w7fi36jw0e5n4h93 & r70hhozfmlgd3eqafzt;    
  wire y_pnmfuono692     = t61y7hkwkrvm7s & ezupw6o2yfm5ojugrc3 & styktg7w7fi36jw0e5n4h93 & qgai63fi1e6hqmwnsi7t; 
  wire x5p2cakvpfx79bot    = t61y7hkwkrvm7s & ezupw6o2yfm5ojugrc3 & styktg7w7fi36jw0e5n4h93 & yzqtbppdh3mlkyfzf0g6at; 

  wire y_0id5h2cb8ukkao;

  
  wire [60-1:0] p8svuggnu7zvtlojt;
  assign p8svuggnu7zvtlojt[3:0]           = 4'd12;
  assign p8svuggnu7zvtlojt[4:4]          = vlfahv69;
  assign p8svuggnu7zvtlojt[10:5      ] = pq5pe3yehrqxr[24:20];
  assign p8svuggnu7zvtlojt[11:11   ] = podz_mnetypiu7   ; 
  assign p8svuggnu7zvtlojt[12:12   ] = fkaztmo9sputf   ; 
  assign p8svuggnu7zvtlojt[13:13  ] = dl4pq4785d2evg  ;
  assign p8svuggnu7zvtlojt[14:14  ] = a90cuq3gcnfvujvq4t  ;
  assign p8svuggnu7zvtlojt[15:15  ] = a7bnvi_up37cgwlgo  ;
  assign p8svuggnu7zvtlojt[16:16  ] = p0wx5tkzaf886os  ;
  assign p8svuggnu7zvtlojt[17:17] = qe8meo02o4s562hq;
  assign p8svuggnu7zvtlojt[18:18] = yxwrh57b5d5hqw19s7waz;
  assign p8svuggnu7zvtlojt[19:19] = pos61lm9pwmw50y3ycsi;
  assign p8svuggnu7zvtlojt[20:20] = p27yz0zu7tm7s9fjd6r;
  assign p8svuggnu7zvtlojt[21:21] = yflkcdpfbgtf0_au_;
  assign p8svuggnu7zvtlojt[22:22] = q7enr9cewlaqzs11e;
  assign p8svuggnu7zvtlojt[23:23] = w2ht8y0gz2gav1oxv_x;
  assign p8svuggnu7zvtlojt[24:24] = k_dh889fnsknt8gtnr;
  assign p8svuggnu7zvtlojt[25:25] = p9ke7v3lz3w4tjmp7;
  assign p8svuggnu7zvtlojt[26:26] = xe7xs7at6t0eaa288;
  assign p8svuggnu7zvtlojt[27:27   ] = ai0h133sxmklw2sh ;
  assign p8svuggnu7zvtlojt[28:28   ] = z2wowpcfaid11_i2 ;
  assign p8svuggnu7zvtlojt[29:29   ] = h53qoytt_1mtyfcas464 ;
  assign p8svuggnu7zvtlojt[30:30   ] = uhcjsl31yez759e ;
  assign p8svuggnu7zvtlojt[56:56   ] = ey6lu8os16zzfpjn ;
  assign p8svuggnu7zvtlojt[57:57   ] = zjlc5cdmk3h_py1d37_o ;
  assign p8svuggnu7zvtlojt[58:58   ] = wkjozhj8gkzn17m ;
  assign p8svuggnu7zvtlojt[59:59   ] = hbc1edn1_8f285is51x ;
  assign p8svuggnu7zvtlojt[31   ] = rf_x1axtwqsgz14s   ;
  assign p8svuggnu7zvtlojt[32   ] = h193fufzl9k9j8_bi   ;
  assign p8svuggnu7zvtlojt[33   ] = vhzlyir7ae3m3dx_o   ;
  assign p8svuggnu7zvtlojt[34   ] = brwqtymgz1q318trw   ;
  assign p8svuggnu7zvtlojt[35   ] = g3eepk0cdmakl1u   ;
  assign p8svuggnu7zvtlojt[36   ] = nybn83l8h8rmm5tk   ;
  assign p8svuggnu7zvtlojt[37   ] = ss1_hx3eo4rnxdbn6   ;
  assign p8svuggnu7zvtlojt[38   ] = i679vkh0e1766qyk   ;
  assign p8svuggnu7zvtlojt[39:39    ] = yjv8gea4klbna3j3p    ; 
  assign p8svuggnu7zvtlojt[40:40     ] = kqdvzyoypaurb     ; 
  assign p8svuggnu7zvtlojt[41:41     ] = slq7c7rnln8nm776     ; 
  assign p8svuggnu7zvtlojt[42:42   ] = wwcr_z51mt1s8b13e   ; 
  assign p8svuggnu7zvtlojt[43:43    ] = xehsykkcziznmy0    ; 
  assign p8svuggnu7zvtlojt[44:44    ] = o1bf95sjlu96k0md    ; 
  assign p8svuggnu7zvtlojt[45:45   ] = h10rn5j_pjeeh_gi   ; 
  assign p8svuggnu7zvtlojt[46:46    ] = u41dwwpt95uk    ; 
  assign p8svuggnu7zvtlojt[47:47    ] = xen0hyummyuh    ; 
  assign p8svuggnu7zvtlojt[48:48   ] = vkh3wnxoirfr15dtj   ; 
  assign p8svuggnu7zvtlojt[49:49  ] = lhx06f20_s0toyo1q7  ; 
  assign p8svuggnu7zvtlojt[50:50     ] = o0rfcptm6iob1mej     ; 
  assign p8svuggnu7zvtlojt[51:51    ] = z3kk91ocqzu25    ; 
  assign p8svuggnu7zvtlojt[52:52    ] = tx04m_rvbl9sow    ; 
  assign p8svuggnu7zvtlojt[53:53     ] = r5qet1mocbtcig     ; 
  assign p8svuggnu7zvtlojt[54:54    ] = y_pnmfuono692    ; 
  assign p8svuggnu7zvtlojt[55:55   ] = x5p2cakvpfx79bot   ; 

  
  assign y_0id5h2cb8ukkao = 
                       | podz_mnetypiu7
                       | fkaztmo9sputf   
                       | dl4pq4785d2evg  
                       | a90cuq3gcnfvujvq4t  
                       | a7bnvi_up37cgwlgo  
                       | p0wx5tkzaf886os  
                       | qe8meo02o4s562hq
                       | yxwrh57b5d5hqw19s7waz
                       | pos61lm9pwmw50y3ycsi
                       | p27yz0zu7tm7s9fjd6r
                       | yflkcdpfbgtf0_au_
                       | q7enr9cewlaqzs11e
                       | w2ht8y0gz2gav1oxv_x
                       | k_dh889fnsknt8gtnr
                       | p9ke7v3lz3w4tjmp7
                       | xe7xs7at6t0eaa288
                       | ai0h133sxmklw2sh 
                       | z2wowpcfaid11_i2 
                       | h53qoytt_1mtyfcas464 
                       | uhcjsl31yez759e 
                       | ey6lu8os16zzfpjn 
                       | zjlc5cdmk3h_py1d37_o 
                       | wkjozhj8gkzn17m 
                       | hbc1edn1_8f285is51x 
                       | rf_x1axtwqsgz14s
                       | h193fufzl9k9j8_bi
                       | vhzlyir7ae3m3dx_o
                       | brwqtymgz1q318trw
                       | g3eepk0cdmakl1u
                       | nybn83l8h8rmm5tk
                       | ss1_hx3eo4rnxdbn6
                       | i679vkh0e1766qyk
                       | yjv8gea4klbna3j3p    
                       | kqdvzyoypaurb     
                       | slq7c7rnln8nm776     
                       | wwcr_z51mt1s8b13e   
                       | xehsykkcziznmy0    
                       | o1bf95sjlu96k0md    
                       | h10rn5j_pjeeh_gi   
                       | u41dwwpt95uk    
                       | xen0hyummyuh    
                       | vkh3wnxoirfr15dtj   
                       | lhx06f20_s0toyo1q7  
                       | o0rfcptm6iob1mej     
                       | z3kk91ocqzu25    
                       | tx04m_rvbl9sow    
                       | r5qet1mocbtcig     
                       | y_pnmfuono692    
                       | x5p2cakvpfx79bot   
                       ;
                        
  assign  mg4yq4mui7ruja[0]              = gdebc5b6o6bv57ax1bw; 
  assign  mg4yq4mui7ruja[1]       = yunpydbojvbs7t1vv3n9ir;
  assign  mg4yq4mui7ruja[2]      = wewa0sb6nm_e_8n25xoi;
  assign  mg4yq4mui7ruja[3]      = f_l92j9mkhdmknnhn2;
  assign  mg4yq4mui7ruja[4]     = woiza4felzgpik5ue3hx8;
  assign  mg4yq4mui7ruja[5]       = rh93dqz7x7e76_rwvdq_gv;
  assign  mg4yq4mui7ruja[6]      = dwf3ct8epliykbwg6fpvn1d;
  assign  mg4yq4mui7ruja[7]      = syyd9204a47y6qq9cyxvn7s;
  assign  mg4yq4mui7ruja[8]   = x4zc788yz37xi4o6fcfpux;
  
  assign  mg4yq4mui7ruja[9]        = ucwkku1t4g36u3iukgb ;
  assign  mg4yq4mui7ruja[10]        = avjo592wbov8cr5i ;
  assign  mg4yq4mui7ruja[11]         = kp1fyknoq74q3vs ;
  assign  mg4yq4mui7ruja[13]   = n4dlb4x1wzqqyr98jl7v8t_apmfb; 
  assign  mg4yq4mui7ruja[14]               = hxv8akm9tnbagx;
  assign  mg4yq4mui7ruja[15]             = qhmdzlcppcq8;
  assign  mg4yq4mui7ruja[17]            = vu8cn0tjzmmmjqj_9 ;
  assign  mg4yq4mui7ruja[18]       = fkdm70orcrtvcpzq7ojzw4s ;
  assign  mg4yq4mui7ruja[19]       = jvifik1nc718375n_1ge ;
  assign  mg4yq4mui7ruja[20]       = v6xqyug4ri5kzkcv8gkoa3z ;
  assign  mg4yq4mui7ruja[21]           = qm17qduoi54r_53z; 
  assign  mg4yq4mui7ruja[22]              = y_0id5h2cb8ukkao;
  assign  mg4yq4mui7ruja[23]             = yg_3i0cfu6iwmj;
  assign  mg4yq4mui7ruja[24]    = ccb88tt72pm4kk3aiztl_;
  assign  mg4yq4mui7ruja[25] = upbbycb5makv3xss7d_ueoxns88bj;
  assign  mg4yq4mui7ruja[26]               = isxv0tqhyam;
  assign  mg4yq4mui7ruja[27]  =  niiot38ff0zsxxncd0u_5fljm__dl;
  assign  mg4yq4mui7ruja[29]  = pm3poaltg6mtmffm_87yhorfj9eort_;
  assign  mg4yq4mui7ruja[28]   = hf3_u19xhtm47jygm346ih5592f;
  assign  mg4yq4mui7ruja[30] = y1fgyae1uzj7ujuxqi3znyfnbb19hjsl;                             
  assign  mg4yq4mui7ruja[31] = sfwi4o77fiwv1s1kb4mmixcewjetb_1;                             
  assign  mg4yq4mui7ruja[32] = oboq9ew68wxfv1zbbzbw6ovxumvp4ms;                             
  assign  mg4yq4mui7ruja[33] = ozipqe_4brzi2opcs5pi232jtqiu7_m6kuv;                             
  assign  mg4yq4mui7ruja[34] = imwjfayr9ztr86owxp26dtq0onjtd6dp;                             
  assign  mg4yq4mui7ruja[35] = n38usa0n35mgmntamkuxh2l5pd2gcwghz;                             
  assign  mg4yq4mui7ruja[36] = gm3156cuu5w0z0iabqd970k351i652n1u;                             
  assign  mg4yq4mui7ruja[37] = n93vkxau7xxglljhnhsxg_4jddx13kcy;                             
  assign  mg4yq4mui7ruja[38] = t88i3logg39o9_7fi_4qgfve8slrofj4j;                             
  assign  mg4yq4mui7ruja[39] = e7ilxivhp9g8urh1klgvakcpqfmwjd5tw;                             
  assign  mg4yq4mui7ruja[40] = hhf5vk7i4v5m5s0diu0q2m6pmxzvm7zeyiv7r;
  assign  mg4yq4mui7ruja[41] = e9gctcgx_15frdmbcrevvtf_2lldmasrmr9gp;
  assign  mg4yq4mui7ruja[42] = wj4suc8dinc_9d5409y_to9toxtea5b3afqoc;
  assign  mg4yq4mui7ruja[43] = o44zcer7fjl2e666o3w3zxacak78idnwavnn;
  assign  mg4yq4mui7ruja[44] = iue4b0u82l97gr25u35a4wkzrr64s8kyxgwm;
  assign  mg4yq4mui7ruja[45] = mr9h2nuumis0_vx1kbbu849xvlx89du725kw;
  assign  mg4yq4mui7ruja[46] = k0ly3yt_k96klqrmoe2jg2fjd6qz2edc5j87l;
  assign  mg4yq4mui7ruja[47] = tivrapwmioo0momgw9hmmlzhrcqyoa8a6wdu2yh;
  assign  mg4yq4mui7ruja[48] = s89z9cptleb2csl1iyj0lg_altgx5k1f6316m1h;
  assign  mg4yq4mui7ruja[49] = oy_6emad9374dtcw5eu89i4o6o5kuiqu26hsgcb;

  
  wire [5-1:0] fd7uuv9az = pq5pe3yehrqxr[31:27];
  
  
  

  assign sibtd2rf5j = t61y7hkwkrvm7s & (vu8cn0tjzmmmjqj_9 | hxv8akm9tnbagx | qhmdzlcppcq8 | y_0id5h2cb8ukkao | yg_3i0cfu6iwmj);
  wire [105-1:0] j2ba3puzp5g9g2fyuo_r3jt82 = {{105-54{1'b0}},wazt073vrvkujb_lpjze6};
  wire [105-1:0] wnflxr48uo4mtm0jalawrfbgut22h = {{105-48{1'b0}},azvwipii1valwcdp80j3_oq};
  wire [105-1:0] h159feqp7mwlb45l1mo2gff4v = {{105-40{1'b0}},no56h0p6kag9edi57joc3m};
  wire [105-1:0] olbxw0wv5dgys5s24i         = {{105-23{1'b0}},  nhqiwwnz4lmleg};
  wire [105-1:0] wtk72spw50t5zncbo1e5       = w98a0gvni829u3;
  wire [105-1:0] v9_h5km97s6fu3_in3n_p       = {{105-62{1'b0}},ykn2abyw7s2voefu};
  wire [105-1:0] jq4qgha4ovygunv2unau        = {{105-60{1'b0}}, p8svuggnu7zvtlojt};
  assign z8t7w6zr5woh649 = 
                       ({105{fkdm70orcrtvcpzq7ojzw4s}} & j2ba3puzp5g9g2fyuo_r3jt82)
                      |({105{jvifik1nc718375n_1ge}} & wnflxr48uo4mtm0jalawrfbgut22h)
                      |({105{v6xqyug4ri5kzkcv8gkoa3z}} & h159feqp7mwlb45l1mo2gff4v)
                      |({105{hxv8akm9tnbagx}}         & olbxw0wv5dgys5s24i)
                      |({105{qhmdzlcppcq8}}       & wtk72spw50t5zncbo1e5)
                      |({105{yg_3i0cfu6iwmj}}       & v9_h5km97s6fu3_in3n_p)
                      |({105{y_0id5h2cb8ukkao}}        & jq4qgha4ovygunv2unau)
                      ;

  wire eshy3jgtzqwpnq = 
      
                        (rr2t_274mgggv4l | dd2765se3n92h_4qm)        |    
                        (ze2pvt1ckieqvubdc | us8ffe1ajwplzv)        |    
                        e0i6g36mshur       |                       
                        k1t9wj3kakgh8lgi      |                       
                        wp21v56lwrh7tyhwwg      |                       
                        wlt11ejucxvlshgz     |                       
                        (nb683t6oih_ek14 | y5khcw8jpof6ude5)      |    
                        (yy2boizah9n6vll94z | cuf6ntg4j_lumj4pox)      |    
                        l1zwxuvb407cnts      |                       
                        ivse5_zisiibgf8oum     |                       
                        (oizf0jkb_iwlm68mrw | wyit9nrrvctc4ii9rb)      |    
                        (i6q7_tpl_4f61n | dqmsf6gtvzuqhis21l)      |    
                        vz7mnovu_m51dq1      |                       
                        jicp1hi2zypaj       |                       
                        rkx2z9tuldgd39zp      |                       
                        (podz_mnetypiu7 | fkaztmo9sputf)       |    
                        (dl4pq4785d2evg | a90cuq3gcnfvujvq4t)     |    
                        a7bnvi_up37cgwlgo     |                       
                        p0wx5tkzaf886os     |                       
                        (styktg7w7fi36jw0e5n4h93 & ezupw6o2yfm5ojugrc3) |    
                        (tfcuen58mdto351cstsry5 & ezupw6o2yfm5ojugrc3) |    
                        lhx06f20_s0toyo1q7     |                       
                        tv4hqiny5afky9w |  vwmbmpalhwfnoi_0g |            
                        hfqcy171lm219z2  |  ecccb2oy3kp6vbt  |dsp656i_shm9fbrjf |  
                        v_b574hro993x |  
                        rf_x1axtwqsgz14s | h193fufzl9k9j8_bi |            
                        vhzlyir7ae3m3dx_o | brwqtymgz1q318trw |            
                        g3eepk0cdmakl1u | nybn83l8h8rmm5tk |            
                        ss1_hx3eo4rnxdbn6 | i679vkh0e1766qyk |            
                        z3kk91ocqzu25       ;                       



  wire s0aynip0upf = (v9zbczh8 | aug3vtovlhu39z) & t6_6ypj94nny67ise0x9;

  wire [19-1:0] r111cw2e83ekvdr;
  assign r111cw2e83ekvdr[3:0          ] = 4'd5;
  assign r111cw2e83ekvdr[4:4         ] = vlfahv69        ;
  assign r111cw2e83ekvdr[5:5   ] = a6x0kl79q36    ;   
  assign r111cw2e83ekvdr[6:6  ] = jgncnwo8lu01   ;
  assign r111cw2e83ekvdr[7:7] = g_oka7qgfr5inx ;
  assign r111cw2e83ekvdr[8:8 ] = zswqi_bpr6dj  ;
  assign r111cw2e83ekvdr[9:9   ] = lpac9vygdosz    ;
  assign r111cw2e83ekvdr[10:10  ] = gu1ryj7evsze   ;
  assign r111cw2e83ekvdr[11:11   ] = ujvx9ip2    ;
  assign r111cw2e83ekvdr[12:12  ] = ph174i8mt   ;
  assign r111cw2e83ekvdr[13:13   ] = sa2f4h4xeakpfnunl;

  assign r111cw2e83ekvdr[14:14  ] = m_5r0ivgcn;
  assign r111cw2e83ekvdr[15:15  ] = vjyxyga4yc;
  assign r111cw2e83ekvdr[16:16 ] = veznwo9f7pzr;
  assign r111cw2e83ekvdr[17:17  ] = re57g9q8nl7bu;
  assign r111cw2e83ekvdr[18:18 ] = cwupd7pgtwtjh;

  assign tkm5u9dl8zav4 = s0aynip0upf;
  assign eaxqugrf_ryu5rxxw41 =  r111cw2e83ekvdr;

  assign t9xs6bqphiru = jgncnwo8lu01 | g_oka7qgfr5inx | zswqi_bpr6dj;
  assign ls1dudpc    = a6x0kl79q36 | m_5r0ivgcn;
  assign tzjssx03b    = lpac9vygdosz | vjyxyga4yc;
  assign kt04okvuth   = gu1ryj7evsze| veznwo9f7pzr;
  assign cni2453cuofb    = ujvx9ip2 | re57g9q8nl7bu;
  assign kq9gup8pu2   = ph174i8mt| cwupd7pgtwtjh;



  wire nn86s_6j0i       = s3qnk2twp6   & ezupw6o2yfm5ojugrc3;
  wire k64nwvru14rm       = s3qnk2twp6   & d24iqtxvb2trplxk2m;
  wire q5tf1gw       = s3qnk2twp6   & t8jc64yc1l6q8eclq_c;
  wire sa1v919c      = s3qnk2twp6   & d0jauc9xnvhr53rq3;
  wire semw666r      = s3qnk2twp6   & tcks0htkit9weu;
  wire k2shv0srgu0krb8ve = s3qnk2twp6 & (w__ro7gwx6w331 | o6hnybbrbqkztojg | dwe8qnpoudm94xa);

  wire u0r8w9ch59lj       = g07txhn20bwh3as  & ezupw6o2yfm5ojugrc3;
  wire c41hgx9ihx       = g07txhn20bwh3as  & d24iqtxvb2trplxk2m;
  wire jitv00eenhhk       = g07txhn20bwh3as  & t8jc64yc1l6q8eclq_c;
  wire ir80nlzybrgunagd7j = g07txhn20bwh3as & (w__ro7gwx6w331 | p2f86tlrac56[2]);

  wire qhv1dh6zaqvg8rb2w    = id7i5ufppar8 & o6hnybbrbqkztojg;
  wire vvjw37emv          = id7i5ufppar8 & w__ro7gwx6w331;

  wire cp2dnt92cia          = hjxhtr2pfh;

  wire pnq529s746a01v0gox = k2shv0srgu0krb8ve;
  wire tg_wq2a0jqwopavmiul = ir80nlzybrgunagd7j;




  wire opeewkej2yt11      = j3paeay4496m & t8jc64yc1l6q8eclq_c & (uk0ahn6nnbba7[6:2] == 5'b00010);
  wire rplybbfmx488      = j3paeay4496m & t8jc64yc1l6q8eclq_c & (uk0ahn6nnbba7[6:2] == 5'b00011);
  wire vjtdrlknn3lxth5 = j3paeay4496m & t8jc64yc1l6q8eclq_c & (uk0ahn6nnbba7[6:2] == 5'b00001);
  wire eryjh8zz18fp00qql0  = j3paeay4496m & t8jc64yc1l6q8eclq_c & (uk0ahn6nnbba7[6:2] == 5'b00000);
  wire go19todx4g7uv_9  = j3paeay4496m & t8jc64yc1l6q8eclq_c & (uk0ahn6nnbba7[6:2] == 5'b00100);
  wire wj_q61p9s8ik6ntb  = j3paeay4496m & t8jc64yc1l6q8eclq_c & (uk0ahn6nnbba7[6:2] == 5'b01100);
  wire sa90h_fldec1y8   = j3paeay4496m & t8jc64yc1l6q8eclq_c & (uk0ahn6nnbba7[6:2] == 5'b01000);
  wire q8qqxf56iuu0hbc  = j3paeay4496m & t8jc64yc1l6q8eclq_c & (uk0ahn6nnbba7[6:2] == 5'b10000);
  wire ixb85e7tad2qw6e7y_  = j3paeay4496m & t8jc64yc1l6q8eclq_c & (uk0ahn6nnbba7[6:2] == 5'b10100);
  wire wolgn4jib9vw24cb = j3paeay4496m & t8jc64yc1l6q8eclq_c & (uk0ahn6nnbba7[6:2] == 5'b11000);
  wire qtmdfs7lvfjchott3al = j3paeay4496m & t8jc64yc1l6q8eclq_c & (uk0ahn6nnbba7[6:2] == 5'b11100);


  wire oo_r3ir9zo8z6zvfbo = j3paeay4496m & 
                  (~(opeewkej2yt11      |
                     rplybbfmx488      |
                     vjtdrlknn3lxth5 |
                     eryjh8zz18fp00qql0  |
                     go19todx4g7uv_9  |
                     wj_q61p9s8ik6ntb  |
                     sa90h_fldec1y8   |
                     q8qqxf56iuu0hbc  |
                     ixb85e7tad2qw6e7y_  |
                     wolgn4jib9vw24cb |
                     qtmdfs7lvfjchott3al )
                  );




  wire cydt9da18h      = rt2gdnok8 & (uk0ahn6nnbba7[6:2] == 5'b00010);
  wire ye6xa_3wfkc4q      = rt2gdnok8 & (uk0ahn6nnbba7[6:2] == 5'b00011);
  wire d896lnaa700uwskj = rt2gdnok8 & (uk0ahn6nnbba7[6:2] == 5'b00001);
  wire t10qyk84kqfrpa  = rt2gdnok8 & (uk0ahn6nnbba7[6:2] == 5'b00000);
  wire nkwt3bpu566hxe5  = rt2gdnok8 & (uk0ahn6nnbba7[6:2] == 5'b00100);
  wire opnkqtu31ik_95tot  = rt2gdnok8 & (uk0ahn6nnbba7[6:2] == 5'b01100);
  wire xs0xi0q3gmrpn2   = rt2gdnok8 & (uk0ahn6nnbba7[6:2] == 5'b01000);
  wire nf82s4nnwk5w2bh1  = rt2gdnok8 & (uk0ahn6nnbba7[6:2] == 5'b10000);
  wire gupca0jjt1piogipv  = rt2gdnok8 & (uk0ahn6nnbba7[6:2] == 5'b10100);
  wire hhsk78rsdy_5ar = rt2gdnok8 & (uk0ahn6nnbba7[6:2] == 5'b11000);
  wire rijags_148du1d = rt2gdnok8 & (uk0ahn6nnbba7[6:2] == 5'b11100);
  
  
  wire sn020cbfgrlm_e = rt2gdnok8 & 
                  (~(cydt9da18h      |
                     ye6xa_3wfkc4q      |
                     d896lnaa700uwskj |
                     t10qyk84kqfrpa  |
                     nkwt3bpu566hxe5  |
                     opnkqtu31ik_95tot  |
                     xs0xi0q3gmrpn2   |
                     nf82s4nnwk5w2bh1  |
                     gupca0jjt1piogipv  |
                     hhsk78rsdy_5ar |
                     rijags_148du1d )
                  );
  
  




  wire   v7s5fo07nb5 = (s3qnk2twp6) | (g07txhn20bwh3as) | yyd3wantj | v_a3dq6 | (mbzx7zhsly5) | nh22c0jbg5o19
                      | j3paeay4496m
                      | u_mgu2iomgss4kbb5q 
                      | no5vijin9fx5kyxd3lop2wg4d 
                      | (hschwo70vh36y   | bx5js_t0gcoh8   | y1x6fpss6_6   | hh5fb5xzanf14) 
                      | (gx2n0dmy9   | yxd3c1kl5vo15   | sbyhjyyw1   | an_cjmmfv) 
                      | (qdqvpvjvmba | pfeg45fn01up | iy0t317_b18b1 | wf8o8lzblge) 
                      | (id7i5ufppar8 |  hjxhtr2pfh | d764kpemvglzpk9 | jm6sitcu2sj | eiqmnomnjfe0 | qi_35cq273ym)
                      | rt2gdnok8
                      ;


  wire [1:0] bplrdqu945g0pwra  = 
                              vlfahv69  ? p2f86tlrac56[1:0] :
                             (d764kpemvglzpk9 | eiqmnomnjfe0 
                            | jm6sitcu2sj | qi_35cq273ym
                            | sbyhjyyw1   | an_cjmmfv 
                            | iy0t317_b18b1 | wf8o8lzblge 
                             ) ? 2'b11 : 2'b10;


  wire       xg3ql287ctjjvi = vlfahv69? p2f86tlrac56[2] : 1'b0;

  wire [29-1:0] a51ngszcxd19m;
  assign a51ngszcxd19m[3:0    ] = 4'd2;
  assign a51ngszcxd19m[4:4   ] = vlfahv69;
  assign a51ngszcxd19m[5:5   ] = s3qnk2twp6  | opeewkej2yt11 | yyd3wantj | mbzx7zhsly5 
                                                   | (hschwo70vh36y  | y1x6fpss6_6 | gx2n0dmy9  | sbyhjyyw1) 
                                                   | (qdqvpvjvmba  | iy0t317_b18b1) 
                                                    | (id7i5ufppar8 | cydt9da18h | d764kpemvglzpk9 | eiqmnomnjfe0)
                                                ;
  assign a51ngszcxd19m[6:6  ] = g07txhn20bwh3as | rplybbfmx488 | v_a3dq6 | nh22c0jbg5o19 
                                                   | u_mgu2iomgss4kbb5q
                                                   | no5vijin9fx5kyxd3lop2wg4d
                                                   | (bx5js_t0gcoh8 | hh5fb5xzanf14 | yxd3c1kl5vo15 | an_cjmmfv) 
                                                   | (pfeg45fn01up  | wf8o8lzblge) 
                                                    | (hjxhtr2pfh | ye6xa_3wfkc4q | jm6sitcu2sj | qi_35cq273ym)
                                                ;
  assign a51ngszcxd19m[28:27] =  2'b00  
                                                   | ({2{(hschwo70vh36y | bx5js_t0gcoh8 | gx2n0dmy9 | yxd3c1kl5vo15 | qdqvpvjvmba | pfeg45fn01up)}} & 2'b10) 
                                                   | ({2{(y1x6fpss6_6 | hh5fb5xzanf14 | sbyhjyyw1 | an_cjmmfv | iy0t317_b18b1 | wf8o8lzblge)}} & 2'b11) 
                                                ;
  assign a51ngszcxd19m[8:7   ] = 
                                                  u_mgu2iomgss4kbb5q ? 2'b11:
                                                  no5vijin9fx5kyxd3lop2wg4d ? 2'b11:
                                                  bplrdqu945g0pwra;
  assign a51ngszcxd19m[9:9  ] = 
                                                  xg3ql287ctjjvi;
  assign a51ngszcxd19m[10:10   ] = opeewkej2yt11 | rplybbfmx488 | cydt9da18h | ye6xa_3wfkc4q;
  assign a51ngszcxd19m[11:11    ] = j3paeay4496m & (~(opeewkej2yt11 | rplybbfmx488))
                                                |  rt2gdnok8 & (~(cydt9da18h | ye6xa_3wfkc4q));
  assign a51ngszcxd19m[12:12] = vjtdrlknn3lxth5 | d896lnaa700uwskj ;
  assign a51ngszcxd19m[13:13 ] = eryjh8zz18fp00qql0  | t10qyk84kqfrpa  ;
  assign a51ngszcxd19m[14:14 ] = wj_q61p9s8ik6ntb  | opnkqtu31ik_95tot  ;
  assign a51ngszcxd19m[15:15  ] = sa90h_fldec1y8   | xs0xi0q3gmrpn2   ;
  assign a51ngszcxd19m[16:16 ] = go19todx4g7uv_9  | nkwt3bpu566hxe5  ;
  assign a51ngszcxd19m[17:17 ] = ixb85e7tad2qw6e7y_  | gupca0jjt1piogipv  ;
  assign a51ngszcxd19m[18:18 ] = q8qqxf56iuu0hbc  | nf82s4nnwk5w2bh1  ;
  assign a51ngszcxd19m[19:19] = qtmdfs7lvfjchott3al | rijags_148du1d ;
  assign a51ngszcxd19m[20:20] = wolgn4jib9vw24cb | hhsk78rsdy_5ar ;
  assign a51ngszcxd19m[21:21 ] = (glv8ztvxphxctm | kvnjxxg7anei8786qg) ? 1'b1 : qt8cr87lzx1u; 
  assign a51ngszcxd19m[23:23 ] = jbkjansoihuv2nv; 
  assign a51ngszcxd19m[22:22   ] = ql2xoldgv6si0j;
  assign a51ngszcxd19m[24:24   ] = aw5pbsduwvhyhb3aka;
  assign a51ngszcxd19m[26:26] = wqpng9lj3ibxslk; 
  assign a51ngszcxd19m[25:25  ] = o2zokol469i9emxjt;




  assign k_y4yq3crp_zqtg = (s3qnk2twp6 | g07txhn20bwh3as | id7i5ufppar8 | hjxhtr2pfh) & 
                      (ga71__f5g1[5-1:0] == 5'b0);

  wire   wib8hsb4py2v2tg_;
  wire   rjob9x0q8su7ed2i;

  wire tcmkugn0bp2nb16 = sbyhjyyw1 | gx2n0dmy9 | qdqvpvjvmba | iy0t317_b18b1;
  wire wxeg7gajnt120 = an_cjmmfv | yxd3c1kl5vo15 | pfeg45fn01up | wf8o8lzblge;
  wire effd0iy0yg9cxfpj = gx2n0dmy9 | yxd3c1kl5vo15 | qdqvpvjvmba | pfeg45fn01up;
  wire hpmp5fw7fq25lvk5p = sbyhjyyw1 | an_cjmmfv | iy0t317_b18b1 | wf8o8lzblge;
  wire nwgcpzroopwqa;

  wire os6z_gmtxe8 = vlfahv69 ? (glv8ztvxphxctm | kvnjxxg7anei8786qg) 
                       : (tcmkugn0bp2nb16 | wxeg7gajnt120);

  wire [12-1:0] ij6wl8uax5l3kq;
  assign ij6wl8uax5l3kq[3:0        ] = 4'd7;
  assign ij6wl8uax5l3kq[4:4       ] = vlfahv69;
  assign ij6wl8uax5l3kq[6:5   ] = 2'd0;
  assign ij6wl8uax5l3kq[9:7   ] = 3'b0;
  assign ij6wl8uax5l3kq[10:10   ] = 1'b0;



  assign ij6wl8uax5l3kq[11:11] = nwgcpzroopwqa; 

  wire ob1elujf = vlfahv69 & (kzyiyt0xi8d | lz1544702tkg0u | o4tc3g036bgoap | cbru05_q5bm7);

  wire [14-1:0] ogm84pywh4cfj1;
  assign ogm84pywh4cfj1[3:0        ] = 4'd7;
  assign ogm84pywh4cfj1[4:4       ] = vlfahv69;
  assign ogm84pywh4cfj1[6:5   ] = 2'd2;
  assign ogm84pywh4cfj1[9:7   ] = k0xug5g[14:12];
  assign ogm84pywh4cfj1[10:10  ] = 1'b1;
  assign ogm84pywh4cfj1[11:11   ] = (kzyiyt0xi8d | lz1544702tkg0u);
  assign ogm84pywh4cfj1[12:12  ] = (o4tc3g036bgoap | cbru05_q5bm7);
  assign ogm84pywh4cfj1[13:13] = (lz1544702tkg0u | cbru05_q5bm7) ;

  wire pnpbz9h07ldh = vlfahv69 & (1'b0
                 | gwoe477gldf8c9e 
                 | my890tb6fuxn0ar 
                 | i_43p0nivqch83l
                 | lg8nys4yk9hgun1
                 | fz4uie4yxvn5  
                 | snxdp3tvw7a  
                 | x0c94xeqpc8nzim7  
                 | j_tdnombv0p5jwn8 
                 | rog98nkwfh96pgah1 
                 | ryz5m33fgnp6ofcw
                 | ig6dxpy3sgfnd
                 | knc4udhhcbv  
                 | vou4ap3g4kukvz7a  
                 | ou19p6zx65a  )  ;

  wire ukjorxd_z0esxtc = vlfahv69 & (1'b0
                 | vzgrcege9g3qyat  
                 | p0u65_oip3cn  
                 | qfgkmomxjwhe   
                 | v3he_44ycy65   
                 | h5gjvo_bpoph5i   
                 | hjq039vacscr  
                 | n6f1xma1ku0cqc9  
                 | ns2ccb8p4kf3o   
                 | wy5oiwkuovruvc   
                 | mtnmu5bzb5z9)  ;

  wire cdlm5zrwv = pnpbz9h07ldh | ukjorxd_z0esxtc;

  wire qic9a7eczdf = ( 
                   j_tdnombv0p5jwn8 
                 | rog98nkwfh96pgah1 
                 | ryz5m33fgnp6ofcw
                 | ig6dxpy3sgfnd
                 | knc4udhhcbv  
                 | vou4ap3g4kukvz7a  
                 | ou19p6zx65a  
                 | hjq039vacscr  
                 | n6f1xma1ku0cqc9  
                 | ns2ccb8p4kf3o   
                 | wy5oiwkuovruvc   
                 | mtnmu5bzb5z9)  ;

  wire [24-1:0] q1nf0s6751pdaj8a;
  assign q1nf0s6751pdaj8a[3:0        ] = 4'd7;
  assign q1nf0s6751pdaj8a[4:4       ] = vlfahv69;
  assign q1nf0s6751pdaj8a[6:5    ] = 2'd1;
  assign q1nf0s6751pdaj8a[9:7     ] = pnpbz9h07ldh ? k0xug5g[14:12] : 3'b0;
  assign q1nf0s6751pdaj8a[10:10  ] = pnpbz9h07ldh ? 1'b1 : 1'b0;
  assign q1nf0s6751pdaj8a[11:11 ] = gwoe477gldf8c9e | j_tdnombv0p5jwn8; 
  assign q1nf0s6751pdaj8a[12:12 ] = my890tb6fuxn0ar | rog98nkwfh96pgah1;
  assign q1nf0s6751pdaj8a[13:13] = i_43p0nivqch83l | ryz5m33fgnp6ofcw;
  assign q1nf0s6751pdaj8a[14:14] = lg8nys4yk9hgun1 | ig6dxpy3sgfnd;
  assign q1nf0s6751pdaj8a[15:15  ] = fz4uie4yxvn5  | knc4udhhcbv ;
  assign q1nf0s6751pdaj8a[16:16  ] = snxdp3tvw7a  | vou4ap3g4kukvz7a ;
  assign q1nf0s6751pdaj8a[17:17  ] = x0c94xeqpc8nzim7  | ou19p6zx65a ;
  assign q1nf0s6751pdaj8a[18:18  ] = vzgrcege9g3qyat  | hjq039vacscr ;
  assign q1nf0s6751pdaj8a[19:19  ] = p0u65_oip3cn  | n6f1xma1ku0cqc9 ;
  assign q1nf0s6751pdaj8a[20:20   ] = qfgkmomxjwhe   | ns2ccb8p4kf3o  ;
  assign q1nf0s6751pdaj8a[21:21   ] = v3he_44ycy65   | wy5oiwkuovruvc  ;
  assign q1nf0s6751pdaj8a[22:22   ] = h5gjvo_bpoph5i   | mtnmu5bzb5z9  ;
  assign q1nf0s6751pdaj8a[23:23] = qic9a7eczdf;



  wire qgo9xkq = vlfahv69 & (1'b0
                 | iz_sm_7y_ixfw1btmz 
                 | uz6maeeehzsn6uzwxk
                 | dywxta8oxdnj1q9i0d 
                 | zqz28qv7052ajkf7
                 | tnkhekmenrbyvq 
                 | gsqes4kpzyh7s4 
                 | th_rx8vbgu0ydrx 
                 | glahkq0rwcrj086j7k1j
                 | i_oja_fou8xg9_ 
                 | jz2t1e591yva8m5
                 | hx05sow34f5nxv 
                 | iboby_h0cqqucgnxw
                 | nu4l8_3i80k9r9huos 
                 | wjhbw3uh3oljyutu2gel
                 | knqkb_9b7915rg 
                 | jlez7xntekztmffn06
                 | q1mnx00q446iezuqt 
                 | bvcgz8q5ffa32w7);


  wire uiogf37b = vlfahv69 & (1'b0
                 | nlb5566a2kkzrak 
                 | t82iq62ywf1u_5
                 | byqkkp26xdsszd
                 | gkj8ltdpe4tcqini4h
                 | l6qpfpq3ro_9gr
                 | nxf52k3xp6im5o6p3
                 | vdmyb8x4qmwi7on2 
                 | tfoxw8ia_xdt0
                 | f128ccj13txxdwpl
                 | u72qi7gmhj37d_h5c
                 | va7j9_tx3li0xd
                 | tr03xi8fsjspsc
                 | qgo9xkq);

  wire [38-1:0] lm7r3hwrkp41v02nig;
  assign lm7r3hwrkp41v02nig[3:0        ] = 4'd7;
  assign lm7r3hwrkp41v02nig[4:4       ] = vlfahv69;
  assign lm7r3hwrkp41v02nig[6:5    ] = 2'd3;
  assign lm7r3hwrkp41v02nig[9:7     ] = qgo9xkq ? k0xug5g[14:12] : 3'b0;
  assign lm7r3hwrkp41v02nig[10:10  ] = qgo9xkq ? 1'b1 : 1'b0;
  assign lm7r3hwrkp41v02nig[11:11 ] = nlb5566a2kkzrak  | vdmyb8x4qmwi7on2  ; 
  assign lm7r3hwrkp41v02nig[12:12] = t82iq62ywf1u_5 | tfoxw8ia_xdt0 ;
  assign lm7r3hwrkp41v02nig[13:13] = byqkkp26xdsszd | f128ccj13txxdwpl ;
  assign lm7r3hwrkp41v02nig[14:14 ] = gkj8ltdpe4tcqini4h ;
  assign lm7r3hwrkp41v02nig[15:15 ] = va7j9_tx3li0xd ;
  assign lm7r3hwrkp41v02nig[16:16] = l6qpfpq3ro_9gr | u72qi7gmhj37d_h5c ;
  assign lm7r3hwrkp41v02nig[17:17 ] = nxf52k3xp6im5o6p3 ;
  assign lm7r3hwrkp41v02nig[18:18 ] = tr03xi8fsjspsc ;
  assign lm7r3hwrkp41v02nig[19:19 ] = iz_sm_7y_ixfw1btmz ;
  assign lm7r3hwrkp41v02nig[20:20] = uz6maeeehzsn6uzwxk;
  assign lm7r3hwrkp41v02nig[21:21 ] = dywxta8oxdnj1q9i0d ;
  assign lm7r3hwrkp41v02nig[22:22] = zqz28qv7052ajkf7;
  assign lm7r3hwrkp41v02nig[23:23 ] = tnkhekmenrbyvq ;
  assign lm7r3hwrkp41v02nig[24:24 ] = gsqes4kpzyh7s4 ;
  assign lm7r3hwrkp41v02nig[25:25 ] = th_rx8vbgu0ydrx ;
  assign lm7r3hwrkp41v02nig[26:26] = glahkq0rwcrj086j7k1j;
  assign lm7r3hwrkp41v02nig[27:27 ] = i_oja_fou8xg9_ ;
  assign lm7r3hwrkp41v02nig[28:28] = jz2t1e591yva8m5;
  assign lm7r3hwrkp41v02nig[30:30 ] = hx05sow34f5nxv ;
  assign lm7r3hwrkp41v02nig[31:31] = iboby_h0cqqucgnxw;
  assign lm7r3hwrkp41v02nig[32:32 ] = nu4l8_3i80k9r9huos ;
  assign lm7r3hwrkp41v02nig[33:33] = wjhbw3uh3oljyutu2gel;
  assign lm7r3hwrkp41v02nig[34:34 ] = knqkb_9b7915rg ;
  assign lm7r3hwrkp41v02nig[35:35] = jlez7xntekztmffn06;
  assign lm7r3hwrkp41v02nig[36:36 ] = q1mnx00q446iezuqt ;
  assign lm7r3hwrkp41v02nig[37:37] = bvcgz8q5ffa32w7;
  assign lm7r3hwrkp41v02nig[29:29] = vdmyb8x4qmwi7on2 | tfoxw8ia_xdt0 | f128ccj13txxdwpl | u72qi7gmhj37d_h5c;

  
  
  
  




  wire pvtposb4yd5tpd95  = lrptc0hyjyd7hdoypa0_g 
                        & y2hcqn22lsrsl 
                        & jnhdayjoseb 
                        & ezupw6o2yfm5ojugrc3 
                        & adw7hffbin 
                        & w0s41titqc28jdt 
                        & d6r44hi25ixatafeu1 
                        & (dlmxb1[1:0] == 2'b00); 

  wire smz1g6gnii8n7mg9_fs  = yf083xcjpnohrzqky4 
                        & sauhc6ef6pqjm_w4 
                        & oezgh2bhqupmgh2 
                        & dwe8qnpoudm94xa 
                        & bgecyjs80sbc 
                        & f_575odq4qxl04 
                        & w3imaozzd_v_wb6wo 
                        & (dlmxb1[1:0] == 2'b11); 

  wire ukx4cgxh08fqx3hu  = mg22fa39qkmi1381_ 
                        & ezupw6o2yfm5ojugrc3 
                        & adw7hffbin     
                        & w0s41titqc28jdt 
                        & d6r44hi25ixatafeu1 
                        & (dlmxb1[1:0] == 2'b00); 

  wire xuqk_ks14k6o5144w  = f9zuwwm5sc91jd4
                        & dwe8qnpoudm94xa 
                        & bgecyjs80sbc 
                        & f_575odq4qxl04 
                        & w3imaozzd_v_wb6wo 
                        & (dlmxb1[1:0] == 2'b11);

  wire ctcwxdialrasri5u6guy = vlfahv69 ?  (pvtposb4yd5tpd95 | smz1g6gnii8n7mg9_fs)
                              :  (ukx4cgxh08fqx3hu | xuqk_ks14k6o5144w);






  wire bqywdsjnr1r6icc0 = 
                      (~adw7hffbin) & (
                    (
                      (~cgfh21c1qcp) & (~g07txhn20bwh3as)
                    & (~dw61vkalbiqitxbxy8n0)
                    & (~waejh__hl02blsw4eau2ir6332zz) 
                    & (~hjxhtr2pfh)
                    )
                   );




  wire chso39421msvbkl9a = isxv0tqhyam | r5qet1mocbtcig | tx04m_rvbl9sow;










  wire hegurso01yv4i =
                     u_mgu2iomgss4kbb5q |
                     no5vijin9fx5kyxd3lop2wg4d |
                  (
                      (~jnhdayjoseb) & (
                    (
                      (~hwj750kj)
                    & (~ccbtxbyh0qmcdfa)
                    & (~h20g0j2jt)
                    & (~dw61vkalbiqitxbxy8n0)
                    & (~waejh__hl02blsw4eau2ir6332zz)
                    & (~nt0rwqyh45801)
                    & (~ae9uh2qsyem1utk9)
                    & (~vv6pnkge7dhr1ay_)
                    )
                   )
                  );







  wire hgjytyuf89rdi = (~y2hcqn22lsrsl) & (
                (
                 (cgfh21c1qcp)
               | (g07txhn20bwh3as)
               | (v9zbczh8)
               | (j3paeay4496m & (~opeewkej2yt11))
               | (t61y7hkwkrvm7s & ~eshy3jgtzqwpnq)
               | (aug3vtovlhu39z)
               | (hjxhtr2pfh)
               | (rt2gdnok8 & (~cydt9da18h))
               | (cicq2g9r_bh93)
                 )
                 );

  wire [64-1:0]  bezlndbgd7ln = { 
                               {(64-12){pq5pe3yehrqxr[31]}} 
                              , pq5pe3yehrqxr[31:20]
                             };

  wire [64-1:0]  en3fz149rzhd = {
                               {(64-12){pq5pe3yehrqxr[31]}} 
                              , pq5pe3yehrqxr[31:25] 
                              , pq5pe3yehrqxr[11:7]
                             };


  wire [64-1:0]  xwc1pi93ll_d7 = {
                               {(64-13){pq5pe3yehrqxr[31]}} 
                              , pq5pe3yehrqxr[31] 
                              , pq5pe3yehrqxr[7] 
                              , pq5pe3yehrqxr[30:25] 
                              , pq5pe3yehrqxr[11:8]
                              , 1'b0
                              };

  wire [64-1:0]  wcpmibamftma = {{(64-32){1'b0}},pq5pe3yehrqxr[31:12],12'b0};
  wire [64-1:0]  sk8lo0tx5lvyk0edhmg = {{(64-32){pq5pe3yehrqxr[31]}},pq5pe3yehrqxr[31:12],12'b0};

  wire [64-1:0]  bmktk5ykhzpq6 = {
                               {(64-21){pq5pe3yehrqxr[31]}} 
                              , pq5pe3yehrqxr[31] 
                              , pq5pe3yehrqxr[19:12] 
                              , pq5pe3yehrqxr[20] 
                              , pq5pe3yehrqxr[30:21]
                              , 1'b0
                              };





  wire lbvhc62mxiulgy5 = it3sb6rq7z2i67 | sa6649too5v5 | s3qnk2twp6 | h877ps0r0cih1_w_ | id7i5ufppar8;
  wire xawot5lgffrfuwnzz = sa6649too5v5;
  wire [64-1:0]  hf_ehpaimuswmut = bezlndbgd7ln;



  wire jtdc8xpvxixw9g = hwj750kj;

  wire etjqvm3qe3vblk3tt1te = ccbtxbyh0qmcdfa;



  wire x170amfl2b09v5m7e = h20g0j2jt;
  wire l9digw11aam6nd6rb9 = h20g0j2jt;
  wire [64-1:0]  qytu41_x5zlegr = bmktk5ykhzpq6;



  wire jqir3okx_oxcqz = cgfh21c1qcp;
  wire o6soq_mfr7s9lh51rhx5 = cgfh21c1qcp | k0glq1z9c20ujfyc;         
  wire [64-1:0]  x8lnalqbfmpei = k0glq1z9c20ujfyc ? e2rml0d5xlemgdqf2a : xwc1pi93ll_d7;



  wire l98vs320d51swn4g = g07txhn20bwh3as | hjxhtr2pfh;









  wire gd9sgaffk92l6drt = mbzx7zhsly5;
  wire [64-1:0]  g2lwvw9vfsdbpofi3 ={
                          {(64-8){1'b0}}
                        , tm0dvbtguid67[3:2]
                        , tm0dvbtguid67[12]
                        , tm0dvbtguid67[6:4]
                        , 2'b0
                         };

  wire w09h3we2skwms5gwum6rj = eiqmnomnjfe0;
  wire [64-1:0]  djngfc30604xfdimoq8 ={
                          {(64-9){1'b0}}
                        , tm0dvbtguid67[4:2]
                        , tm0dvbtguid67[12]
                        , tm0dvbtguid67[6:5]
                        , 3'b0
                         };







  wire b0i56ck3zq4jygridon5w4 = mhz85qp | rqj6hf1k9f | w5wv66al4ks3x
                   | afnn1is_f9szbi | h__4na2w1 | bs3b85ifu | srcanpuv42e7t;
  wire [64-1:0]  xsp528jeqsyil8ctqv ={
                          {(64-6){tm0dvbtguid67[12]}}
                        , tm0dvbtguid67[12]
                        , tm0dvbtguid67[6:2]
                         };



  wire ruoecoltz5fh1u_uioq = qvq4uyy0b;
  wire [64-1:0]  vnzuwr41a04js8 ={
                          {(64-18){tm0dvbtguid67[12]}}
                        , tm0dvbtguid67[12]
                        , tm0dvbtguid67[6:2]
                        , 12'b0
                         };



  wire gvzpjholr_265fkk_gjsaa = einxry70u73t166q;
  wire [64-1:0]  b6h2el009zfreguoxk ={
                          {(64-10){tm0dvbtguid67[12]}}
                        , tm0dvbtguid67[12]
                        , tm0dvbtguid67[4]
                        , tm0dvbtguid67[3]
                        , tm0dvbtguid67[5]
                        , tm0dvbtguid67[2]
                        , tm0dvbtguid67[6]
                        , 4'b0
                         };



  wire m1p7je1f8iqvuiqtsxy = nh22c0jbg5o19;
  wire [64-1:0]  igsqeqei9b_m ={
                          {(64-8){1'b0}}
                        , tm0dvbtguid67[8:7]
                        , tm0dvbtguid67[12:9]
                        , 2'b0
                         };

  wire jhnz8_4pcxii6op9f_2o = qi_35cq273ym;
  wire [64-1:0]  dq9y438n_c9145r2 ={
                          {(64-9){1'b0}}
                        , tm0dvbtguid67[9:7]
                        , tm0dvbtguid67[12:10]
                        , 3'b0
                         };


  wire ukevfivu49g_lnhx = tdceg4r4ocywxjcsuv;
  wire [64-1:0]  d3ni905810iog5yn ={
                          {(64-10){1'b0}}
                        , tm0dvbtguid67[10:7]
                        , tm0dvbtguid67[12]
                        , tm0dvbtguid67[11]
                        , tm0dvbtguid67[5]
                        , tm0dvbtguid67[6]
                        , 2'b0
                         };



  wire w_gnrh8qm5y15liydhp = yyd3wantj;
  wire [64-1:0]  azcp5tz0ja9e ={
                          {(64-7){1'b0}}
                        , tm0dvbtguid67[5]
                        , tm0dvbtguid67[12]
                        , tm0dvbtguid67[11]
                        , tm0dvbtguid67[10]
                        , tm0dvbtguid67[6]
                        , 2'b0
                         };

  wire dpp1njvi_j743ql7v_op = d764kpemvglzpk9;                 
  wire [64-1:0]  ukb_03_4r5h4pu ={
                          {(64-8){1'b0}}
                        , tm0dvbtguid67[6]
                        , tm0dvbtguid67[5]
                        , tm0dvbtguid67[12]
                        , tm0dvbtguid67[11]
                        , tm0dvbtguid67[10]
                        , 3'b0
                         };


  wire c1_xssiqdzyhatzdgcwr = v_a3dq6;
  wire [64-1:0]  grxnrl07y_4cziq ={
                          {(64-7){1'b0}}
                        , tm0dvbtguid67[5]
                        , tm0dvbtguid67[12]
                        , tm0dvbtguid67[11]
                        , tm0dvbtguid67[10]
                        , tm0dvbtguid67[6]
                        , 2'b0
                         };

   wire qhz11v1fatt4mcjxq0m4a = jm6sitcu2sj;
   wire [64-1:0]  i6jkk5pbwa_884xd1 ={
                          {(64-8){1'b0}}
                        , tm0dvbtguid67[6]
                        , tm0dvbtguid67[5]
                        , tm0dvbtguid67[12]
                        , tm0dvbtguid67[11]
                        , tm0dvbtguid67[10]
                        , 3'b0
                         };




  wire dll6xk9dzqf_mh1dtz = tez8bez5l4r | zh62ppn61_4yw4;
  wire [64-1:0]  ucjofgpggsfb0 ={
                          {(64-9){tm0dvbtguid67[12]}}
                        , tm0dvbtguid67[12]
                        , tm0dvbtguid67[6:5]
                        , tm0dvbtguid67[2]
                        , tm0dvbtguid67[11:10]
                        , tm0dvbtguid67[4:3]
                        , 1'b0
                         };
  wire [64-1:0]  xoxse1yov4vm01rl = ucjofgpggsfb0;




  wire s4kndwtbl8fxmiyi3m = ei1me6y0 | e_qxxtaevvw;
  wire [64-1:0]  hx6p43b2pspg_ ={
                          {(64-12){tm0dvbtguid67[12]}}
                        , tm0dvbtguid67[12]
                        , tm0dvbtguid67[8]
                        , tm0dvbtguid67[10:9]
                        , tm0dvbtguid67[6]
                        , tm0dvbtguid67[7]
                        , tm0dvbtguid67[2]
                        , tm0dvbtguid67[11]
                        , tm0dvbtguid67[5:3]
                        , 1'b0
                         };
  wire [64-1:0]  q6dj3cn7jeic88g0ok = hx6p43b2pspg_;



  wire [64-1:0]  onxwi3lt3vee8230ahq9 = 64'b0;








  wire [64-1:0]  egbzq3jp2wqrziqrgkpxo  = bezlndbgd7ln;
  wire [64-1:0]  t89ie00ykt7rqgf5ul_1zt = en3fz149rzhd;
  wire [64-1:0]  tqeq1dm5bhi = 
                     ({64{lbvhc62mxiulgy5}} & bezlndbgd7ln)
                   | ({64{l98vs320d51swn4g}} & en3fz149rzhd)
                   | ({64{jqir3okx_oxcqz}} & xwc1pi93ll_d7)
                   | ({64{jtdc8xpvxixw9g}} & wcpmibamftma)
                   | ({64{etjqvm3qe3vblk3tt1te}} & sk8lo0tx5lvyk0edhmg)
                   | ({64{x170amfl2b09v5m7e}} & bmktk5ykhzpq6)
                   | ({64{u_mgu2iomgss4kbb5q}} & ({{(64-5){1'b0}},ga71__f5g1}<<2))  
                   | ({64{no5vijin9fx5kyxd3lop2wg4d}} & ({{(64-5){1'b0}},ga71__f5g1}<<2))  
                   ;

  wire  utnmorebychmpkqe = 
                     lbvhc62mxiulgy5
                   | l98vs320d51swn4g
                   | jqir3okx_oxcqz
                   | jtdc8xpvxixw9g
                   | etjqvm3qe3vblk3tt1te
                   | x170amfl2b09v5m7e
                   | u_mgu2iomgss4kbb5q
                   | no5vijin9fx5kyxd3lop2wg4d
                   ;

  wire [64-1:0]  ksfckote0z60c = 
                     ({64{gd9sgaffk92l6drt   }} & g2lwvw9vfsdbpofi3)
                   | ({64{b0i56ck3zq4jygridon5w4  }} & xsp528jeqsyil8ctqv)
                   | ({64{ruoecoltz5fh1u_uioq }} & vnzuwr41a04js8)
                   | ({64{gvzpjholr_265fkk_gjsaa}} & b6h2el009zfreguoxk)
                   | ({64{m1p7je1f8iqvuiqtsxy   }} & igsqeqei9b_m)
                   | ({64{ukevfivu49g_lnhx   }} & d3ni905810iog5yn)
                   | ({64{w_gnrh8qm5y15liydhp    }} & azcp5tz0ja9e)
                   | ({64{c1_xssiqdzyhatzdgcwr    }} & grxnrl07y_4cziq)
                   | ({64{dll6xk9dzqf_mh1dtz    }} & ucjofgpggsfb0)
                   | ({64{s4kndwtbl8fxmiyi3m    }} & hx6p43b2pspg_)
                   | ({64{dpp1njvi_j743ql7v_op  }} & ukb_03_4r5h4pu)
                   | ({64{qhz11v1fatt4mcjxq0m4a  }} & i6jkk5pbwa_884xd1)
                   | ({64{w09h3we2skwms5gwum6rj }} & djngfc30604xfdimoq8)
                   | ({64{jhnz8_4pcxii6op9f_2o }} & dq9y438n_c9145r2)
                   ;

  wire z5j5j7h24q3p52 = 
                     gd9sgaffk92l6drt   
                   | b0i56ck3zq4jygridon5w4  
                   | ruoecoltz5fh1u_uioq 
                   | gvzpjholr_265fkk_gjsaa
                   | m1p7je1f8iqvuiqtsxy   
                   | ukevfivu49g_lnhx   
                   | w_gnrh8qm5y15liydhp    
                   | c1_xssiqdzyhatzdgcwr    
                   | dll6xk9dzqf_mh1dtz    
                   | s4kndwtbl8fxmiyi3m   
                   | dpp1njvi_j743ql7v_op
                   | qhz11v1fatt4mcjxq0m4a
                   | w09h3we2skwms5gwum6rj
                   | jhnz8_4pcxii6op9f_2o
                   ;


  assign qt8cr87lzx1u = vlfahv69 ? utnmorebychmpkqe : z5j5j7h24q3p52; 

  assign t05leas4w4r = vlfahv69 ? tqeq1dm5bhi : ksfckote0z60c;

  
  assign nwgcpzroopwqa = os6z_gmtxe8;

  wire [64-1:0]  u5l2osbbofl1q4 = glv8ztvxphxctm ? egbzq3jp2wqrziqrgkpxo : t89ie00ykt7rqgf5ul_1zt;
  wire [64-1:0]  sc_kd_kbclahr_e76 = 
                     ({64{pfeg45fn01up }} & igsqeqei9b_m)
                   | ({64{wf8o8lzblge }} & dq9y438n_c9145r2)
                   | ({64{yxd3c1kl5vo15   }} & grxnrl07y_4cziq)
                   | ({64{an_cjmmfv   }} & i6jkk5pbwa_884xd1)
                   | ({64{gx2n0dmy9   }} & azcp5tz0ja9e)
                   | ({64{sbyhjyyw1   }} & ukb_03_4r5h4pu)
                   | ({64{qdqvpvjvmba }} & g2lwvw9vfsdbpofi3)
                   | ({64{iy0t317_b18b1 }} & djngfc30604xfdimoq8)
                   ;
  assign pxhhgm9746n = vlfahv69 ? u5l2osbbofl1q4 : sc_kd_kbclahr_e76;

  wire b7nkstim3k = 
              1'b0
            | uiogf37b
            | ob1elujf
              ;
  assign g5usf8ixwjaxjs1m = 
              ({48{ob1elujf}} & {{48-14{1'b0}},ogm84pywh4cfj1})
            | ({48{uiogf37b}} & {{48-38{1'b0}},lm7r3hwrkp41v02nig})
              ;
  assign hhj5975j18r0n =  ({48{cdlm5zrwv}} & {{48-24{1'b0}},q1nf0s6751pdaj8a});
  assign d40y0va2l7xzj = cdlm5zrwv;

















  assign vfye1vj155_k = ei82smlw45m;
  assign vujduks2o30 = v7s5fo07nb5;
  assign y4zqru1tedm = khaw8p;
  assign q1coyps2cz7xe = a7bzgrh;
  assign oli3_udj80h6urj   = b7nkstim3k;



  assign zj0wqwminaxn = ({{48-47{1'b0}},deq9tleqxy3fq} & {48{vfye1vj155_k}}) 
                      | ({{48-29{1'b0}},a51ngszcxd19m} & {48{vujduks2o30}}) 
                      | ({{48-34{1'b0}},loymwnjzrl_cl} & {48{y4zqru1tedm}}) 
                      | ({{48-27{1'b0}},krezi5k4lo8g} & {48{q1coyps2cz7xe}})




                      ;

  wire wri2knqd9wtnw = 
              ei82smlw45m
            | v7s5fo07nb5
            | khaw8p
            | b7nkstim3k
            | cdlm5zrwv
            | a7bzgrh
            | s0aynip0upf
            | sibtd2rf5j 
            ;

  assign qzdlalytscynhz1 =   al4xeg8mukgfg
                       | piwiqvrjoq
                       | s1woka0byzgo
                       | wi_dfzp70x09hm1m
                       | jdyqycv3wdp2sgy
                       | fpwql5ik7_sp0
                       ;

  wire fzxbs1cvbln1tpmeb_h =
                         (zziyl6t8rs22kz2 | nt0rwqyh45801)
                       | ((fb2hmea7xsh48i | ae9uh2qsyem1utk9) & ~jnhdayjoseb)
                       | ((k7_rcb9pbl | vv6pnkge7dhr1ay_) & ~jnhdayjoseb)
                       ;

  wire [11:0] e1go3iu = pq5pe3yehrqxr[31:20];

  wire zjd3xkagpssdo = fzxbs1cvbln1tpmeb_h & 
                        (
                            (e1go3iu == 12'h7cc)
                          | (e1go3iu == 12'h5cc)
                          | (e1go3iu == 12'h4cc)
                        )
                        ;

  assign ch8qv98q9xu469etyz8oj = 
              1'b0

            | l143yo227i5fe5s3    
            | cicq2g9r_bh93     
            | zjd3xkagpssdo 
            ;



  wire oc5hvlivuu5m4il_  = lr08s8a1cosklchm4m;
  wire mlmxilw0ul2smb4qj  = mbzx7zhsly5 | qdqvpvjvmba | iy0t317_b18b1 | mhz85qp | br9ybmw_8qr_xw4ojzr | rqj6hf1k9f | w5wv66al4ks3x | eiqmnomnjfe0 | srcanpuv42e7t; 
  wire d5eruydc6areuii2hl = nh22c0jbg5o19 | pfeg45fn01up | wf8o8lzblge | qi_35cq273ym; 
  wire cfx_w6vuaoga0no4 = tdceg4r4ocywxjcsuv; 
  wire kq82kshd_pizpgc  = yyd3wantj | gx2n0dmy9 | sbyhjyyw1 | d764kpemvglzpk9; 
  wire zi1eyt7b9_t6nrk  = v_a3dq6 | yxd3c1kl5vo15 | an_cjmmfv | pjq11l4lomf3lrph | jm6sitcu2sj | cm7ij9pf198f0ifu | ai1ohlxb9k0vgo1d9; 
  wire uvzwbt2hqdfu1uhwlwk  = tez8bez5l4r | zh62ppn61_4yw4 | h__4na2w1 | afnn1is_f9szbi | bs3b85ifu | ai1ohlxb9k0vgo1d9; 
  wire bdi73zoss0yjl_lzgm  = ei1me6y0 | e_qxxtaevvw; 








  wire os3ot61nnenwcn07o   = oc5hvlivuu5m4il_ & 1'b1;
  wire c62bp44094ap3hls93y   = oc5hvlivuu5m4il_ & 1'b1;
  wire ajcak8n6efgb0a7    = oc5hvlivuu5m4il_ & 1'b1;
  wire [5-1:0] ptls2qbpekw776 = ekodeh8usegq ? 5'd0 : ag9ylluguwcr[5-1:0];
  wire [5-1:0] kqalxxzfv7s85 = tbilhd3n1v[5-1:0];

  wire [5-1:0] r8qjp6txwnbzt  = (wgc_484cnth5 | w72sj0ys3h3)? 
                 {{5-1{1'b0}},tm0dvbtguid67[12]} : z7cl6tvk[5-1:0];







  wire z18i84zj8pggjnu0ax   = mlmxilw0ul2smb4qj & 1'b1;
  wire zjvhftiagb7l65bh5i   = mlmxilw0ul2smb4qj & 1'b0;
  wire emvc9gbmzqk07ivf8bbc    = mlmxilw0ul2smb4qj & 1'b1;
  wire [5-1:0] d1_1deih4nf7 = (mbzx7zhsly5 | qdqvpvjvmba | iy0t317_b18b1 | eiqmnomnjfe0) ? 5'd2 :
                                  (mhz85qp | qvq4uyy0b) ? 5'd0 : ag9ylluguwcr[5-1:0];
  wire [5-1:0] t7w49hivsdeeyh_0 = 5'd0;
  wire [5-1:0] cvbuf0xszkg8z2t  = z7cl6tvk[5-1:0];



  wire x9c_afdnfztrc0iq4bhv  = d5eruydc6areuii2hl & 1'b1;
  wire cv0piv5zky6kq_5rvsn  = d5eruydc6areuii2hl & 1'b1;
  wire edbnrxdg88apcxf9_wz   = d5eruydc6areuii2hl & 1'b0;
  wire [5-1:0] vywos882h0078 = 5'd2;
  wire [5-1:0] z1fntw6i8wctgcl7r = tbilhd3n1v[5-1:0];
  wire [5-1:0] g203zwhpqmo7  = 5'd0;



  wire q9n7zhbv_nvwvm2qr2z = cfx_w6vuaoga0no4 & 1'b1;
  wire usm8jjd3d6kllywh9w6 = cfx_w6vuaoga0no4 & 1'b0;
  wire io39eu_nclgfwg1dh4eq4  = cfx_w6vuaoga0no4 & 1'b1;
  wire [5-1:0] y10pdwkv_hm6nu3  = 5'd2;
  wire [5-1:0] sooa2hj7jwt64i  = 5'd0;
  wire [5-1:0] tvzetpi1oen5ik  = oduuhk6i[5-1:0];



  wire tpzgpeqjh4w3ruqiwiux  = kq82kshd_pizpgc & 1'b1;
  wire wqwc2zh6986p0sdox  = kq82kshd_pizpgc & 1'b0;
  wire x8wzvkf7gc6hluh4hx   = kq82kshd_pizpgc & 1'b1;
  wire [5-1:0] liq97mheu0vd41is = yq79t1_13[5-1:0];
  wire [5-1:0] w7tuyx3s7209e = 5'd0;
  wire [5-1:0] c1lj39gyj2y  = oduuhk6i[5-1:0];




  wire mx7zleq35h8yivtuy  = zi1eyt7b9_t6nrk & 1'b1;
  wire w663a70cvxnae9fzz  = zi1eyt7b9_t6nrk & 1'b1;
  wire tb6dx9vbazjt_ikq5   = zi1eyt7b9_t6nrk & pjq11l4lomf3lrph | cm7ij9pf198f0ifu | ai1ohlxb9k0vgo1d9;
  wire [5-1:0] p6n7b7fda8iworcx = yq79t1_13[5-1:0];
  wire [5-1:0] wc5_xepdh0nvxo = cjywp5cfm[5-1:0];
  wire [5-1:0] e9ak1p3yk1_1  = yq79t1_13[5-1:0];




  wire v73s5mmrt7tt3gqn7gqvy  = uvzwbt2hqdfu1uhwlwk & 1'b1;
  wire itidxzq9m2o2306pyw077  = uvzwbt2hqdfu1uhwlwk & (tez8bez5l4r | zh62ppn61_4yw4);
  wire brrszlfkyivox7jern   = uvzwbt2hqdfu1uhwlwk & (~(tez8bez5l4r | zh62ppn61_4yw4));
  wire [5-1:0] pb5vat5kfwq0 = yq79t1_13[5-1:0];
  wire [5-1:0] j4x2ke88_rem8083g = 5'd0;
  wire [5-1:0] d0cjbhhdw6oe  = yq79t1_13[5-1:0];




  wire a0xx9d_tpq8imwhtff  = bdi73zoss0yjl_lzgm & 1'b0;
  wire vl183kzeu77tapzyno  = bdi73zoss0yjl_lzgm & 1'b0;
  wire tlncpd0m_kefu0aje   = bdi73zoss0yjl_lzgm & 1'b1;
  wire [5-1:0] hbo5xxllemuw = 5'd0;
  wire [5-1:0] e_sgv6k4y4pmgw89 = 5'd0;
  wire [5-1:0] s5izacjghu1  = ei1me6y0 ? 5'd0 : 5'd1;









  wire j9zngxhw7hhb7wr81 = os3ot61nnenwcn07o | z18i84zj8pggjnu0ax | x9c_afdnfztrc0iq4bhv;
  wire jmima8oe0kbtp = c62bp44094ap3hls93y | zjvhftiagb7l65bh5i | cv0piv5zky6kq_5rvsn;
  wire pqvvwub0du2hsy2pbnk  = ajcak8n6efgb0a7  | emvc9gbmzqk07ivf8bbc  | edbnrxdg88apcxf9_wz;

  wire irbju9_cuzmdf155y4 = q9n7zhbv_nvwvm2qr2z|tpzgpeqjh4w3ruqiwiux|mx7zleq35h8yivtuy|v73s5mmrt7tt3gqn7gqvy|a0xx9d_tpq8imwhtff;
  wire axnh5gjxafoa13jl10 = usm8jjd3d6kllywh9w6|wqwc2zh6986p0sdox|w663a70cvxnae9fzz|itidxzq9m2o2306pyw077|vl183kzeu77tapzyno;
  wire m2ulf0uhnahhennrj  = io39eu_nclgfwg1dh4eq4 |x8wzvkf7gc6hluh4hx |tb6dx9vbazjt_ikq5 |brrszlfkyivox7jern |tlncpd0m_kefu0aje ;

  wire y37z_dzbgh = (j9zngxhw7hhb7wr81 | irbju9_cuzmdf155y4);
  wire rfxb0v1yejd7l = (jmima8oe0kbtp | axnh5gjxafoa13jl10);
  wire gwc5qjrcohbdez = 1'b0;
  wire yjigfdj36u7d3yg = (pqvvwub0du2hsy2pbnk  | m2ulf0uhnahhennrj);


  assign u2apzx0s0_ms = 
         ({5{os3ot61nnenwcn07o }} & ptls2qbpekw776)
       | ({5{z18i84zj8pggjnu0ax }} & d1_1deih4nf7)
       | ({5{x9c_afdnfztrc0iq4bhv}} & vywos882h0078)
       | ({5{q9n7zhbv_nvwvm2qr2z}} & y10pdwkv_hm6nu3)
       | ({5{tpzgpeqjh4w3ruqiwiux}}  & liq97mheu0vd41is)
       | ({5{mx7zleq35h8yivtuy}}  & p6n7b7fda8iworcx)
       | ({5{v73s5mmrt7tt3gqn7gqvy}}  & pb5vat5kfwq0)
       | ({5{a0xx9d_tpq8imwhtff}}  & hbo5xxllemuw)
       ;

  assign cyoz2x_qbs1p = 
         ({5{c62bp44094ap3hls93y }} & kqalxxzfv7s85)
       | ({5{zjvhftiagb7l65bh5i }} & t7w49hivsdeeyh_0)
       | ({5{cv0piv5zky6kq_5rvsn}} & z1fntw6i8wctgcl7r)
       | ({5{usm8jjd3d6kllywh9w6}} & sooa2hj7jwt64i)
       | ({5{wqwc2zh6986p0sdox}}  & w7tuyx3s7209e)
       | ({5{w663a70cvxnae9fzz}}  & wc5_xepdh0nvxo)
       | ({5{itidxzq9m2o2306pyw077}}  & j4x2ke88_rem8083g)
       | ({5{vl183kzeu77tapzyno}}  & e_sgv6k4y4pmgw89)
       ;

  assign h_3trq2o2w5gb = 
         ({5{ajcak8n6efgb0a7 }} & r8qjp6txwnbzt)
       | ({5{emvc9gbmzqk07ivf8bbc }} & cvbuf0xszkg8z2t)
       | ({5{edbnrxdg88apcxf9_wz}} & g203zwhpqmo7)
       | ({5{io39eu_nclgfwg1dh4eq4}} & tvzetpi1oen5ik)
       | ({5{x8wzvkf7gc6hluh4hx}}  & c1lj39gyj2y)
       | ({5{tb6dx9vbazjt_ikq5}}  & e9ak1p3yk1_1)
       | ({5{brrszlfkyivox7jern}}  & d0cjbhhdw6oe)
       | ({5{tlncpd0m_kefu0aje}}  & s5izacjghu1)
       ;


  wire r0g29vl2l15pr0c5y = gkfxs8wvvzhw35g2w
                 
                 | fklgk6eyb2vd8   
                 | zfotdct2of6_kc  
                 | k1oqlvc677n04h94z31 
                 | wean5xmif_myv  
                 | qzptr55gc1d815k 
                 | fouln9y77frzodomf   
                 | ot7hpozxj594mxo0o8  
                 | q9uit_5jup8pgp6l 
                 | hked2y47eglmii  
                 | utvej5knrsiltp5b    
                 | o0rfcptm6iob1mej    
                 | z3kk91ocqzu25 
                 | tv4hqiny5afky9w
                 | vwmbmpalhwfnoi_0g
                 | s_6vyiuywqqrd9say
                 | k7c8gfhghnfklxr2
                 | we6wj_afzuesr1zwnl
                 | jzbjl5cnc_hb5hixv
                 | qusz_xa0ku_toij493
                 | bi0wblozr4jb8yf4
                 ;

  wire ie85o8yuqac_w = fklgk6eyb2vd8   
                     | zfotdct2of6_kc  
                     | k1oqlvc677n04h94z31 
                     | wean5xmif_myv  
                     | qzptr55gc1d815k 
                     | fouln9y77frzodomf   
                     | ot7hpozxj594mxo0o8  
                     | q9uit_5jup8pgp6l 
                     | hked2y47eglmii  
                     | utvej5knrsiltp5b
                     | we6wj_afzuesr1zwnl
                     | jzbjl5cnc_hb5hixv
                     | qusz_xa0ku_toij493
                     | bi0wblozr4jb8yf4
                        ;   


  wire vw9hu_0ki = r0g29vl2l15pr0c5y
                 ;


  wire cod__ro1xnfzpp = ie85o8yuqac_w
                 ;













  assign rig48lgqgq8oxt = vlfahv69 ? 
                            (
                          u_mgu2iomgss4kbb5q ? 5'd2 :
                          no5vijin9fx5kyxd3lop2wg4d ? 5'd2 :
                            ga71__f5g1[5-1:0]
                            )
                            : u2apzx0s0_ms;

  assign zaub9z0lm4s93y = vlfahv69 ? 
                            (
							aihiftly[5-1:0]
							)
							: cyoz2x_qbs1p;

  
  
  
  
  assign j_69hsshtbv  = isxv0tqhyam   ? adjmfzwj55ej [5-1:0] : 
                       r5qet1mocbtcig  ? adjmfzwj55ej [5-1:0] : 
                       tx04m_rvbl9sow ? fd7uuv9az[5-1:0] : 
                       5'b0; 







  assign kd6v2vk601xpnm  = vlfahv69 ? 
                            (
							adjmfzwj55ej [5-1:0] 
							)
							: h_3trq2o2w5gb ;



   
   
   
   
   
   
   
   
   

  assign wib8hsb4py2v2tg_     = sbyhjyyw1 | gx2n0dmy9 
                         | iy0t317_b18b1 | qdqvpvjvmba ;
  assign rjob9x0q8su7ed2i    = an_cjmmfv | yxd3c1kl5vo15 
                         | wf8o8lzblge | pfeg45fn01up;
  wire c8ozh5_4o07          = wib8hsb4py2v2tg_
                         | rjob9x0q8su7ed2i;

  assign g_o2wra9n9s         = t6u2o2tra | c8ozh5_4o07;

  
  
  wire ar1cmuouyh1 = hschwo70vh36y | bx5js_t0gcoh8 | y1x6fpss6_6 | hh5fb5xzanf14 | hh5s1lrugs7 | wcsiqmn9v7po
               | c8ozh5_4o07
               ;
  assign m05tjqf24b1fabuu0e = rnx27onf2lbe & 
                            ( b7nkstim3k   
                            | cdlm5zrwv  
                            | ar1cmuouyh1) 
                            ;



  wire b3_j_0uzawl4fqhs6 = c8ozh5_4o07 & y37z_dzbgh;  
  wire a4hwlysrb9k5o37 = c8ozh5_4o07 & rfxb0v1yejd7l;
  wire dyw44w8jyc2ky0629zh;

  wire [5-1:0] njp6apzwktb8b6wm641 = u2apzx0s0_ms;
  wire [5-1:0] edfzs8oj_2g75isz = cyoz2x_qbs1p;
  wire [5-1:0] mcwlcrcptl761luzw5  = h_3trq2o2w5gb ;

  wire h8xbg9ob5pg5n_n5 = 1'b0;
  wire [5-1:0] udmsy586rsyu5j09u0 = 5'b0;

  wire fufjdaoqszpwah561178; 

  
  wire xpnihwic7a27noexvq = t6u2o2tra;
                    
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  wire j50bt7tjt4wz8hkuvv = t6u2o2tra &
                (
                 (~hschwo70vh36y)
               & (~y1x6fpss6_6)
               & (~o4tc3g036bgoap)
               & (~cbru05_q5bm7)
               & (~dywxta8oxdnj1q9i0d)
               & (~zqz28qv7052ajkf7)
               & (~iz_sm_7y_ixfw1btmz)
               & (~uz6maeeehzsn6uzwxk)
               & (~tnkhekmenrbyvq)
               & (~gsqes4kpzyh7s4)
               & (~i_oja_fou8xg9_)
               & (~jz2t1e591yva8m5)
               & (~th_rx8vbgu0ydrx)
               & (~glahkq0rwcrj086j7k1j)
               & (~nu4l8_3i80k9r9huos)
               & (~wjhbw3uh3oljyutu2gel)
               & (~hx05sow34f5nxv)
               & (~iboby_h0cqqucgnxw)
               & (~q1mnx00q446iezuqt)
               & (~bvcgz8q5ffa32w7)
               & (~knqkb_9b7915rg)
               & (~jlez7xntekztmffn06)
               & (~gkj8ltdpe4tcqini4h)
               & (~va7j9_tx3li0xd)
               & (~l6qpfpq3ro_9gr)
               & (~nxf52k3xp6im5o6p3)
               & (~u72qi7gmhj37d_h5c)
               & (~tr03xi8fsjspsc)
                 );

  
  wire rhttudaoog18_uuoooxeob = t6u2o2tra & (qwppxd4zz
                                    | wh7hmrmzlb 
                                    | eueft5qh43m7e
                                    | jn7op2_63ozfv);

    
    
  wire [5-1:0] k4_jx9ixctuib2g1b  = pq5pe3yehrqxr[31:27];
  assign jc4yg1pkylr2gonwcd = vlfahv69 ? ga71__f5g1[5-1:0] : njp6apzwktb8b6wm641;
  assign nd3cgvec1pogf2 = vlfahv69 ? aihiftly[5-1:0] : edfzs8oj_2g75isz;
  assign f7crsrzernrwgmepy = vlfahv69 ? k4_jx9ixctuib2g1b[5-1:0] : udmsy586rsyu5j09u0;
  assign pw085ct76po3c  = vlfahv69 ? adjmfzwj55ej [5-1:0] : mcwlcrcptl761luzw5 ;
  
  
  
  
  
  
  
    
    
    
    
    
    
    
    
    
    
    
  
  
    
    
  
  
    
    
    
  
  
    
    

  wire l4p2yfrqb9vqu331  = t6u2o2tra & (
                             (~glv8ztvxphxctm)
                           & (~kvnjxxg7anei8786qg)
                           & (~dywxta8oxdnj1q9i0d )
                           & (~zqz28qv7052ajkf7)
                           & (~i_oja_fou8xg9_ )
                           & (~jz2t1e591yva8m5)
                           & (~nu4l8_3i80k9r9huos )
                           & (~wjhbw3uh3oljyutu2gel)
                           & (~q1mnx00q446iezuqt )
                           & (~bvcgz8q5ffa32w7)
                           & (~nxf52k3xp6im5o6p3)
                           & (~tr03xi8fsjspsc)
                           );
  wire brx6nla_mtrays  = t6u2o2tra;
  wire j23vj00z182h  = t6u2o2tra;
  wire oj48f6biuilerfy   = t6u2o2tra & (
                             (~iz_sm_7y_ixfw1btmz )
                           & (~uz6maeeehzsn6uzwxk)
                           & (~th_rx8vbgu0ydrx )
                           & (~glahkq0rwcrj086j7k1j)
                           & (~hx05sow34f5nxv )
                           & (~iboby_h0cqqucgnxw)
                           & (~knqkb_9b7915rg )
                           & (~jlez7xntekztmffn06)
                           & (~gkj8ltdpe4tcqini4h)
                           & (~va7j9_tx3li0xd)
                           & (~qfgkmomxjwhe)
                           & (~v3he_44ycy65)
                           & (~h5gjvo_bpoph5i)
                           & (~ns2ccb8p4kf3o)
                           & (~wy5oiwkuovruvc)
                           & (~mtnmu5bzb5z9)
                           & (~u72qi7gmhj37d_h5c)
                           & (~l6qpfpq3ro_9gr)
                           & (~u72qi7gmhj37d_h5c)
                           );
  
  
  
  wire phs3h9_sv3ea6q  = c8ozh5_4o07 & (~wib8hsb4py2v2tg_) & (~rjob9x0q8su7ed2i);
  wire mn5von2vdgtowoe  = c8ozh5_4o07;
  wire cbfgecuirt4z_t  = c8ozh5_4o07;
  wire dvzltftlrzgl   = c8ozh5_4o07;


  assign dyw44w8jyc2ky0629zh  = c8ozh5_4o07 & yjigfdj36u7d3yg &
                         (~((~dvzltftlrzgl) & (h_3trq2o2w5gb == 5'b0))) 
                         ;

  
  
  
  assign fufjdaoqszpwah561178 = t6u2o2tra &
                    (
                      (~kvnjxxg7anei8786qg)
                    ) &
                    (~((~oj48f6biuilerfy) & adw7hffbin))
                    ;

  assign nykwng_3anppxi  = vlfahv69 ? (xpnihwic7a27noexvq) : (b3_j_0uzawl4fqhs6);
  assign shpynlimbt55rj4  = vlfahv69 ? (j50bt7tjt4wz8hkuvv) : (a4hwlysrb9k5o37);
  assign jycwup76klyed6d2  = vlfahv69 ? (rhttudaoog18_uuoooxeob) : (h8xbg9ob5pg5n_n5);
  assign i7pubsxfsb4uys  = vlfahv69 ? (fufjdaoqszpwah561178) : (dyw44w8jyc2ky0629zh );
  assign fgm5kq4y725x6yylw = vlfahv69 ? (l4p2yfrqb9vqu331) : (phs3h9_sv3ea6q);
  assign awld9ngcypgfxa = vlfahv69 ? (brx6nla_mtrays) : (mn5von2vdgtowoe);
  assign v5m66onlnmxeejfhn = vlfahv69 ? (j23vj00z182h) : (cbfgecuirt4z_t);
  assign kfz3mojvfh2fsfd  = vlfahv69 ? (oj48f6biuilerfy ) : (dvzltftlrzgl );

  assign sb8ax73d3ud = vlfahv69 ? hegurso01yv4i : (y37z_dzbgh & (~(u2apzx0s0_ms == 5'b0))); 
  assign f9_w27gbcq__ = vlfahv69 ? hgjytyuf89rdi : (rfxb0v1yejd7l & (~(cyoz2x_qbs1p == 5'b0)));
  assign iq9sj_i8z1k712   =  chso39421msvbkl9a; 
  assign b6cv9yeaga7hf = vlfahv69 ? bqywdsjnr1r6icc0 : (yjigfdj36u7d3yg & (~(h_3trq2o2w5gb  == 5'b0)));

  assign mg0onistbzu9ys = (rig48lgqgq8oxt == 5'b0);
  assign g3btysb7vvv = (zaub9z0lm4s93y == 5'b0);
  assign yjgkn7vcv = (j_69hsshtbv == 5'b0);  

  wire hqxuxwgpn_xbzk1;














      
  assign hqxuxwgpn_xbzk1 = 1'b0;

  assign nnng_p6632p = vlfahv69;

  assign bdhv0j4zhtx9nxmz = 
                     ({64{e_qxxtaevvw | ei1me6y0     }} & q6dj3cn7jeic88g0ok)
                   | ({64{lr08s8a1cosklchm4m      }} & onxwi3lt3vee8230ahq9)
                   | ({64{tez8bez5l4r | zh62ppn61_4yw4 }} & xoxse1yov4vm01rl)
                   | ({64{h20g0j2jt              }} & qytu41_x5zlegr)
                   | ({64{sa6649too5v5             }} & hf_ehpaimuswmut)
                   | ({64{o6soq_mfr7s9lh51rhx5      }} & x8lnalqbfmpei)
                   ;

  assign ng_pudjzgnamv0es = vlfahv69 ? ga71__f5g1[5-1:0] : ag9ylluguwcr[5-1:0]; 


  assign fqizcmmfg   = u2k4dyp52s_m;
  assign tbuacpjktio   = djvj1e_;
  assign ciftsjs2bvaxns   = bktu0z1mk56;


  assign dwci8hbxok739 = v91kaxeokzy6fv5 | g0rwtpabeiisocfnwg
                       | (r773brf2qafg123x)
                       | (ebxkh3mj83gh00a86o_rb)
                       | (r1pa5yctc1vd7e650n)
                       | (plr5quy6x6fvmq27ye)
                       ; 

  assign fpwql5ik7_sp0 = 
            (ctcwxdialrasri5u6guy) 
          | (hqxuxwgpn_xbzk1) 
          | (kg80830otj0fcd2qp2u90)
          | (epmy5pkue90oo6im57xozi)
          | (oa000fsbi9vz2933)
          | (x9cbta8yo_b811qozvyp0tqoa)
          | (g0rwtpabeiisocfnwg)
          | (v91kaxeokzy6fv5)
          | (r773brf2qafg123x)
          | (ebxkh3mj83gh00a86o_rb)
          | (r1pa5yctc1vd7e650n)
          | (plr5quy6x6fvmq27ye)
          | rb8rv_jwet5lap0p
          | w15cfmvs_rdfsulo
          | elg6c3h_r04v5e71
          | (ww_v_rhq1pd2_fg)
          | k2shv0srgu0krb8ve 
          | oo_r3ir9zo8z6zvfbo
          | m05tjqf24b1fabuu0e
          | qzjna_8yrjwqibq75b9s 
          | ir80nlzybrgunagd7j 
          | piay0j_yijhago5y 




          | wa2rqb81bsgzs2g9adv
          | (~wri2knqd9wtnw);

  wire d3e2e1oz1q = 1'b0;


  assign zk9uk90j08ogqpn[0] = 1'b0;

  assign zk9uk90j08ogqpn[1] = 1'b1;

  assign zk9uk90j08ogqpn[2] = 1'b1;

  assign zk9uk90j08ogqpn[3] = v7s5fo07nb5 & a51ngszcxd19m[5:5];

  assign zk9uk90j08ogqpn[4] = v7s5fo07nb5 & a51ngszcxd19m[6:6]; 

  assign zk9uk90j08ogqpn[5] = v7s5fo07nb5 & a51ngszcxd19m[11:11]; 

  assign zk9uk90j08ogqpn[6] = sm_lqinid6ej;

  assign zk9uk90j08ogqpn[7] = hqkcyoh04f5d5j;

  assign zk9uk90j08ogqpn[8] = j_ku88w81rg;

  assign zk9uk90j08ogqpn[9] = j_ku88w81rg;

  assign zk9uk90j08ogqpn[10] = o8rwk067;



  assign zk9uk90j08ogqpn[11] = r1on2k03r;






  wire fo1wd_wpluhuucji = (rig48lgqgq8oxt == 5'd1);
  wire b3wi4y0jobpbh_bhc3rl = (rig48lgqgq8oxt == 5'd5);
  wire qurxq4mqvhmg4q = (kd6v2vk601xpnm == 5'd1);
  wire ujkxu7tcwu6bne8 = (kd6v2vk601xpnm == 5'd5);
  wire v9yeadvpvxx5m0w4i4swx = fo1wd_wpluhuucji | b3wi4y0jobpbh_bhc3rl;
  wire m8emmeleqvsylkfd0ip = qurxq4mqvhmg4q | ujkxu7tcwu6bne8;
  assign zk9uk90j08ogqpn[12] = r1on2k03r & (bdhv0j4zhtx9nxmz == 64'b0) & (
                             ((~m8emmeleqvsylkfd0ip) & v9yeadvpvxx5m0w4i4swx)
                           | (qurxq4mqvhmg4q & b3wi4y0jobpbh_bhc3rl)
                           | (ujkxu7tcwu6bne8 & fo1wd_wpluhuucji)
                          );


  assign zk9uk90j08ogqpn[13] = r1on2k03r | o8rwk067 | j_ku88w81rg;

  assign zk9uk90j08ogqpn[14] = 
                             1'b0
                             ;

  assign zk9uk90j08ogqpn[15] = s0aynip0upf & (t9xs6bqphiru | ls1dudpc);

  assign zk9uk90j08ogqpn[16] = s0aynip0upf & (tzjssx03b | kt04okvuth | cni2453cuofb | kq9gup8pu2);

  assign zk9uk90j08ogqpn[17] = glv8ztvxphxctm;

  assign zk9uk90j08ogqpn[18] = kvnjxxg7anei8786qg;

  assign zk9uk90j08ogqpn[19] = fz4uie4yxvn5 | snxdp3tvw7a | knc4udhhcbv | vou4ap3g4kukvz7a;

  assign zk9uk90j08ogqpn[20] = x0c94xeqpc8nzim7 | ou19p6zx65a;


  assign zk9uk90j08ogqpn[21] = t6u2o2tra & (qwppxd4zz | wh7hmrmzlb | eueft5qh43m7e | jn7op2_63ozfv);


  assign zk9uk90j08ogqpn[22] = (kzyiyt0xi8d | o4tc3g036bgoap | lz1544702tkg0u | cbru05_q5bm7);

  assign zk9uk90j08ogqpn[23] = t6u2o2tra & (~(|zk9uk90j08ogqpn[22:17]));
  assign zk9uk90j08ogqpn[31:24] = 8'b0;


endmodule                                      



module qh5_zkb1tn0pxt6hr3yb # (
  parameter onr7l = 32,
  parameter d5y59uh9zri = {onr7l{1'b0}}
)(

  input               abwn, 
  input      [onr7l-1:0] q461tw,
  output     [onr7l-1:0] p4dxkq4k,

  input               gf33atgy,
  input               ru_wi
);

reg [onr7l-1:0] nkvgr6w73w;

always @(posedge gf33atgy or negedge ru_wi)
begin : y37z8h3v53a3
  if (ru_wi == 1'b0)
    nkvgr6w73w <= d5y59uh9zri;
  else if (abwn == 1'b1)
    nkvgr6w73w <= q461tw;
end

assign p4dxkq4k = nkvgr6w73w;


endmodule



module sav90_q6tp_eioxey5390qd # (


  parameter tcebpmbl7g = 0,
  parameter mhdlk = 1,
  parameter onr7l = 32
) (
  input           bw6ftrau0, 
  output          eef2g8, 
  input  [onr7l-1:0] qbjvs30wtb,
  output          wqljp, 
  input           h9378, 
  output [onr7l-1:0] dqgck5s,

  input           gf33atgy,
  input           ru_wi
);

  genvar i;
  generate 

  if(mhdlk == 0) begin: kum1oxhw1b434q

      assign wqljp = bw6ftrau0;
      assign eef2g8 = h9378;
      assign dqgck5s = qbjvs30wtb;

  end
  else begin: r1f9lplxw0lya5z

      wire d35brwhbkm;
      wire xlzi7_mjg;
      wire xayqet0sd;
      wire ycgzbt;
      wire d0x7t39v;


      assign d35brwhbkm = bw6ftrau0 & eef2g8;

      assign xlzi7_mjg = wqljp & h9378;

      assign xayqet0sd = d35brwhbkm | xlzi7_mjg;
      assign d0x7t39v = d35brwhbkm | (~xlzi7_mjg);

      ux607_gnrl_dfflr #(1) hdti_6iaq (xayqet0sd, d0x7t39v, ycgzbt, gf33atgy, ru_wi);

      assign wqljp = ycgzbt;

      ux607_gnrl_dfflr #(onr7l) tn7qvilprku (d35brwhbkm, qbjvs30wtb, dqgck5s, gf33atgy, ru_wi);

      if(tcebpmbl7g == 1) begin:lvfon_zgkwp229

          assign eef2g8 = (~ycgzbt);
      end
      else begin:ulbqsqnmhe2qhizmyx

          assign eef2g8 = (~ycgzbt) | xlzi7_mjg;
      end
  end
  endgenerate


endmodule 


































module v3jar7rg0a6jqc(
  input  r5hpbriny8m67sv9e_ylgo1,
  input  dyl5g2vgrvy4mb3,





  input  vi03qlql8tkd5,


  input  p1oz3zlyx9z099ko, 
  output i7xpott8rcin, 

  input  i4ph1cg8ey91ao,

  input v367rhzcrd1qq5y,
  input m6ow3ped_b3ynpgtz,
  input po8t3bdmxflhl2,
  input acploblvq3_mum6ni,
  input d5hyfhqo_lj0prgy,
  input pf_xchk7690b64ux,
  input [48-1:0]  nog5k2tkaj_,

  input kshl17el0r504ln0s0,


  input  so8hgqibdpmm,
  input  jyc3e55o28bdrj7ce,
  input  jjab0msl5gufous,
  input  y4er8_lympr8x7vr4,
  input  fxa5t2739h1y,
  input  ng2go_dzj8ezoh,
  input  [5-1:0] pdyldj59mo6vg0bdw,
  input  [5-1:0] dxnb4vitu85cv,
  input  [5-1:0] y0sg1fz2ziwsp,
  input  [64-1:0] xfxtnu32e4,
  input  [64-1:0] bzyabkjyg5aufwj,
  input  [64-1:0] be99yq3n56,
  input  l2t6z9zsi2w0_zq,
  input  [3-1:0] k1hmos4y13oq40h,
  input  [5-1:0] ir18j9t6197l06,
  input  [64-1:0] a1nhqrkfzavps,
  input  [31:0] d0fq7icjv8j5ogee,
  input  [64-1:0] ee8ig_qwdt,
  input  [64-1:0] kn1fenl59sz01m7vnq2em_s,
  input  [4*8-1:0] u_rd99v1d167myvqms9,
  input  yauc7c8wjjqclo3tp,
  input  [2-1:0] m_h2ikgwk1idzghe517,
  input  [9-1:0] sjpycsle28a3pm_p,
  input  vuxawlqfs_00v7_hzu3nxvoz,


  output [7:0] kbdkmakcambtuegb3yt,
  input  [7:0] u9fj6h2fgqotisf,
  input  [2:0] z2kxp5om4aw87pz8o18n1z6h,
  output [2:0] i6zm27hf33zy3u5g9qudq24sqm285,

  input  hyt20f5h_uwl66fhu4_,
  input  qmscup3rxdd9panua6h,
  input  odgwr675x09tn ,
  input  lzddtts2zym6c0cpur ,
  input  i11dangz7fq7x35giy ,
  input  zyh78crm605f5vguk,
  input  p_cayjjoaokcjaec,
  input  ciy8of6we8nbld  ,
  input  dcpzocokm__mx7iua  ,
  input  isem4fqob1u88i  ,
  input  rqmodrsg4hiv3yd ,
  input  e6dhhsva7_jc3yex ,
  input  m01780lmcvgmej7gv  ,
  input  vmc4uk3dtr_i3b6a1ojb,

  input ssbpxp6oebc9u,
  input mp__ij57saap5pzjguck,
  input bzxq5cchssdayz9w,
  input j35b4l1vciavqz_c8d,
  input q3fqrzgv4ce7343pb4,
  input [5-1:0] lou99zfk5t2fgui5tdozk,
  input [5-1:0] vx_07j3zzi0_m3lyq2tj,
  input [5-1:0] zo2kgt18lgbbaee80oq,
  input [5-1:0] cez5fjfkhrstof7vn,
  input woaibn5hs0f9zh9obi,
  input rczetx728pgbbuyhj,
  input l4y91rsecb8o3de_m,
  input i90ggmn3seqiequ3ikr,
  input  [64-1:0] dg8l11o4gz7pp4nz6q,
  input  [64-1:0] l_w_v2dy7wxfnyy_ka5,
  input  [64-1:0] zrckh33wcln3qe0gwm,

  input  glf9eqlzf6ocu2fgv_jen,
  output fn921s9pkxbuyodk3cs,



  output d3le01r9nrj56s4d, 
  input  awd7cj8qhsnpdq2i,

  input  mhnv1zj1t2xbsvq6pgtez4d,
  input  h76iv7j9x_gukyjc7q75qp_kags,

  output [64-1:0] fssz5redtt2z0j3bm,
  output [64-1:0] vahtdoye9yd23j,
  output [64-1:0] tc85_x5h95y20zrlyv5,
  output [3-1:0] cqiq85nw82tognls5,
  output e8htsab8ol_n9_vmg55h,
  output v8h7kn3z48bhc41oj0m,
  output [5-1:0] s_ngsncbxs5sazdn09m2,
  output [64-1:0] tml6nm8cttakxkfl21,
  output [31:0] qjdagljhhzu7oqkdf8dt,
  output [64-1:0] pj2f1w77r_add,
  output [64-1:0] euzjqpru0y77ampkkzy_xt,
  output [4*8-1:0] mizeob9j8ozttr2_5f1bf4zfgw0j,
  output hl3g_tq2rbkqa9ohkpb,
  output [2-1:0] zrnrmtty0nzt9spsnhdcm1fcb,
  output [9-1:0]  m9w2x58qenx6t_2bi2,
  output sw9yrs02t82mjdszv19xlcnijsm,
  output [4-1:0] ta29h0x4_ymr6ur6mk04,
  output lgm4pk95gcg3msfburvh,
  output r9xo5zxa6yk5sahklgriapc,
  output qhr7po23q4sobg2liu8pg ,
  output fat5whs4wafix5rmfhm4837957 ,
  output wtormxdkxhzy97pmh ,
  output dskiex0swz5vysk4mc5 ,
  output w313qpi6k9c_3uaxaj_ew ,
  output hzx0lxqvh33f51vttk0y  ,
  output vzwsikmnhz1uumkd9  ,
  output vfq4rm5ouxjqvse7  ,
  output p0q6b5s2pyhh9h5qc724n ,
  output m755tv316f55fgbeul39qh,
  output bvwm3a9jzm7y_sjdaeqvzzvxeg,



  input  hwu6b9ql3l7sw43wkk0lg,
  input  a4rzfgrj8wj0hf3kl4wtn,
  input  dp3lxnqfh_zuqs0qfwzb8,
  input  [4-1:0] g5uxvsehmtgyorg3wb ,
  output jya9awf7h3oxy2ame3,
  input  gjbc27bxx6tkh_1w1,
  output i9h3d3za76przvk_l70p,
  output euc_83pmnhwvr32xx,
  output o2psmcgly2h0shgva5,
  output f9fubli1q2_q74eh ,

  output rev7x95ee0q6067 ,
  output bpr67a65mrtg6l5byk3 ,
  output qe_d8g8bvqcuzvaepz ,
  output l56hg65h6fdq8htrj6gb ,


  output hrlh00uvgxvc0v3fhap ,
  output xnnfhu8lpo04_jagyvmf ,
  output keve1s8kiyssv8a ,

  output [5-1:0] fnkzuyagjhoinc95_,
  output [5-1:0] x70ugsspg9qc0ccmj,
  output [5-1:0] bhpc3d1wahnkux0bil5x,
  output [5-1:0] wtrlpn7minfboagr ,


  output feq1g7m2cy1erl,

  input  gf33atgy,
  input  ru_wi
  );

  wire zhf3ql_4fi_c5_b1;




  assign zhf3ql_4fi_c5_b1 = 1'b0;

  assign feq1g7m2cy1erl = 1'b0;









  wire ac3235afm = acploblvq3_mum6ni;
  wire h16aj5yf = d5hyfhqo_lj0prgy;

  wire obeilvz6aywpv3jnunz = h76iv7j9x_gukyjc7q75qp_kags;
  wire u9ys3fhcgd7kbaxni5ea = mhnv1zj1t2xbsvq6pgtez4d;


  wire zymbxusz8g0f4apj7   = po8t3bdmxflhl2 &
                               ( nog5k2tkaj_ [20:20] | nog5k2tkaj_ [21:21]);   
  wire ljzvtkybvc4         = po8t3bdmxflhl2 & nog5k2tkaj_ [21:21];   
  wire okhq1zhvfjuf         = po8t3bdmxflhl2 & nog5k2tkaj_ [22:22]; 

  wire ckx7zudt_jkvcyxrqbh_6wyl8_7v = zymbxusz8g0f4apj7 | okhq1zhvfjuf;




  wire w860ns6z_bj6yyaj; 

  wire   j746sidtcglv5f5n = awd7cj8qhsnpdq2i;


  assign d3le01r9nrj56s4d = w860ns6z_bj6yyaj; 

































  wire fu959zi =  ((hwu6b9ql3l7sw43wkk0lg)   |
                   (a4rzfgrj8wj0hf3kl4wtn)   |
                   (dp3lxnqfh_zuqs0qfwzb8)
				   ); 


















  wire cm2y65s0 = (
                    1'b0
				  ); 

  wire fqieg3m = fu959zi | cm2y65s0; 

  wire cztyzemcgla7e0ev = pf_xchk7690b64ux;


  wire uoq13ng8ai8cg = kshl17el0r504ln0s0;















  wire uoq92ktpn3xml4sibfj = 







               & (cztyzemcgla7e0ev ? vi03qlql8tkd5 : 1'b1) 
               & (uoq13ng8ai8cg ? vi03qlql8tkd5 : 1'b1) 
               & ((ckx7zudt_jkvcyxrqbh_6wyl8_7v) ? (vi03qlql8tkd5 & (~r5hpbriny8m67sv9e_ylgo1)) : 1'b1)

               & (~zhf3ql_4fi_c5_b1)
               & (~feq1g7m2cy1erl)


               
               
               & gjbc27bxx6tkh_1w1 
               ;

  assign w860ns6z_bj6yyaj = uoq92ktpn3xml4sibfj & p1oz3zlyx9z099ko; 
  assign i7xpott8rcin     = uoq92ktpn3xml4sibfj & j746sidtcglv5f5n; 






  wire [64-1:0] l0mrvs75tc02qy = {{64-64{1'b0}},dg8l11o4gz7pp4nz6q};
  wire [64-1:0] wv8yw1ke55mr = {{64-64{1'b0}},l_w_v2dy7wxfnyy_ka5};
  wire [64-1:0] coq3ctgsd9iar8 = {{64-64{1'b0}},zrckh33wcln3qe0gwm};

  wire [64-1:0] qpscc8xem = {{64-64{1'b0}},(xfxtnu32e4 & {64{~so8hgqibdpmm}})};
  wire [64-1:0] u3wdadynlf = {{64-64{1'b0}},(bzyabkjyg5aufwj & {64{~jyc3e55o28bdrj7ce}})};
  wire [64-1:0] igvq6tvqkm = {{64-64{1'b0}},(be99yq3n56 & {64{~jjab0msl5gufous}})};

  wire [64-1:0] kb70bgh44hh7uig8d = i9h3d3za76przvk_l70p ? l0mrvs75tc02qy : qpscc8xem ;
  wire [64-1:0] lrgxvtpcvkq20zjin5 = euc_83pmnhwvr32xx ? wv8yw1ke55mr : u3wdadynlf ;
  wire [64-1:0] pvkagzonx0zz8b7on = o2psmcgly2h0shgva5 ? coq3ctgsd9iar8 :  
                                                        igvq6tvqkm
                                              ;









  assign fssz5redtt2z0j3bm   = kb70bgh44hh7uig8d;
  assign vahtdoye9yd23j   = lrgxvtpcvkq20zjin5;
  assign tc85_x5h95y20zrlyv5   = pvkagzonx0zz8b7on;
  assign cqiq85nw82tognls5 = k1hmos4y13oq40h;
  assign e8htsab8ol_n9_vmg55h = f9fubli1q2_q74eh & l56hg65h6fdq8htrj6gb; 
  assign v8h7kn3z48bhc41oj0m = l2t6z9zsi2w0_zq;
  assign s_ngsncbxs5sazdn09m2 = ir18j9t6197l06;
  assign fn921s9pkxbuyodk3cs   = glf9eqlzf6ocu2fgv_jen;





  assign jya9awf7h3oxy2ame3 = d3le01r9nrj56s4d & awd7cj8qhsnpdq2i; 


  assign tml6nm8cttakxkfl21  = a1nhqrkfzavps;
  assign pj2f1w77r_add   = ee8ig_qwdt;
  assign euzjqpru0y77ampkkzy_xt = kn1fenl59sz01m7vnq2em_s;
  assign sw9yrs02t82mjdszv19xlcnijsm = vuxawlqfs_00v7_hzu3nxvoz;
  assign mizeob9j8ozttr2_5f1bf4zfgw0j = u_rd99v1d167myvqms9;
  assign hl3g_tq2rbkqa9ohkpb = yauc7c8wjjqclo3tp;
  assign zrnrmtty0nzt9spsnhdcm1fcb = m_h2ikgwk1idzghe517;
  assign m9w2x58qenx6t_2bi2 = sjpycsle28a3pm_p;

  assign kbdkmakcambtuegb3yt = u9fj6h2fgqotisf;
  assign i6zm27hf33zy3u5g9qudq24sqm285 = z2kxp5om4aw87pz8o18n1z6h;
  assign ta29h0x4_ymr6ur6mk04 = g5uxvsehmtgyorg3wb;
  assign lgm4pk95gcg3msfburvh= hyt20f5h_uwl66fhu4_;
  assign r9xo5zxa6yk5sahklgriapc= qmscup3rxdd9panua6h;
  assign qhr7po23q4sobg2liu8pg = odgwr675x09tn;
  assign fat5whs4wafix5rmfhm4837957 = lzddtts2zym6c0cpur;
  assign wtormxdkxhzy97pmh = i11dangz7fq7x35giy;
  assign dskiex0swz5vysk4mc5 = zyh78crm605f5vguk;
  assign w313qpi6k9c_3uaxaj_ew = p_cayjjoaokcjaec;
  assign hzx0lxqvh33f51vttk0y  = ciy8of6we8nbld   ;
  assign vzwsikmnhz1uumkd9  = dcpzocokm__mx7iua   ;
  assign vfq4rm5ouxjqvse7  = isem4fqob1u88i   ;
  assign p0q6b5s2pyhh9h5qc724n = rqmodrsg4hiv3yd  ;
  assign m755tv316f55fgbeul39qh   = m01780lmcvgmej7gv;
  assign bvwm3a9jzm7y_sjdaeqvzzvxeg = vmc4uk3dtr_i3b6a1ojb;

  assign i9h3d3za76przvk_l70p = ssbpxp6oebc9u ? (mp__ij57saap5pzjguck & woaibn5hs0f9zh9obi) : 1'b0;
  assign euc_83pmnhwvr32xx = ssbpxp6oebc9u ? (bzxq5cchssdayz9w & rczetx728pgbbuyhj) : 1'b0;
  assign o2psmcgly2h0shgva5 = ssbpxp6oebc9u ? (j35b4l1vciavqz_c8d & l4y91rsecb8o3de_m) : 1'b0;
  assign f9fubli1q2_q74eh  = ssbpxp6oebc9u ? (q3fqrzgv4ce7343pb4 & i90ggmn3seqiequ3ikr ) : 1'b0;

  assign rev7x95ee0q6067  = ssbpxp6oebc9u ? mp__ij57saap5pzjguck : y4er8_lympr8x7vr4;
  assign bpr67a65mrtg6l5byk3  = ssbpxp6oebc9u ? bzxq5cchssdayz9w : fxa5t2739h1y;
  assign qe_d8g8bvqcuzvaepz  = ssbpxp6oebc9u ? j35b4l1vciavqz_c8d :
                                                          ng2go_dzj8ezoh 
                                                         ;
  assign l56hg65h6fdq8htrj6gb  = ssbpxp6oebc9u ? q3fqrzgv4ce7343pb4 : l2t6z9zsi2w0_zq;

  assign hrlh00uvgxvc0v3fhap  = ssbpxp6oebc9u ? 1'b0 : so8hgqibdpmm;
  assign xnnfhu8lpo04_jagyvmf  = ssbpxp6oebc9u ? 1'b0 : jyc3e55o28bdrj7ce;
  assign keve1s8kiyssv8a  = ssbpxp6oebc9u ? 1'b0 :
                                                 jjab0msl5gufous 
                                             ;


  assign fnkzuyagjhoinc95_ = ssbpxp6oebc9u ? lou99zfk5t2fgui5tdozk : pdyldj59mo6vg0bdw;
  assign x70ugsspg9qc0ccmj = ssbpxp6oebc9u ? vx_07j3zzi0_m3lyq2tj : dxnb4vitu85cv;
  assign bhpc3d1wahnkux0bil5x = ssbpxp6oebc9u ? zo2kgt18lgbbaee80oq : y0sg1fz2ziwsp;
  assign wtrlpn7minfboagr  = ssbpxp6oebc9u ? cez5fjfkhrstof7vn  : ir18j9t6197l06;



  assign qjdagljhhzu7oqkdf8dt = d0fq7icjv8j5ogee; 



endmodule                                      





`define UX607_EXU_DIVCORE__V


module jvwuov7by1m8upbjlyy6 (
  input [68-1:0] rydw,
  input [68-1:0] d4y,
  input [68-1:0] iev4j_o4,
  input [68-1:0] hfl_1crp,
  input [68-1:0] h891r,
  input [68-1:0] m48h,
  input [68-1:0] r04h,
  input k2xz1iocfj4qk7btop,
  
  output [68-1:0] kktrbu07,
  output [68-1:0] kf9hl8c_,
  output [68-1:0] spfqyly64 ,
  output [68-1:0] dqm4y5o,
  output [68-1:0] tzwq6o86 
  );

wire [68-1:0] ctoy95b;
wire [68-1:0] zlq70vuuuc;
wire [68-1:0] ujdzwwros_3b ;
wire [68-1:0] olgpxn;
wire [68-1:0] vdmf0obdru6b;

wire ktu7z7eeks17;
wire oxt4ewm09j ;
wire p5l63dwt7156pi;

qp2s59tux3j91cdjqs bwajrce_x9amgczb8w362txq7h(
  .rydw     (rydw),
  .d4y     (d4y),
  .w0m_yvp2sos8e(ktu7z7eeks17),
  .dtgamdbpa4gj (oxt4ewm09j ),
  .ysl1y4xf1(p5l63dwt7156pi)
);

assign ujdzwwros_3b[68-1-1:0] = h891r[68-1:1] ;
assign ujdzwwros_3b[68-1] = 1'b1 ;

c2dm5oqn6257o319rma1kr9 p1cgh45s12e714v00acvr85vmw56(
  .rydw     (rydw),
  .d4y     (d4y),
  .iev4j_o4 (iev4j_o4),
  .hfl_1crp (hfl_1crp),
  .ysl1y4xf1(p5l63dwt7156pi),
  .w0m_yvp2sos8e(ktu7z7eeks17),
  .dtgamdbpa4gj (oxt4ewm09j ),
  .xphx    (ctoy95b),
  .fap75    (zlq70vuuuc)
);

assign olgpxn  = (p5l63dwt7156pi ? r04h : m48h) & ujdzwwros_3b | ~{68{oxt4ewm09j}} & ~ujdzwwros_3b ;
assign vdmf0obdru6b = (ktu7z7eeks17 ? m48h : r04h) & ujdzwwros_3b | {68{oxt4ewm09j}} & ~ujdzwwros_3b ;

wire [68-1:0] r5utfvc7oz     =ctoy95b;
wire [68-1:0] vqxjyefxtk     =zlq70vuuuc;
wire [68-1:0] ptl5g3zjau =iev4j_o4;
wire [68-1:0] ptvzkd3c5gfz85 =hfl_1crp;
wire [68-1:0] iily74b8    =ujdzwwros_3b;
wire [68-1:0] idpqk     =olgpxn;
wire [68-1:0] vpvwojcah    =vdmf0obdru6b;

wire [68-1:0] iy7_96w4xsmu7xh;
wire [68-1:0] rude3zls82mq;
c2dm5oqn6257o319rma1kr9 ltfzoc5jxilrl4i1_1dpfan_xq1j0(
  .rydw     (rydw),
  .d4y     (d4y),
  .iev4j_o4 (iev4j_o4),
  .hfl_1crp (hfl_1crp),
  .ysl1y4xf1(1'b0),
  .w0m_yvp2sos8e(1'b0),
  .dtgamdbpa4gj (1'b1 ),
  .xphx    (iy7_96w4xsmu7xh),
  .fap75    (rude3zls82mq)
);

wire y022y5lgu5q5z_i;
wire tqt6kzwmx2e3h2 ;
wire y2hpqatjf4b06o47va;

qp2s59tux3j91cdjqs urg8v842scsuz_5ktdmq0o2z(
  .rydw     (iy7_96w4xsmu7xh),
  .d4y     (rude3zls82mq),
  .w0m_yvp2sos8e(y022y5lgu5q5z_i),
  .dtgamdbpa4gj (tqt6kzwmx2e3h2 ),
  .ysl1y4xf1(y2hpqatjf4b06o47va)
);

wire [68-1:0] z1f2orfwb02yxhy;
wire [68-1:0] hj63u9fp059ch;
c2dm5oqn6257o319rma1kr9 b0d9dp6lebs3pxu1cpqcs9n2viyf(
  .rydw     (rydw),
  .d4y     (d4y),
  .iev4j_o4 (iev4j_o4),
  .hfl_1crp (hfl_1crp),
  .ysl1y4xf1(1'b0),
  .w0m_yvp2sos8e(1'b1),
  .dtgamdbpa4gj (1'b0 ),
  .xphx    (z1f2orfwb02yxhy),
  .fap75    (hj63u9fp059ch)
);

wire wufvkpcwv_7l53;
wire ilnldo2qebgfdabgfq ;
wire zrotme_c1tv9ggx;

qp2s59tux3j91cdjqs l_hv4zym21ow5ws9kxx588(
  .rydw     (z1f2orfwb02yxhy),
  .d4y     (hj63u9fp059ch),
  .w0m_yvp2sos8e(wufvkpcwv_7l53),
  .dtgamdbpa4gj (ilnldo2qebgfdabgfq ),
  .ysl1y4xf1(zrotme_c1tv9ggx)
);

wire [68-1:0] xyoecfug3y_5s3;
wire [68-1:0] njxu97ibzwrkjyek;
c2dm5oqn6257o319rma1kr9 glccozti43ihspkqq8127vmj3yz6(
  .rydw     (rydw),
  .d4y     (d4y),
  .iev4j_o4 (iev4j_o4),
  .hfl_1crp (hfl_1crp),
  .ysl1y4xf1(1'b1),
  .w0m_yvp2sos8e(1'b0),
  .dtgamdbpa4gj (1'b0 ),
  .xphx    (xyoecfug3y_5s3),
  .fap75    (njxu97ibzwrkjyek)
);

wire uqcuak_gzilz7mrpz0;
wire nk0icy0xeofyyx1w_l ;
wire otcdnhpg8mwltf;

qp2s59tux3j91cdjqs djuuhh3zwc97c6u6q6r9hsoosnq(
  .rydw     (xyoecfug3y_5s3),
  .d4y     (njxu97ibzwrkjyek),
  .w0m_yvp2sos8e(uqcuak_gzilz7mrpz0),
  .dtgamdbpa4gj (nk0icy0xeofyyx1w_l ),
  .ysl1y4xf1(otcdnhpg8mwltf)
);

wire i_nnb5tc7xe6=(ktu7z7eeks17&wufvkpcwv_7l53) | (p5l63dwt7156pi&uqcuak_gzilz7mrpz0) | (oxt4ewm09j&y022y5lgu5q5z_i);
wire z1ot6fwfi2ihrl =(ktu7z7eeks17&ilnldo2qebgfdabgfq ) | (p5l63dwt7156pi&nk0icy0xeofyyx1w_l ) | (oxt4ewm09j&tqt6kzwmx2e3h2 );
wire aarvtm8rud8z0k4=(ktu7z7eeks17&zrotme_c1tv9ggx) | (p5l63dwt7156pi&otcdnhpg8mwltf) | (oxt4ewm09j&y2hpqatjf4b06o47va);
wire [68-1:0] mi_b4b0k5uuzd41;
wire [68-1:0] bghobt3obp5;


assign spfqyly64[68-1-1:0] = iily74b8[68-1:1] ;
assign spfqyly64[68-1] = 1'b1 ;

c2dm5oqn6257o319rma1kr9 jzbq22qrcr629tqzyd3b2zt(
  .rydw     (r5utfvc7oz),
  .d4y     (vqxjyefxtk),
  .iev4j_o4 (ptl5g3zjau),
  .hfl_1crp (ptvzkd3c5gfz85),
  .ysl1y4xf1(aarvtm8rud8z0k4),
  .w0m_yvp2sos8e(i_nnb5tc7xe6),
  .dtgamdbpa4gj (z1ot6fwfi2ihrl ),
  .xphx    (mi_b4b0k5uuzd41),
  .fap75    (bghobt3obp5)
);

assign dqm4y5o  = k2xz1iocfj4qk7btop ? olgpxn  : (aarvtm8rud8z0k4 ? vpvwojcah : idpqk) & spfqyly64 | ~{68{z1ot6fwfi2ihrl}} & ~spfqyly64 ;
assign tzwq6o86 = k2xz1iocfj4qk7btop ? vdmf0obdru6b : (i_nnb5tc7xe6 ? idpqk : vpvwojcah) & spfqyly64 | {68{z1ot6fwfi2ihrl}} & ~spfqyly64 ;

assign kktrbu07 = k2xz1iocfj4qk7btop ? ctoy95b : mi_b4b0k5uuzd41;
assign kf9hl8c_ = k2xz1iocfj4qk7btop ? zlq70vuuuc : bghobt3obp5;

endmodule



module c2dm5oqn6257o319rma1kr9(
  input [68-1:0] rydw,
  input [68-1:0] d4y,
  input [68-1:0] iev4j_o4,
  input [68-1:0] hfl_1crp,
  input ysl1y4xf1,
  input w0m_yvp2sos8e,
  input dtgamdbpa4gj,
  output [68-1:0] xphx,
  output [68-1:0] fap75
);
wire [68-1:0] scerhy06y;
wire [68-1:0] kybl1x84k6ea;
assign scerhy06y = {rydw[68-1-1:0], 1'b0} ;
assign kybl1x84k6ea [68-1:1] = d4y[68-1-1:0] ;
assign kybl1x84k6ea [0] = w0m_yvp2sos8e ;
wire [68-1:0] rjjjs3lcw9 = hfl_1crp & {68{w0m_yvp2sos8e & ~dtgamdbpa4gj}} 
                        | iev4j_o4 & {68{~w0m_yvp2sos8e & ~dtgamdbpa4gj}} ;

l3hw_f8igiui51siqdj 
#(.onr7l(68)) 
ag_zmq4ehicv__fmnmhhofu8sp1(
      .frgfco(scerhy06y), 
      .ii(kybl1x84k6ea), 
      .fij51v(rjjjs3lcw9), 
      .c(fap75),
      .s(xphx)
) ;
endmodule 



module qp2s59tux3j91cdjqs(
  input [68-1:0] rydw,
  input [68-1:0] d4y,
  output w0m_yvp2sos8e,
  output dtgamdbpa4gj ,
  output ysl1y4xf1
);

wire [3:0] wv9;
assign wv9 = rydw[68-1-1:68-1-4] + d4y[68-1-1:68-1-4] ;
assign w0m_yvp2sos8e = ~wv9[3] ;
assign dtgamdbpa4gj = &wv9[3:0];
assign ysl1y4xf1 = wv9[3] & ~(wv9[2] & wv9[1] & wv9[0]) ;

endmodule



                



module crj9jaav6wgkqbu1 #(
  parameter onr7l=64,
  parameter hw3qvr=6
)(
  input [onr7l-1:0] bjh,
  output [hw3qvr-1:0] ht70
);

wire [onr7l-1:0] cvf2uttd2wy;

assign cvf2uttd2wy[onr7l-1] = bjh[onr7l-1];

genvar j;
generate 
 for (j=onr7l-2; j>=0; j=j-1) begin: m_j0ywdyf2
    assign cvf2uttd2wy[j] = (|bjh[onr7l-1:j]);
 end
endgenerate

wire [onr7l-1:0] i = cvf2uttd2wy & {1'b1,~cvf2uttd2wy[onr7l-1:1]};

assign ht70[0]=( i[00] | i[02] | i[04] | i[06] | i[08] |
                i[10] | i[12] | i[14] | i[16] | i[18] |
                i[20] | i[22] | i[24] | i[26] | i[28] |
                i[30] | i[32] | i[34] | i[36] | i[38] |
                i[40] | i[42] | i[44] | i[46] | i[48] |
                i[50] | i[52] | i[54] | i[56] | i[58] |
                i[60] | i[62] );

assign ht70[1]=( i[00] | i[01] | i[04] | i[05] | 
                i[08] | i[09] | i[12] | i[13] | 
                i[16] | i[17] | i[20] | i[21] | 
                i[24] | i[25] | i[28] | i[29] | 
                i[32] | i[33] | i[36] | i[37] |
                i[40] | i[41] | i[44] | i[45] | 
                i[48] | i[49] | i[52] | i[53] | 
                i[56] | i[57] | i[60] | i[61] );

assign ht70[2]=( i[00] | i[01] | i[02] | i[03] | 
                i[08] | i[09] | i[10] | i[11] | 
                i[16] | i[17] | i[18] | i[19] | 
                i[24] | i[25] | i[26] | i[27] | 
                i[32] | i[33] | i[34] | i[35] |
                i[40] | i[41] | i[42] | i[43] | 
                i[48] | i[49] | i[50] | i[51] | 
                i[56] | i[57] | i[58] | i[59] );

assign ht70[3]=( i[00] | i[01] | i[02] | i[03] | i[04] | i[05] | i[06] | i[07] | 
                i[16] | i[17] | i[18] | i[19] | i[20] | i[21] | i[22] | i[23] | 
                i[32] | i[33] | i[34] | i[35] | i[36] | i[37] | i[38] | i[39] | 
                i[48] | i[49] | i[50] | i[51] | i[52] | i[53] | i[54] | i[55] );

assign ht70[4]=( i[00] | i[01] | i[02] | i[03] | i[04] | i[05] | i[06] | i[07] |
                i[08] | i[09] | i[10] | i[11] | i[12] | i[13] | i[14] | i[15] | 
                i[32] | i[33] | i[34] | i[35] | i[36] | i[37] | i[38] | i[39] |
                i[40] | i[41] | i[42] | i[43] | i[44] | i[45] | i[46] | i[47] );

assign ht70[5]=( i[00] | i[01] | i[02] | i[03] | i[04] | i[05] | i[06] | i[07] |
                i[08] | i[09] | i[10] | i[11] | i[12] | i[13] | i[14] | i[15] | 
                i[16] | i[17] | i[18] | i[19] | i[20] | i[21] | i[22] | i[23] |
                i[24] | i[25] | i[26] | i[27] | i[28] | i[29] | i[30] | i[31] );

endmodule

module t9iz7s9l43z8zrzmf #(
  parameter onr7l=32,
  parameter hw3qvr=5
)(
  input [onr7l-1:0] bjh,
  output [hw3qvr-1:0] ht70
);

wire [onr7l-1:0] cvf2uttd2wy;

assign cvf2uttd2wy[onr7l-1] = bjh[onr7l-1];

genvar j;
generate 
 for (j=onr7l-2; j>=0; j=j-1) begin: m_j0ywdyf2
    assign cvf2uttd2wy[j] = (|bjh[onr7l-1:j]);
 end
endgenerate

wire [onr7l-1:0] i = cvf2uttd2wy & {1'b1,~cvf2uttd2wy[onr7l-1:1]};

assign ht70[0]=( i[00] | i[02] | i[04] | i[06] | i[08] |
                i[10] | i[12] | i[14] | i[16] | i[18] |
                i[20] | i[22] | i[24] | i[26] | i[28] |
                i[30] );
                 

assign ht70[1]=( i[00] | i[01] | i[04] | i[05] | 
                i[08] | i[09] | i[12] | i[13] | 
                i[16] | i[17] | i[20] | i[21] | 
                i[24] | i[25] | i[28] | i[29] );
                

assign ht70[2]=( i[00] | i[01] | i[02] | i[03] | 
                i[08] | i[09] | i[10] | i[11] | 
                i[16] | i[17] | i[18] | i[19] | 
                i[24] | i[25] | i[26] | i[27] ); 
                

assign ht70[3]=( i[00] | i[01] | i[02] | i[03] | i[04] | i[05] | i[06] | i[07] | 
                i[16] | i[17] | i[18] | i[19] | i[20] | i[21] | i[22] | i[23] ); 
                

assign ht70[4]=( i[00] | i[01] | i[02] | i[03] | i[04] | i[05] | i[06] | i[07] |
                i[08] | i[09] | i[10] | i[11] | i[12] | i[13] | i[14] | i[15] ); 


endmodule



























module a3zxpqwwtl53hi(

  
  
  
  
  input                                   z4za08k83of9q, 
  output                                  d9f119ap_n00k, 
  input  [64-1:0]                 dq0a9sotg74w,
  input  [64-1:0]                 netnmrvccmf,
  input  [64-1:0]                 qaxmne8xc_,
  input  [19-1:0] v48iyoy1fdeh,
  input  [4-1:0]           gcl2zxzh4brhr,

  output                                  ogtxqxlymgsff9qr,

  
  
  
  output                  jfgbmn4y_79lt81, 
  input                   tsa8otson44it2, 
  output [64-1:0] du9nxa6qo7knx2et1gw6,
  output                  h7szh92q4s7x6vx_,   

  
  
  
  output                        isz7jw04u7k3s7b398, 
  input                         q4_7fnx90rztwn6_8dybi, 
  output [64-1:0]       zq2e9j_emlri_qjtg,
  output                        qv749hsiom75nyn49v,   
  output [4-1:0] gw6s_h2ymbn1ds50q8,
  
  input  gf33atgy,
  input  ru_wi
  );

  wire pn5sglj4k8u17arywgn;

    
  assign h7szh92q4s7x6vx_  = 1'b1;
  assign du9nxa6qo7knx2et1gw6 = 64'b0;

  assign d9f119ap_n00k = 
           (tsa8otson44it2)  
         & (pn5sglj4k8u17arywgn); 

  wire   gr5ok7alh29knnfzuu0 = z4za08k83of9q & tsa8otson44it2;
  assign jfgbmn4y_79lt81 = z4za08k83of9q & pn5sglj4k8u17arywgn;

 localparam jwxxo5dwz741q1 = 64*2 + 19 + 4;

 wire [jwxxo5dwz741q1-1:0] nks3h78aq1ssl9a;
 wire [jwxxo5dwz741q1-1:0] oa9guo_6_;

 wire [64-1:0] artnbioj;
 wire [64-1:0] emfjxicm;
 wire [4-1:0] qbpmsk2;
 wire [19-1:0] ql3pltf;
 wire [19-1:0] s5e1ijt4hac;

 assign nks3h78aq1ssl9a ={
                       dq0a9sotg74w
                     , netnmrvccmf
                     , v48iyoy1fdeh
                     , gcl2zxzh4brhr
                     };
 
 assign             {
                       artnbioj
                     , emfjxicm
                     , ql3pltf
                     , qbpmsk2
                     } = oa9guo_6_;

 wire jjzotrbn; 
 wire hw1_k1jmu; 

 ux607_gnrl_pipe_stage # (
  .CUT_READY(1),
  .DP(1),
  .DW(jwxxo5dwz741q1)
 ) k75wa_p8zgd6rkhhbze (
   .i_vld(gr5ok7alh29knnfzuu0), 
   .i_rdy(pn5sglj4k8u17arywgn), 
   .i_dat(nks3h78aq1ssl9a  ),
   .o_vld(jjzotrbn), 
   .o_rdy(hw1_k1jmu), 
   .o_dat(oa9guo_6_ ),
 
   .clk  (gf33atgy  ),
   .rst_n(ru_wi)  
  );


  wire [67-1:0] wanhh3qu4ohss9m;
  wire [67-1:0] vwbsb33jbcgdblb;
  wire                                c6mg4aw3ydy52bnar ;
  wire                                rzgepy3r4ibso2v3ea7r ;
  wire [67-1:0] cpl0d1l0rfztufu;

  wire          tcioj21iaq52vw3;
  wire [64:0] d8cf11_gw8vhq;
  wire [64:0] r87cg11xdmmo6m1i;

  wire          ehlal_jbp2qi9wkr8;
  wire [64:0] ych1yr4tro3wfb7hy;
  wire [64:0] x20j55p_9ns4u;


  assign s5e1ijt4hac[3:0          ] = ql3pltf[3:0 ];
  assign s5e1ijt4hac[4:4         ] = ql3pltf[4:4];
  assign s5e1ijt4hac[5:5   ] = 1'b0;
  assign s5e1ijt4hac[6:6  ] = 1'b0;
  assign s5e1ijt4hac[7:7] = 1'b0;
  assign s5e1ijt4hac[8:8 ] = 1'b0;
  assign s5e1ijt4hac[9:9   ] = ql3pltf[9:9   ];
  assign s5e1ijt4hac[10:10  ] = ql3pltf[10:10  ];
  assign s5e1ijt4hac[11:11   ] = ql3pltf[11:11   ];
  assign s5e1ijt4hac[12:12  ] = ql3pltf[12:12  ];
  assign s5e1ijt4hac[13:13   ] = ql3pltf[13:13   ];
  assign s5e1ijt4hac[14:14  ] = ql3pltf[14:14  ];
  assign s5e1ijt4hac[15:15  ] = ql3pltf[15:15  ];
  assign s5e1ijt4hac[16:16 ] = ql3pltf[16:16 ];
  assign s5e1ijt4hac[17:17  ] = ql3pltf[17:17  ];
  assign s5e1ijt4hac[18:18 ] = ql3pltf[18:18 ];


  wire                        sti6zw89hiczcu_iz ; 
  wire                        qnzni53zqm9butd ; 
  wire [64-1:0]       nfwuyk8cl0ce6umv4v  ;
  wire                        b6648sfmn8rxay   ;   
  wire [4-1:0] c5t7d65j1bt68x7 = qbpmsk2 ;
  

  uflzl0cx7tik0xzqybt c4q88mqbrzua266_ol7k9hq(

      .kg5ogiwmi4x2jcasma      (jjzotrbn),
      .rbjqmkcrkr7uyq4dauq      (hw1_k1jmu),
                           
      .w56hh_dniqksvhf        (artnbioj      ),
      .q6e0lb86_tx2afeh        (emfjxicm      ),
      .i5vvhea8kczaa        (64'b0      ),
      .umfak1vbx2r1b       (s5e1ijt4hac),
      .l3kh5v32kt2mkcqz6t   (),
      .i1gdm9hju_gidl       (4'b0),
                          

          
      .dnmtm28bd2t         (1'b0    ),

      .qqrzyv7p9gfzn99      (sti6zw89hiczcu_iz    ),
      .ori3109ceulwf9p      (qnzni53zqm9butd    ),
      .p3nl1p59c7tkqhr5l8rl  (nfwuyk8cl0ce6umv4v),
      .sw6cd2q81orxwjah_hdqq9   (b6648sfmn8rxay ),

      .alse1t6spxo4msbspebwy3y  (wanhh3qu4ohss9m),
      .x0er7wym12k2zbbkwic3tk  (vwbsb33jbcgdblb),
      .g35fohnhd6cn9np610_  (c6mg4aw3ydy52bnar),
      .nn3y8_8tdpg0r00cfh22  (rzgepy3r4ibso2v3ea7r),
      .tvohxqv2vynsps11_n8jcm1  (cpl0d1l0rfztufu),
      
      .b9_gjh0acfnkvdnxisky4    (tcioj21iaq52vw3  ),
      .kjts4h4q5dfneeyrrdrxw    (d8cf11_gw8vhq  ),
      .sco_wqinvslwrh      (r87cg11xdmmo6m1i    ),
     
      .sj_mdw9rcnoy3tw08nw    (ehlal_jbp2qi9wkr8  ),
      .bx56_yppcspoez2oo86i    (ych1yr4tro3wfb7hy  ),
      .tjsikyyrigiuo_      (x20j55p_9ns4u    ),

      .gf33atgy                 (gf33atgy               ),
      .ru_wi               (ru_wi             ) 
  );

 localparam lgs5lf2mxxr_do2xuk_ = 64+4;
 wire [lgs5lf2mxxr_do2xuk_-1:0] zx4e1q4vx0hpooq = {nfwuyk8cl0ce6umv4v, c5t7d65j1bt68x7};
 wire [lgs5lf2mxxr_do2xuk_-1:0] houn75bo0_82oq7b;
 ux607_gnrl_pipe_stage # (
  .CUT_READY(0),
  .DP(1),
  .DW(lgs5lf2mxxr_do2xuk_)
 ) g3rauzz0reiwsdvzwra35i (
   .i_vld(sti6zw89hiczcu_iz), 
   .i_rdy(qnzni53zqm9butd), 
   .i_dat(zx4e1q4vx0hpooq ),
   .o_vld(isz7jw04u7k3s7b398), 
   .o_rdy(q4_7fnx90rztwn6_8dybi), 
   .o_dat(houn75bo0_82oq7b ),
 
   .clk  (gf33atgy  ),
   .rst_n(ru_wi)  
  );
  assign {zq2e9j_emlri_qjtg,gw6s_h2ymbn1ds50q8} = houn75bo0_82oq7b;
  assign qv749hsiom75nyn49v = 1'b0;
  
  
  
  ux607_gnrl_dffl #(64+1) l_umgyq0nvgdi2z2 (tcioj21iaq52vw3, d8cf11_gw8vhq, r87cg11xdmmo6m1i, gf33atgy, ru_wi);
  ux607_gnrl_dffl #(64+1) ld1t7i795rr21jgz (ehlal_jbp2qi9wkr8, ych1yr4tro3wfb7hy, x20j55p_9ns4u, gf33atgy, ru_wi);

    
  
  

  wire [67-1:0] ti2vpd9jde = wanhh3qu4ohss9m;
  wire [67-1:0] xfvd9b_1bqsugi = vwbsb33jbcgdblb;

  wire knqibikmye3;
  wire [67-1:0] atsytx8oasf;
  wire [67-1:0] d_h0rtp1mu2fy;
  wire [67-1:0] wrcjvt7pl1j_;

  wire qqjhj5cz1ue = c6mg4aw3ydy52bnar ;
  wire gn6aq7h3cy = rzgepy3r4ibso2v3ea7r ;

  wire nuhvvo7aaoun4df0 = qqjhj5cz1ue | gn6aq7h3cy; 
  

     
  assign atsytx8oasf = {67{nuhvvo7aaoun4df0}} & (ti2vpd9jde);
  assign d_h0rtp1mu2fy = {67{nuhvvo7aaoun4df0}} & (gn6aq7h3cy ? (~xfvd9b_1bqsugi) : xfvd9b_1bqsugi);
  assign knqibikmye3 = nuhvvo7aaoun4df0 & gn6aq7h3cy;

  assign wrcjvt7pl1j_ = atsytx8oasf + d_h0rtp1mu2fy + {{67-1{1'b0}},knqibikmye3};

  assign cpl0d1l0rfztufu = wrcjvt7pl1j_;

  
  assign ogtxqxlymgsff9qr  = 1'b0;

endmodule                                      






















module qaszx6xv9r9g8927s (
  output  tywculgjyor8ndw,
  output  btwmhh91h50d5flgwx4o6pwu,

  input   a02zzbowpjn06h,
  input   se2buoxmq91dbic3y2m5hu,
  output   e9u0rtvt8jrygyc8s,

  output av1w8ld09cfofn,
  output im2b5l0h98avl6t4sj,
  output bw65wl7fvekfymd8vqx,
  output [64-1:0] pecbpcoa04vq,
  output [64-1:0] tb_snaxyfs,
  output [64-1:0] zc4mldgm25r,
  output [32-1:0] d23wb5yh1iyvf,
  output [1:0] srim3bfnzhve,
  output cy3nuhzm_v2p73mt,
  output fvqwdz2hdbb,

  input feq1g7m2cy1erl,


  input rvr30vvllni,

  input   w2fpnf5fg1byp6,

  output [11:0] k3cmpuswk7in0u4,


  input  [64-1:0] k84xk2u4clez     ,
  input                      jd2_q1xken6mnd8v ,
  input                      tb198r6lzk1sr77g4 ,
  input  [64-1:0] cvvsn7xc8qg5uk     ,
  input                      jp82o1hu0f41an   ,



  output  tw5xnp59d8x,
  output  y_0q8d40rrzolo1y6,
  output  qwcb6hcmvfqmf032z,
  input   ao17frh5wnr0wddz3,
  input   woon4h3ivznl_qiu7i_9,
  input   [4-1:0] p25dd0cxz7nmi6w9ebukmr,
  output  [4-1:0] uvgy9al0j8prciqsh,
  output  f8pn1x6gurodpy04d3j1ihn,
  output  mmludd_fnt2yevok8a1a0,
  input   buwj9_8l8bwj80kkinq9p,

  input   apid0ys34zyekptw7un,
  output  um8zsjyxn_4p,  

  input   h7fseh5_df0hbx,

  output  c8w01x5rfmr6shqzb,
  input   p7rj2v1hvh0nab6ei       ,
  input   fe8u85vitwnfnuszhl          ,
  input   stx6pefjqd_oqqg5gej9       ,
  input   u3qmzjrm6inkod3m3ghp     ,
  input   wkyo2nrlaz9sq3m1chcysnofuenz ,
  input   vmkmkz3cm8cgbet959d4pw_0ti,
  input   gnn94t_31a_j59f483ym5f68sb    ,     
  input   zb322_7v29pmo4jvmvow3qi8  ,

  input   qsn_nfmbj97wz1r3s59t2 ,
  input   uuvo0ter1b1y6j1xfc ,
  input   hjysp7ahvean99t41k89pt ,
  input   ggvuzlnuknlvg4a50n4hy7ok ,
  input [5-1:0] frfbo512g1_94ncrem_be859f, 
  input [64-1:0] lt3biawnyshgr5rw4q5chcg6u7rc,
  input   j6g8r7rblr88am07jc3i5 ,
  input   klz7l8_75czqn63zb ,
  input   esb6gep_3iit0w ,
  input   iq2e_b4p5qjp2ryy5sktbl6kd0 ,
  input   om206h86cfrb69iqc9pzq3fq1 ,
  input   yk85cwkls6hcvp4_g70j2 ,
  input   cj2z8_7e4hw2s1u6mhckmpm4i ,
  input   rpt826mhm0kwty9qlty6rt1 ,
  input   pmcsf3olv_ztinoakqw67nno42plkv ,
  input   dgigaix0xkzcg64kbmiqjlagh1cqid2 ,
  input   m2av7b78yjzgy1j3a9inerkjyzrkdg9 ,
  input   z2tyajok7rez0sc5ugh28p8o0rsrq ,
  input   o2rr0tomxjme9ua4btx71i4hsfz ,
  input   [64-1:0] n7orghfl8x_7wsaisuhpw9o,
  input   [64-1:0] wql66zm9cb_1pzbk,
  input   [32-1:0] skcwu9hiw7zl59wu,
  input   ij7ql6t124xbofcx,
  input   z2574r4ajgr7u7mtpb_wpetx,
  input   fof2qu1zf51j1nid7vs4,
  input   umg0x8yb1yqjkaw34l6t,

  input   [64-1:0] lovkp0eqfnxtb7,


  input   fi9wz0kme0ey_bxavdqx_9,
  input   tmhbzyv2b510vt_9qkb16hdwa,
  input   nqoqg40hg82wgdbsfubvu4fg,
  input   hcx0jkab_j87_6j7phxnsz,
  input   t0zuyah73tpfg_dtxy56ug9ej,
  input [64-1:0] sq0y2gv0vwpq_6ckk9b89gybz,
  output  i32x_jtt7bvmr9lu2p,
  input   mxa77etukhs8o_5z6962l19,
  input   cd4v4c_rw906kt5,
  input   idat72abxke4z9s,
  input   hv4wuttuo9jk_cqa8sxqwt , 
  input   ac8_dky9fhpbsxu0b9t88ag8 , 

  input   [64-1:0] r_8f7p3tznijza5y03ko,



  output  ip4b_cj6h98z45oey8l,

























  output  oyiml9jn3w6vt88yja9asjx,
  output  glime27x19feqrvvsa2nmeh5f,


  output  ljd_sv9l5ykkrwitvxjydqd5n55,  
  output  wrg2t13vafz_5z44ejdmrpmnk1,  
  output  g7cxea_49xi94dndcklkkq,  
  output  vj6p6j6avq664060js8d_wit_7a,  


  output  [64-1:0] vfga_wjq02bdlelajwej,  


  input   o7hoht1pqz01v7,
  input   [64-1:0] kbv2bs_lxmvu,

  input   [64-1:0] unbt3q05xijb,
  input   [64-1:0] hawbmpz6j7pzibqr,

  input   jw4fsjecr0u919fr7,
  input   fh49u69v0he,
  input   af5qc04tmn51e4u2h1z,

  output  [64-1:0] wtd_nuaeb_mpye,
  output  [64-1:0] elth4vimq_j,


  output  [64-1:0] xd66pm611ai1dg,
  output  x7eg618xaszd4f21cl_g,
  output  r9uxubpl2h2alj1q,
  output  jlud6jeuxe0espga,

  input   [64-1:0] pldoasxyzlvx2,
  input   [64-1:0] bde41te346q515l,

  output  sf0uuehfhfa,
  output  hvy2cpsp75f3,
  output  k3z202os,
  output  z35xlcc6bt4,
  output  [64-1:0] ew08uu2kn2p9e11s,
  output  xv08lot3vi9dag4vs0,
  output  [64-1:0] mtc04rctrfyb,
  output  if5jz8qk0aqefy3v35o,



  input   fcjh1nct4r,
  input   [9:0] b4lwcgm6l21pi,
  input   zwcbp7zqfei5xz,
  input   dn8riluj40uunvq5,
  output  dz0zrf512290tvcy4q,
  input   [64-1:0]  z0yhjfv_e0yaa2r,

  output  z1l80uwh6vyyg34,
  input   rn1o3sl83,

  input   uc5qxb4d2b28ye5,
  output  o2qkf90r783,




  input   s5f_36xvqrtq7,


  input   x6eltyshbu5,
  input   lt3v_fm0ipu,
  input   v3ne7glf8d8,
  input   v9dnbgjy6c0vf,
  input   hmzw4exmjn8k921c,

  input   siifnhwgancn8,
  input   mfzl2fqml69hx,
  input   aw0hbwfkx3f63s,
  input   u83p4flbuvkqt26z,
  input   tvglhc8o_izdq,

  input   pydatzxqqi,

  input   c4ughu0qm5sfai,

  input   w632tcbtqncn6,
  input   ai169tbqp4seb3,
  input   b0zz_ornhz010,
  input   yw4o4kdms07_32,
  input   ezl3jzeqhltgj7h,
  input   w529wbj853,
  input   i9xvsmm45fp0f58,
  input   [64-1:0]     r4bs4k_53n5wp,


  input   jqsukc5b5drcc1e78,
  input   gnn46rd7vvofruqij,
  input   vkyge0q4mfc5,
  input   [64-1:0]     cppkd01vpwwnlfy,
  input   [64-1:0]  d3hccrck1fl7jjf6,
  input   [64-1:0]     h_qwsgi7nk2,

  output  [64-1:0]     u25pqekq4df,
  output                       dhjwho76fa8hqc,
  output  [64-1:0]     xel6gw173w5x0,
  output                       icauf4l_12_c2xkj53lf,
  output  [64-1:0]     v8ydjtlz16x9tx,
  output                       e_z6d7r9kxqg32te,
  output  [64-1:0]  p5jpgn4rvarpo,
  output                       z2g63deibg1b1quqr,
  output  [64-1:0]     tlgcdv86voe9,
  output                       u_ufp_wg29ieoklxxz1,

  output  [64-1:0] qeb3z0x5,
  output  ibhfuwrztbm8p4gg,
  output  [3-1:0] i8_5wt0vppx,
  output  osv2437qj_3nuf,


  output  b7g_vsn0zoewh6g1,
  output  [2-1:0] onnv64ydiajl,


  input   c5ewdqztjw9za,
  input   rn2mt6nngsc9w5cz,
  input   t5trf35s8vy,
  input   zbac123pv78sbz3,
  input   z4e_m564fxae0kpbjr,
  input   hixy2y36a1pn0,
  input   ozwene1gdpatk6g,

  input  [64*4-1:0] azll7rq5fab5ou,
  input  [64*4-1:0] n6a0r_0zddzrme8,
  output ns0i7siujgkrghjpqv6,

  input   um28jgd2x4mbs,

  input   aw82i964do,
  input   y8_gkxsfle,
  input   cwwkpmk260lrt,

  output  qo5p9t6s74zxpo,

  input   dk2xhkj77a,
  input   gf33atgy,
  input   ru_wi
  );
  localparam urjif1vu4pqgqxt4x8 = 51;
  localparam m_rz39tx6bnugdx = (urjif1vu4pqgqxt4x8<=2)?1:(urjif1vu4pqgqxt4x8<=4)?2:(urjif1vu4pqgqxt4x8<=8)?3:(urjif1vu4pqgqxt4x8<=16)?4:(urjif1vu4pqgqxt4x8<=32)?5:(urjif1vu4pqgqxt4x8<=64)?6:(urjif1vu4pqgqxt4x8<=128)?7:(urjif1vu4pqgqxt4x8<=256)?8:(urjif1vu4pqgqxt4x8<=512)?9:(urjif1vu4pqgqxt4x8<=1024)?10:(urjif1vu4pqgqxt4x8<=2048)?11:(urjif1vu4pqgqxt4x8<=4096)?12:-1;
  localparam v_1vibiyou7ysbpkunv = (urjif1vu4pqgqxt4x8  < 32) ? 7 : (m_rz39tx6bnugdx + 2);



  wire y5pha1zmcujhhs6sq = 1'b0;
  wire ar2xblav711he9vqcjg8nxq = 1'b0;
  wire e1645180ujgpiuebeqa = 1'b0;
  wire evla4t4m7kx62w598l = 1'b0;
  wire oxberxo5xs4cqy454m0 = 1'b0;

  wire bkjtjv8qktytwklm1;
  wire mp89sr5uys176dofb6r;

  assign tywculgjyor8ndw = bkjtjv8qktytwklm1 | mp89sr5uys176dofb6r;






  wire bet3r1ns0njrwezuu;
  wire cn7vi2ekbeqvap2074co5n33s;






  wire xjzmsfojv82w58 = (y_0q8d40rrzolo1y6 & tw5xnp59d8x & qwcb6hcmvfqmf032z & woon4h3ivznl_qiu7i_9)
                            & (mmludd_fnt2yevok8a1a0 & buwj9_8l8bwj80kkinq9p)
                            & (~a02zzbowpjn06h) 
                          ;


  wire q7r68kfb621_p;
  wire r18u32nuzxrk;
  wire z5sexv2;



  wire o7ou0irmq_m20mo9iaidwbxx3f;



  wire sjiqvq4geh18r8dpd = 1'b0
      | tw5xnp59d8x 
      ;
  wire x76a6w0qgnegw5;

  wire m0hir9b4vzdlau = xjzmsfojv82w58 & (~sjiqvq4geh18r8dpd) & (~x76a6w0qgnegw5);
  wire ajfpr1hse233eo9zr = m0hir9b4vzdlau | sjiqvq4geh18r8dpd;

  wire vnijg2dqxrwcg = m0hir9b4vzdlau & (~sjiqvq4geh18r8dpd);


  ux607_gnrl_dfflr #(1) d_wpq5kp_cyqpize (ajfpr1hse233eo9zr, vnijg2dqxrwcg, r18u32nuzxrk, dk2xhkj77a, ru_wi);
  assign tw5xnp59d8x = r18u32nuzxrk;

  wire sl491lvt7orov19r0 = ajfpr1hse233eo9zr ? vnijg2dqxrwcg : r18u32nuzxrk;
  wire vhwvqw2isian0 = sl491lvt7orov19r0;

  wire mv5lq3jts3ftcrxz2h = (sl491lvt7orov19r0 & apid0ys34zyekptw7un);
  ux607_gnrl_dffr #(1) vlpctplxjxzbkce (mv5lq3jts3ftcrxz2h, um8zsjyxn_4p, dk2xhkj77a, ru_wi);


  wire mf_9_fzjbuyej45vf = sjiqvq4geh18r8dpd & r18u32nuzxrk;
  wire sbkebsnoxe_flm = x76a6w0qgnegw5;
  wire b3r1_vbhjziooe2conb = mf_9_fzjbuyej45vf | sbkebsnoxe_flm;
  wire i7uaj2m98c9j2d = mf_9_fzjbuyej45vf & (~sbkebsnoxe_flm);
  ux607_gnrl_dfflr #(1) d9lwa0k0ug1dqwzgfi (b3r1_vbhjziooe2conb, i7uaj2m98c9j2d, x76a6w0qgnegw5, dk2xhkj77a, ru_wi);










  wire stoyzmp_n_xpa90k = esb6gep_3iit0w & fh49u69v0he;
  wire wolnms170782my7_gk = stoyzmp_n_xpa90k & (~pydatzxqqi);
  wire u5a92wwchl7sg75h;
  wire [4-1:0] wh00ey3j8j7cuxdpqnag;




  wire a_fwigc8tf1pwpa_h4rd = ip4b_cj6h98z45oey8l; 
  wire rwe32f8r_3ajh9xkq = x76a6w0qgnegw5 | (u5a92wwchl7sg75h & a_fwigc8tf1pwpa_h4rd);

  wire fedy8pl1rxkooxtsv_0 = wolnms170782my7_gk | rwe32f8r_3ajh9xkq;

  wire ok_yh0erb9nokqy54 = wolnms170782my7_gk & (~rwe32f8r_3ajh9xkq);
  ux607_gnrl_dfflr #(1) osvptmp0c77j7j401vj2q (fedy8pl1rxkooxtsv_0, ok_yh0erb9nokqy54, u5a92wwchl7sg75h, gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(4) w5aawf29_9_jt6v69y2a9un (fedy8pl1rxkooxtsv_0, p25dd0cxz7nmi6w9ebukmr, wh00ey3j8j7cuxdpqnag, gf33atgy, ru_wi);



  assign y_0q8d40rrzolo1y6 = u5a92wwchl7sg75h
                          & tb198r6lzk1sr77g4 



                            ;



  assign qwcb6hcmvfqmf032z = u5a92wwchl7sg75h  
                          & tb198r6lzk1sr77g4   



                            ;
  assign f8pn1x6gurodpy04d3j1ihn = u5a92wwchl7sg75h; 
  assign uvgy9al0j8prciqsh = wh00ey3j8j7cuxdpqnag;

  assign mmludd_fnt2yevok8a1a0 = u5a92wwchl7sg75h
                          & tb198r6lzk1sr77g4 



                            ;

  wire kynmn08sx90nf4lm2aki6okl = 
                                (qwcb6hcmvfqmf032z ? 1'b1 : jd2_q1xken6mnd8v)   
                              & (!se2buoxmq91dbic3y2m5hu)

                              & (qwcb6hcmvfqmf032z ? tb198r6lzk1sr77g4 : ~tb198r6lzk1sr77g4)
                              & (~jp82o1hu0f41an)  
                              ;





  wire rjjrzh_tco6hcost86;























  wire zxz41rcq69i2tnl6wx1lz2t = kynmn08sx90nf4lm2aki6okl; 

  wire wmeyhl03a273zu2s7qupf5h = rjjrzh_tco6hcost86
                              & zxz41rcq69i2tnl6wx1lz2t;



  assign i32x_jtt7bvmr9lu2p = zxz41rcq69i2tnl6wx1lz2t;
























  wire u9s6l7o34d25v4npe6zl = (~rjjrzh_tco6hcost86) 
                              & kynmn08sx90nf4lm2aki6okl  
                              ;

  wire xo1uoocz53uginn8n        = y5pha1zmcujhhs6sq 
                              & u9s6l7o34d25v4npe6zl;




  wire ya4_xt1c2gbjveqcssfkrflo3yj4kza = (~rjjrzh_tco6hcost86) & (~y5pha1zmcujhhs6sq) 
                              & kynmn08sx90nf4lm2aki6okl  

                              & (~feq1g7m2cy1erl) 
                              ;

  wire usl0bxdbhf2_xj;
  wire lpofewte8nxu7_o;
  wire tg6dvyjbvr4lk8_esf1fjt = (usl0bxdbhf2_xj  | lpofewte8nxu7_o)
                              & ya4_xt1c2gbjveqcssfkrflo3yj4kza;
  wire v406rha54c4fv52jvro_wx_ = (usl0bxdbhf2_xj                  )  
                              & ya4_xt1c2gbjveqcssfkrflo3yj4kza;
  wire tg0gz600v1f7omqs_85rx6cnq3 = (                  lpofewte8nxu7_o)  
                              & ya4_xt1c2gbjveqcssfkrflo3yj4kza;




  wire ytk71a3aqo1gspmy46_28lj = (~rjjrzh_tco6hcost86) & (~y5pha1zmcujhhs6sq) & (~usl0bxdbhf2_xj) 
                              & kynmn08sx90nf4lm2aki6okl  

                              & (~feq1g7m2cy1erl) 
                              ;

  wire jukbv9h11v1o8cebnq        = z5sexv2
                              & ytk71a3aqo1gspmy46_28lj;



  wire q8aazbn3lcj5_rsvwyrh36o_glp_ermqiwjm = 
                              & (~z5sexv2) & (~rjjrzh_tco6hcost86) & (~y5pha1zmcujhhs6sq) & (~usl0bxdbhf2_xj) 
                              & kynmn08sx90nf4lm2aki6okl  

                              & (~feq1g7m2cy1erl) 
                              ;

  wire g1hkbyqaj8r_janme7jrc8rxe_rrb  = cn7vi2ekbeqvap2074co5n33s
                              & q8aazbn3lcj5_rsvwyrh36o_glp_ermqiwjm;







  wire w_406g1gnqqywd5j20dbpxvcebcs6jcb = 1'b1





                              ;

  wire kdpaa43ha_zuq8zsbp5o7u8a  = bkjtjv8qktytwklm1  
                              & w_406g1gnqqywd5j20dbpxvcebcs6jcb;





  wire i28kzhzarq9ngflg   = p7rj2v1hvh0nab6ei & mp89sr5uys176dofb6r;

  wire asclifx_kw21p4ynudz9aaaukgl6a4 = 



                                (~bkjtjv8qktytwklm1) ;



  wire m0ugsckv2bvgxdilc4lz   = i28kzhzarq9ngflg
                              & asclifx_kw21p4ynudz9aaaukgl6a4;












  assign c8w01x5rfmr6shqzb = w_406g1gnqqywd5j20dbpxvcebcs6jcb;

  wire pbtbpfm39qh0vekjwkog  = g1hkbyqaj8r_janme7jrc8rxe_rrb | kdpaa43ha_zuq8zsbp5o7u8a;


  wire   jbod2vk5w_ts8f0pmlikw9b7;


  assign o7ou0irmq_m20mo9iaidwbxx3f  = (tg6dvyjbvr4lk8_esf1fjt | xo1uoocz53uginn8n | wmeyhl03a273zu2s7qupf5h | pbtbpfm39qh0vekjwkog | jukbv9h11v1o8cebnq | m0ugsckv2bvgxdilc4lz);
  wire all_excp_flush_type;
  assign all_excp_flush_type = tg6dvyjbvr4lk8_esf1fjt | xo1uoocz53uginn8n | wmeyhl03a273zu2s7qupf5h | m0ugsckv2bvgxdilc4lz;

  assign ip4b_cj6h98z45oey8l  = (o7ou0irmq_m20mo9iaidwbxx3f) & (~tw5xnp59d8x) 

                            | x76a6w0qgnegw5
                              ;
  wire   kv0a6wk1ng1nyfl1xjkh34 = jbod2vk5w_ts8f0pmlikw9b7 & m0ugsckv2bvgxdilc4lz
                                 & (~tg6dvyjbvr4lk8_esf1fjt)
                                 & (~xo1uoocz53uginn8n)
                                 & (~wmeyhl03a273zu2s7qupf5h)
                                 ;

  assign glime27x19feqrvvsa2nmeh5f = 
             rjjrzh_tco6hcost86 | 
             usl0bxdbhf2_xj | 
             y5pha1zmcujhhs6sq | 
             cn7vi2ekbeqvap2074co5n33s |
             z5sexv2          ;

  assign oyiml9jn3w6vt88yja9asjx = 
             bkjtjv8qktytwklm1 |
             m0ugsckv2bvgxdilc4lz;

  wire wlotcqomlz6de0sr4ukuhgbwpu3n;
  wire r2ovgzxgcrqk7dmnynz6j1zh_61qmz = 
             rjjrzh_tco6hcost86 | 
             usl0bxdbhf2_xj | lpofewte8nxu7_o |
             y5pha1zmcujhhs6sq | 
             wlotcqomlz6de0sr4ukuhgbwpu3n |
             z5sexv2          ;



  assign qo5p9t6s74zxpo = r2ovgzxgcrqk7dmnynz6j1zh_61qmz; 


  wire cxij98yy3k4hy34_9o = ip4b_cj6h98z45oey8l;



  wire d7lhla0f70idm9pt;
  wire l89rffl8xklfzh4_e;
  wire n703xx6o97u6y;
  wire r5sqfkv0bsgn5k6la      = all_excp_flush_type & cxij98yy3k4hy34_9o;

  wire d7gc7q1qy89t05;
  wire xv76y4hz81uw_gu;
  wire gxmbdujixw2_0t7d527dq  =   (jukbv9h11v1o8cebnq & d7gc7q1qy89t05 & (~d7lhla0f70idm9pt) & (~n703xx6o97u6y) & cxij98yy3k4hy34_9o)
                             | (jukbv9h11v1o8cebnq & xv76y4hz81uw_gu & (~l89rffl8xklfzh4_e) & (~n703xx6o97u6y) & cxij98yy3k4hy34_9o);
  wire z1ri4yxi78_p8hx8y       = jukbv9h11v1o8cebnq & ( n703xx6o97u6y) & cxij98yy3k4hy34_9o;
  assign dz0zrf512290tvcy4q    = gxmbdujixw2_0t7d527dq;
  wire dbg_entry_taken_ena;
  assign dbg_entry_taken_ena = pbtbpfm39qh0vekjwkog & cxij98yy3k4hy34_9o;


  wire [64-1:0] n5_4v2cdhby2lv =  {unbt3q05xijb[64-1:2],2'b0};
  wire [64-1:0] faqz95ne3ps3e1o7d9 =  {hawbmpz6j7pzibqr[64-1:2],2'b0};
  wire [64-1:0] wsufrwtxevzipw =  {h_qwsgi7nk2[64-1:2],2'b0};
  wire [64-1:0] sco4chgj6vsbyoxn2j =  {kbv2bs_lxmvu[64-1:2],2'b0};
  wire [64-1:0] tx81df88wvd5cnr5h5 =  {cppkd01vpwwnlfy[64-1:2],2'b0};


  assign z1l80uwh6vyyg34 = z1ri4yxi78_p8hx8y;

  wire s74_qw0a41imkgkdcsf0rdhta;
  wire tf2ird6le5az6cmue2y6_;
  wire av15ikbsl_f;
  wire dbk9rh15g1;
  wire gvvhhfwk9lgdcu = 1'b1;

  wire [64-1:0] uolend5_94trunxfp6p5;

  assign {
      vfga_wjq02bdlelajwej,
      ljd_sv9l5ykkrwitvxjydqd5n55,
      wrg2t13vafz_5z44ejdmrpmnk1,
      g7cxea_49xi94dndcklkkq,
      vj6p6j6avq664060js8d_wit_7a
  } = 
      pbtbpfm39qh0vekjwkog ? {
          (32'h00000000 
            ),
              aw82i964do, 
              y8_gkxsfle, 
              1'b1,    
              1'b0  
          }:
      (all_excp_flush_type & kv0a6wk1ng1nyfl1xjkh34 & pydatzxqqi) ? {
          32'h00000000, 
              aw82i964do, 
              y8_gkxsfle, 
              pydatzxqqi, 
              1'b0  
         }:
      (all_excp_flush_type & pydatzxqqi) ? { 
          (32'h00000000 + 64'd4
            ),
              aw82i964do, 
              y8_gkxsfle, 
              pydatzxqqi, 
              1'b0  
         }:
      (jukbv9h11v1o8cebnq & n703xx6o97u6y) ? {
          faqz95ne3ps3e1o7d9,
              1'b1, 
              1'b0, 
              pydatzxqqi, 
              1'b0  
          } :
      (all_excp_flush_type & (~pydatzxqqi)) ? 
          ( 
           av15ikbsl_f ? {
             n5_4v2cdhby2lv,
                1'b1, 
                1'b0, 
                pydatzxqqi, 
                1'b0  
                } : {  
             wsufrwtxevzipw,
                1'b0, 
                1'b1, 
                pydatzxqqi, 
                1'b0  
                }  
          ) : 
        
      (jukbv9h11v1o8cebnq & d7gc7q1qy89t05 & (~dn8riluj40uunvq5) & (~n703xx6o97u6y) & (~d7lhla0f70idm9pt) ) ? {
            n5_4v2cdhby2lv ,
              1'b1, 
              1'b0, 
              pydatzxqqi, 
              1'b0  
          }:
      (jukbv9h11v1o8cebnq & xv76y4hz81uw_gu & (~dn8riluj40uunvq5) & (~n703xx6o97u6y) & (~l89rffl8xklfzh4_e) ) ? {
            wsufrwtxevzipw ,
              1'b0, 
              1'b1, 
              pydatzxqqi, 
              1'b0  
          }:
      (jukbv9h11v1o8cebnq & d7gc7q1qy89t05 & ( dn8riluj40uunvq5) & (~n703xx6o97u6y) & (~d7lhla0f70idm9pt) ) ? 
          (
            zwcbp7zqfei5xz ? {
              z0yhjfv_e0yaa2r,
              1'b1, 
              1'b0, 
              pydatzxqqi, 
              1'b1  
              } : 
            (o7hoht1pqz01v7 ? {
                   sco4chgj6vsbyoxn2j,
                   1'b1, 
                   1'b0, 
                   pydatzxqqi, 
                   1'b0  
               }: {  
                   n5_4v2cdhby2lv,
                   1'b1, 
                   1'b0, 
                   pydatzxqqi, 
                   1'b0  
                  }
               )  
          ) :
      (jukbv9h11v1o8cebnq & xv76y4hz81uw_gu & ( dn8riluj40uunvq5) & (~n703xx6o97u6y) & (~l89rffl8xklfzh4_e) ) ? 
          (
            zwcbp7zqfei5xz ? {
              d3hccrck1fl7jjf6,
              1'b0, 
              1'b1, 
              pydatzxqqi, 
              1'b1  
              } : 
            (vkyge0q4mfc5 ? {
                   tx81df88wvd5cnr5h5,
                   1'b0, 
                   1'b1, 
                   pydatzxqqi, 
                   1'b0  
               }: {  
                   wsufrwtxevzipw,
                   1'b0, 
                   1'b1, 
                   pydatzxqqi, 
                   1'b0  
                  }
               )  
          ) :
    
    
        (jukbv9h11v1o8cebnq & d7gc7q1qy89t05 & (~n703xx6o97u6y) & d7lhla0f70idm9pt ) ? {
                   uolend5_94trunxfp6p5,  
                   aw82i964do, 
                   y8_gkxsfle, 
                   pydatzxqqi, 
                   1'b0  
        } :
        (jukbv9h11v1o8cebnq & (~d7gc7q1qy89t05) & (~n703xx6o97u6y) & l89rffl8xklfzh4_e ) ? {
                   uolend5_94trunxfp6p5,  
                   aw82i964do, 
                   y8_gkxsfle, 
                   pydatzxqqi, 
                   1'b0  
        } :

          x76a6w0qgnegw5 ? {
                   uolend5_94trunxfp6p5,  
                   aw82i964do, 
                   y8_gkxsfle, 
                   pydatzxqqi, 
                   1'b0  
          }:{
                   n5_4v2cdhby2lv,
                   1'b1, 
                   1'b0, 
                   pydatzxqqi, 
                   1'b0  
                      } ;








  assign rjjrzh_tco6hcost86 = mxa77etukhs8o_5z6962l19;











  wire iynsf81xhrevxqe;
  wire rv1zybj1x67i66vbcgxki; 
  wire ij_6ovykpmdmrocvmn9udt; 

  wire kkbon6pdajchuxp;

  wire dd8pb3i1ec_uv5  ;
  wire s62ahm8e0we20r;
  qy_752rpwt4qqgs1gejira_te o61okcsx2t8btek447pam71bv (
    .j2f1_e0en      (pydatzxqqi),
    .aw82i964do      (aw82i964do), 
    .y8_gkxsfle      (y8_gkxsfle), 
    .azll7rq5fab5ou  (azll7rq5fab5ou   ),
    .dd8pb3i1ec_uv5  (dd8pb3i1ec_uv5  ),
    .s62ahm8e0we20r(s62ahm8e0we20r) 
  );

  wire h1zbk0qylhay7  ;

  assign ns0i7siujgkrghjpqv6 = (dbg_entry_taken_ena & kkbon6pdajchuxp)
                          | (r5sqfkv0bsgn5k6la & tg6dvyjbvr4lk8_esf1fjt & lpofewte8nxu7_o);
  
  
  
  wire nwl5lb3sma2kq78h = (~pydatzxqqi) & dd8pb3i1ec_uv5 & fh49u69v0he & (~dbg_entry_taken_ena);
  wire k0b98g3lj9szavjv9s = dbg_entry_taken_ena;
  wire xw8kra1vkkd21sk = nwl5lb3sma2kq78h | k0b98g3lj9szavjv9s;
  wire a5zxmoc94eq0hd6n26l = nwl5lb3sma2kq78h | (~k0b98g3lj9szavjv9s);
  ux607_gnrl_dfflr #(1) i624ky0quv0f1ys0ehgji (xw8kra1vkkd21sk, a5zxmoc94eq0hd6n26l, h1zbk0qylhay7, gf33atgy, ru_wi);

  wire ydz4q0fm5jvlahtf = h1zbk0qylhay7 | ((~pydatzxqqi) & dd8pb3i1ec_uv5 & jp82o1hu0f41an);

  wire ghbecqx593k3jui1e0b4 = (~pydatzxqqi) & s62ahm8e0we20r & fh49u69v0he & (~dbg_entry_taken_ena);
  wire rnjxs9qkjtqk_qq1 = r5sqfkv0bsgn5k6la;
  wire e6bcpnpomcng_r7x_ = ghbecqx593k3jui1e0b4 | rnjxs9qkjtqk_qq1;
  wire c5vih93g_pvfeeik = ghbecqx593k3jui1e0b4 | (~rnjxs9qkjtqk_qq1);
  ux607_gnrl_dfflr #(1) ihn82x5t9wvt9qdntb9i (e6bcpnpomcng_r7x_, c5vih93g_pvfeeik, lpofewte8nxu7_o, gf33atgy, ru_wi);



  
  
  
  
  wire vimkwxm8wxk8 = (~pydatzxqqi) & t5trf35s8vy & fh49u69v0he & (~dbg_entry_taken_ena) 
                      ;
  wire i26xa6gy6g6urr = dbg_entry_taken_ena;
  wire nu7da44khhl97840 = vimkwxm8wxk8 | i26xa6gy6g6urr;
  wire vtlq33kwc6mr = vimkwxm8wxk8 | (~i26xa6gy6g6urr);
  ux607_gnrl_dfflr #(1) itdw07c90jzyy75a (nu7da44khhl97840, vtlq33kwc6mr, iynsf81xhrevxqe, gf33atgy, ru_wi);

  wire a6m20tbmqogxskxqk2 = iynsf81xhrevxqe | ((~pydatzxqqi) & t5trf35s8vy & jp82o1hu0f41an);

 
  
  wire xgewxr6whza7hq;
  wire lptjbws412hnq = (~pydatzxqqi) & c4ughu0qm5sfai & rn2mt6nngsc9w5cz;
  wire avr43wmkvapsg = dbg_entry_taken_ena;
  wire cnfwj2f_p5i9haz = lptjbws412hnq | avr43wmkvapsg;
  wire m3ukybgp1gj8b = lptjbws412hnq & (~avr43wmkvapsg);
     
  ux607_gnrl_dfflr #(1) iq9qktodub_fa_3e16dx (cnfwj2f_p5i9haz, m3ukybgp1gj8b, xgewxr6whza7hq, dk2xhkj77a, ru_wi);

  wire nkyy10bp7u39xhsj = xgewxr6whza7hq | lptjbws412hnq;
  



  wire vjddv91epk5owamk = 1'b0;

  wire ietrigger_2dm_req_r;
  wire efxi850xz4_6cjr;
  wire sqv_vy58z6wkj_9z6; 
  wire dv16dpuz618c30za;
  wire xnziswi3rasuzqr; 

  wire hb3jz3_tihbfjg65curfxye;
 
  wire xa1l_abwrg85pdl8v8qfvrnz2 = (~pydatzxqqi) 
                       & efxi850xz4_6cjr
                       & gxmbdujixw2_0t7d527dq
                       ;
  
  wire n2jw5a4wxzlt258gkyog1e = dbg_entry_taken_ena;
  wire mxwbkm4d_h8wshcz93z8_ = xa1l_abwrg85pdl8v8qfvrnz2 | n2jw5a4wxzlt258gkyog1e;
  wire uov3bg1pa0nf503cyj_e64 = xa1l_abwrg85pdl8v8qfvrnz2 | (~n2jw5a4wxzlt258gkyog1e);
  ux607_gnrl_dfflr #(1) eatnpv3ny1j4dfja25m4qympm8 (mxwbkm4d_h8wshcz93z8_, uov3bg1pa0nf503cyj_e64, hb3jz3_tihbfjg65curfxye, gf33atgy, ru_wi);

  wire wvdg5kuzog0nneud5ocquvl4;
 
  wire fiqq_93fue_d4t0chcw3mn = (~pydatzxqqi) 
                       & sqv_vy58z6wkj_9z6
                       & gxmbdujixw2_0t7d527dq
                       ;
  
  wire nosya4fxy1b5hdx0ozknai_k3o = r5sqfkv0bsgn5k6la;
  wire hhiroca8wx2kd63havneej = fiqq_93fue_d4t0chcw3mn | nosya4fxy1b5hdx0ozknai_k3o;
  wire ovf6txzxn9gt_l8rpjjvbx9 = fiqq_93fue_d4t0chcw3mn | (~nosya4fxy1b5hdx0ozknai_k3o);
  ux607_gnrl_dfflr #(1) od5vjfmcjltc9_f1okjy15fokifh (hhiroca8wx2kd63havneej, ovf6txzxn9gt_l8rpjjvbx9, wvdg5kuzog0nneud5ocquvl4, gf33atgy, ru_wi);

  wire b0hxibua7idgqwtycep9;
 
  wire f_s51co7ag9qa0r65n0dt00 = (~pydatzxqqi) 
                       & dv16dpuz618c30za
                       & r5sqfkv0bsgn5k6la
                       ;
  
  wire jcrn6okn9qfl3103og38xx9m = dbg_entry_taken_ena;
  wire b1l46smcne7osj05_iqf3dwy = f_s51co7ag9qa0r65n0dt00 | jcrn6okn9qfl3103og38xx9m;
  wire k8vxwl3a697y4et4if7mds = f_s51co7ag9qa0r65n0dt00 | (~jcrn6okn9qfl3103og38xx9m);
  ux607_gnrl_dfflr #(1) qvlj3afmlft_mbfzqcygvd6mxgv (b1l46smcne7osj05_iqf3dwy, k8vxwl3a697y4et4if7mds, b0hxibua7idgqwtycep9, gf33atgy, ru_wi);

  wire jpp_xn78vvlrfu2ofdtlxm_4;
 
  wire r7o79i_n2yhrz7yc_zbd8p1 = (~pydatzxqqi) 
                       & xnziswi3rasuzqr
                       & r5sqfkv0bsgn5k6la
                       ;
  
  wire lxj25qm5rs2zmw6i0vhjxb1pz6e = r5sqfkv0bsgn5k6la;
  wire eo1gj6qt_gu_bdjckme3z60p = r7o79i_n2yhrz7yc_zbd8p1 | lxj25qm5rs2zmw6i0vhjxb1pz6e;
  wire nyhsikwoa5z8q4fc1pgc2lewgwn = r7o79i_n2yhrz7yc_zbd8p1 | (~lxj25qm5rs2zmw6i0vhjxb1pz6e);
  ux607_gnrl_dfflr #(1) r_m713fqirqeora7uqigfczhdz_ (eo1gj6qt_gu_bdjckme3z60p, nyhsikwoa5z8q4fc1pgc2lewgwn, jpp_xn78vvlrfu2ofdtlxm_4, gf33atgy, ru_wi);



  wire jgdzznlamq4mykbg3iszr = wvdg5kuzog0nneud5ocquvl4 | jpp_xn78vvlrfu2ofdtlxm_4;
  assign ietrigger_2dm_req_r   = hb3jz3_tihbfjg65curfxye   | b0hxibua7idgqwtycep9  ;

  assign usl0bxdbhf2_xj = jgdzznlamq4mykbg3iszr; 


  wire dbg_trig_req;
  wire dbg_exc2dbg_req;



    wire x6r5iqjhi4m5203iz8k = 1'b0;
  wire aoanpm_v6evzqd4 = nkyy10bp7u39xhsj       & (~x6r5iqjhi4m5203iz8k) ; 
  assign dbg_exc2dbg_req = vjddv91epk5owamk       & (~x6r5iqjhi4m5203iz8k) & (~nkyy10bp7u39xhsj) ;
  wire fk4wnf38_vuoydu  = ietrigger_2dm_req_r & (~x6r5iqjhi4m5203iz8k) & (~nkyy10bp7u39xhsj)  & (~vjddv91epk5owamk) ;
  wire eq9_qziyj0kl7v    = c5ewdqztjw9za            & (~x6r5iqjhi4m5203iz8k) & (~nkyy10bp7u39xhsj)  & (~vjddv91epk5owamk) & (~ietrigger_2dm_req_r) ;
  wire ftbwgnjeq_iu    = iynsf81xhrevxqe          & (~x6r5iqjhi4m5203iz8k) & (~nkyy10bp7u39xhsj)  & (~vjddv91epk5owamk) & (~ietrigger_2dm_req_r) & (~c5ewdqztjw9za);
  assign kkbon6pdajchuxp  = h1zbk0qylhay7        & (~x6r5iqjhi4m5203iz8k) & (~nkyy10bp7u39xhsj)& (~vjddv91epk5owamk) & (~ietrigger_2dm_req_r) & (~c5ewdqztjw9za) & (~iynsf81xhrevxqe);
  assign dbg_trig_req = ij_6ovykpmdmrocvmn9udt  & (~x6r5iqjhi4m5203iz8k) & (~nkyy10bp7u39xhsj)  & (~vjddv91epk5owamk) & (~ietrigger_2dm_req_r) & (~c5ewdqztjw9za) & (~iynsf81xhrevxqe) & (~h1zbk0qylhay7);
  wire kz5i_8mxfpdjge1u = rv1zybj1x67i66vbcgxki  & (~x6r5iqjhi4m5203iz8k) & (~nkyy10bp7u39xhsj)  & (~vjddv91epk5owamk) & (~ietrigger_2dm_req_r) & (~c5ewdqztjw9za) & (~iynsf81xhrevxqe) & (~h1zbk0qylhay7) & (~ij_6ovykpmdmrocvmn9udt) ;

  wire ez7p69p7r34w1cv4hspa9f  = a6m20tbmqogxskxqk2;
  wire u1z2rhoobjnpx2jl8rcm  = ydz4q0fm5jvlahtf;



  wire nuutbfpu8f4qqs5h3z  = pydatzxqqi;

  assign q7r68kfb621_p = cn7vi2ekbeqvap2074co5n33s | bkjtjv8qktytwklm1;

  assign bkjtjv8qktytwklm1 = (~nuutbfpu8f4qqs5h3z) & (
                                              dbg_trig_req
                                            | kz5i_8mxfpdjge1u
                                            );

  assign cn7vi2ekbeqvap2074co5n33s = (~nuutbfpu8f4qqs5h3z) & (

                                              x6r5iqjhi4m5203iz8k
                                            | eq9_qziyj0kl7v
                                            | dbg_exc2dbg_req
                                            | fk4wnf38_vuoydu
                                            | kkbon6pdajchuxp
                                            | aoanpm_v6evzqd4
                                            | ftbwgnjeq_iu
                                            );

  assign wlotcqomlz6de0sr4ukuhgbwpu3n = (~nuutbfpu8f4qqs5h3z) & (

                                              x6r5iqjhi4m5203iz8k
                                            | eq9_qziyj0kl7v
                                            | dbg_exc2dbg_req
                                            | fk4wnf38_vuoydu
                                            | u1z2rhoobjnpx2jl8rcm 
                                            | aoanpm_v6evzqd4
                                            | ez7p69p7r34w1cv4hspa9f 
                                            );











  wire   oi9ysx1fe1e6o6ozcfe = s5f_36xvqrtq7 | (~aw82i964do);
  assign d7lhla0f70idm9pt = (u5a92wwchl7sg75h & ((~oi9ysx1fe1e6o6ozcfe) 
                                              | h7fseh5_df0hbx) 
                                              );

  wire   h84s5qlh46hifajxj9n = (w632tcbtqncn6 & (~aw82i964do) & y8_gkxsfle) | ((~aw82i964do) & (~y8_gkxsfle));
  








  assign l89rffl8xklfzh4_e =  u5a92wwchl7sg75h & 
                            (
                                 (~h84s5qlh46hifajxj9n) 
                               | h7fseh5_df0hbx 
                            );

  wire zsg9re2v0e3y4ik5bekzg2 =  t5trf35s8vy ? (~ozwene1gdpatk6g) : 1'b0;




  wire lvgwfqq1fbs  = pydatzxqqi | zsg9re2v0e3y4ik5bekzg2 | cwwkpmk260lrt;

  wire c64nh23l7  = pydatzxqqi | zsg9re2v0e3y4ik5bekzg2;

  
  
  
  
  
  
  
  
  
  wire gz7m6d_jp54  = pydatzxqqi | zsg9re2v0e3y4ik5bekzg2 | 
                   (
                       d7gc7q1qy89t05 ?       
                      ((~oi9ysx1fe1e6o6ozcfe)   
                     & (~d7lhla0f70idm9pt)) :   
                       (xv76y4hz81uw_gu       

                     & (~h84s5qlh46hifajxj9n)   
                     & (~l89rffl8xklfzh4_e)   
                   ))
                   ;

  wire ym57gq2j35jz7   = (v3ne7glf8d8   & aw0hbwfkx3f63s); 
  wire tqt7qc7ciiqou6m   = (lt3v_fm0ipu   & mfzl2fqml69hx); 
  wire q89equ1ce16bt5   = (x6eltyshbu5   & siifnhwgancn8);
  wire k45zf0g_j1rcvg1d72 = (v9dnbgjy6c0vf & u83p4flbuvkqt26z); 
  wire cgx9nttfofebj23k4  = (hmzw4exmjn8k921c  & tvglhc8o_izdq );
  assign s74_qw0a41imkgkdcsf0rdhta = ym57gq2j35jz7 | tqt7qc7ciiqou6m | q89equ1ce16bt5 | k45zf0g_j1rcvg1d72 | cgx9nttfofebj23k4;

  wire t9sjp9l7wcp8ii   = (ezl3jzeqhltgj7h   & ai169tbqp4seb3); 
  wire o2f1c5d_jgdk_65   = (i9xvsmm45fp0f58   & yw4o4kdms07_32); 
  wire upjfj9ci9jnkqdc   = (w529wbj853   & b0zz_ornhz010);
  assign tf2ird6le5az6cmue2y6_ = t9sjp9l7wcp8ii | o2f1c5d_jgdk_65 | upjfj9ci9jnkqdc;

  wire ztqjcc14uirynsx = dn8riluj40uunvq5 ? fcjh1nct4r : (
                   s74_qw0a41imkgkdcsf0rdhta   
                 | tf2ird6le5az6cmue2y6_   
                 );

  assign n703xx6o97u6y = (~lvgwfqq1fbs) & feq1g7m2cy1erl; 
  wire qlc_ro_yd0vr   = (~gz7m6d_jp54) & ztqjcc14uirynsx;
  wire ptj40008gk    = (~c64nh23l7) & uc5qxb4d2b28ye5; 


  wire a7_9q7k_ywckdao = (d7lhla0f70idm9pt & h7fseh5_df0hbx);
  assign z5sexv2 = a7_9q7k_ywckdao ? (ptj40008gk | n703xx6o97u6y) :

                                  (qlc_ro_yd0vr | n703xx6o97u6y);


  assign bet3r1ns0njrwezuu = z5sexv2; 


  wire [64-1:0] l69ubuy_qz;

  assign k3cmpuswk7in0u4 = l69ubuy_qz[11:0];

  assign l69ubuy_qz[64-1] = n703xx6o97u6y ? 1'b0 : 1'b1;
  assign l69ubuy_qz[64-2:12] = {(64-13){1'b0}};
  assign l69ubuy_qz[11:0]  =  
                           n703xx6o97u6y    ? {w2fpnf5fg1byp6 ? 12'hFFF : 12'h001} :  
                           dn8riluj40uunvq5 ? {{12-10{1'b0}},b4lwcgm6l21pi} :
                           (
                           cgx9nttfofebj23k4  ? 12'd18 :
                           k45zf0g_j1rcvg1d72 ? 12'd16 :
                           ym57gq2j35jz7   ? 12'd11 :  
                           tqt7qc7ciiqou6m   ? 12'd3  :  
                           q89equ1ce16bt5   ? 12'd7  :  
                           t9sjp9l7wcp8ii   ? 12'd9  :  
                           o2f1c5d_jgdk_65   ? 12'd1  :  
                           upjfj9ci9jnkqdc   ? 12'd5  :  
                                         12'b0);










  wire zv3yqd89ktm50jultzaxa;
  wire q3xnqi83t13ql96xa2lnj9e;
  wire l6t30n2cfj_wzt549dhwjl8x3 = klz7l8_75czqn63zb & (~q3xnqi83t13ql96xa2lnj9e);
  wire azsxdi_wqzat2q = (
                      (aw82i964do ? (~zbac123pv78sbz3) : y8_gkxsfle ? (~z4e_m564fxae0kpbjr) :(~hixy2y36a1pn0)) 

                     | pydatzxqqi
                     );
  assign jbod2vk5w_ts8f0pmlikw9b7 = (l6t30n2cfj_wzt549dhwjl8x3 & (azsxdi_wqzat2q));
  wire mp4bdzd27nl7gsjskmzri3cgojs = jbod2vk5w_ts8f0pmlikw9b7
                                | zv3yqd89ktm50jultzaxa
                                ;


  wire of8jbhv7emsqm5tw2qqov4t = l6t30n2cfj_wzt549dhwjl8x3 & (~azsxdi_wqzat2q);

  assign rv1zybj1x67i66vbcgxki = p7rj2v1hvh0nab6ei & of8jbhv7emsqm5tw2qqov4t;
  assign btwmhh91h50d5flgwx4o6pwu = rv1zybj1x67i66vbcgxki;





  wire c7o1ubuxo5fr_pgdh4pfb = (~pydatzxqqi) & 
                    ( 
                    | gnn94t_31a_j59f483ym5f68sb
                    | wkyo2nrlaz9sq3m1chcysnofuenz
                    );
  assign zv3yqd89ktm50jultzaxa = (~pydatzxqqi) & 
                    ( 
                    | zb322_7v29pmo4jvmvow3qi8
                    | vmkmkz3cm8cgbet959d4pw_0ti
                    );
  assign ij_6ovykpmdmrocvmn9udt = p7rj2v1hvh0nab6ei & c7o1ubuxo5fr_pgdh4pfb;




  assign q3xnqi83t13ql96xa2lnj9e = 
            ( u3qmzjrm6inkod3m3ghp 
            | qsn_nfmbj97wz1r3s59t2 
            | uuvo0ter1b1y6j1xfc 
            | hjysp7ahvean99t41k89pt 
            | ggvuzlnuknlvg4a50n4hy7ok 

            | j6g8r7rblr88am07jc3i5
            | iq2e_b4p5qjp2ryy5sktbl6kd0  
            | om206h86cfrb69iqc9pzq3fq1  
            | yk85cwkls6hcvp4_g70j2  
            | cj2z8_7e4hw2s1u6mhckmpm4i  
            | rpt826mhm0kwty9qlty6rt1  
            | nqoqg40hg82wgdbsfubvu4fg
            | hcx0jkab_j87_6j7phxnsz
            | t0zuyah73tpfg_dtxy56ug9ej
            );

  assign mp89sr5uys176dofb6r = 
            ( q3xnqi83t13ql96xa2lnj9e 
            | mp4bdzd27nl7gsjskmzri3cgojs
            ) & (~c7o1ubuxo5fr_pgdh4pfb);











  wire i8gj0xp7yt1_pz2mb5mvqdemh    = m0ugsckv2bvgxdilc4lz & fe8u85vitwnfnuszhl;
  wire wbletfvgmj22tsfe41_moe80ay = m0ugsckv2bvgxdilc4lz & stx6pefjqd_oqqg5gej9;


  wire shf9huvtyxgf86qaw8npjh6mvfdk13 = om206h86cfrb69iqc9pzq3fq1 
                                  & (~yk85cwkls6hcvp4_g70j2)
                                  & (~cj2z8_7e4hw2s1u6mhckmpm4i)
                                  ;

  wire yyd7bchda2at_6ombe9lj_7yb      = (m0ugsckv2bvgxdilc4lz & mp4bdzd27nl7gsjskmzri3cgojs);
  wire o5rg5rzrjydokq_ibohf3u3xc12       = (m0ugsckv2bvgxdilc4lz & j6g8r7rblr88am07jc3i5);
  wire mg31i1mqkc18cng71t81u4am419lz6 = (m0ugsckv2bvgxdilc4lz & iq2e_b4p5qjp2ryy5sktbl6kd0);
  wire k6_34kl5n41c6xlwcq130vu4g3dp0mq_  = (m0ugsckv2bvgxdilc4lz & shf9huvtyxgf86qaw8npjh6mvfdk13);
  wire lewchw0ezo4jt8v22yrw8w56kl4bfb_  = (m0ugsckv2bvgxdilc4lz & yk85cwkls6hcvp4_g70j2);
  wire eqywl573zop4xk9qcqxsg8hofl60nlh31  = (m0ugsckv2bvgxdilc4lz & cj2z8_7e4hw2s1u6mhckmpm4i);
  wire f1zgxm6uf8gjzesiiqgbeeey3j409   = (m0ugsckv2bvgxdilc4lz & rpt826mhm0kwty9qlty6rt1 & (~om206h86cfrb69iqc9pzq3fq1));
  wire uxe2yyr6wh0nuxu79x89lzay9r     = t0zuyah73tpfg_dtxy56ug9ej & 
                                        (
                                           1'b1 
                                         & ~nqoqg40hg82wgdbsfubvu4fg
                                         & ~hcx0jkab_j87_6j7phxnsz
                                        )
                                        ;
  wire wh5ybgwfpmtfo57_js_ngl7k98u5elwp2  = (m0ugsckv2bvgxdilc4lz & fi9wz0kme0ey_bxavdqx_9 & uxe2yyr6wh0nuxu79x89lzay9r);
  wire zha0bsafnp8bvf2f0hpach3w54b41ix  = (m0ugsckv2bvgxdilc4lz & tmhbzyv2b510vt_9qkb16hdwa & uxe2yyr6wh0nuxu79x89lzay9r);
  wire fds7hg2n4wmvmzq9ld13kq5gpv4t8k  = (m0ugsckv2bvgxdilc4lz & fi9wz0kme0ey_bxavdqx_9 & nqoqg40hg82wgdbsfubvu4fg);
  wire xgtje2gxllohikwc3j_ql2fchhhe3hl  = (m0ugsckv2bvgxdilc4lz & tmhbzyv2b510vt_9qkb16hdwa & nqoqg40hg82wgdbsfubvu4fg);
  wire i0_i17y0yq11bismg5yaqrk1h4wi9iad9  = (m0ugsckv2bvgxdilc4lz & fi9wz0kme0ey_bxavdqx_9 & hcx0jkab_j87_6j7phxnsz);
  wire z0heerx232q93x2y8ewx75q0swerv  = (m0ugsckv2bvgxdilc4lz & tmhbzyv2b510vt_9qkb16hdwa & hcx0jkab_j87_6j7phxnsz);


  wire adi1tne59q4fj9gpvzopu1cjh9peva    = (i8gj0xp7yt1_pz2mb5mvqdemh    & u3qmzjrm6inkod3m3ghp);
  wire rxvfzl0wv05oaumybran7wvqdf3ww0     = (i8gj0xp7yt1_pz2mb5mvqdemh    & qsn_nfmbj97wz1r3s59t2);
  wire b08xw227fs65cv4t3ljg_650u5g5wn     = (i8gj0xp7yt1_pz2mb5mvqdemh    & uuvo0ter1b1y6j1xfc);
  wire bj2wyn7rse20tace3s37xhus8h0ppn_aq = (wbletfvgmj22tsfe41_moe80ay & u3qmzjrm6inkod3m3ghp);
  wire jlva726ka65z9up1cmfrkh0wz38dvcv7  = (wbletfvgmj22tsfe41_moe80ay & qsn_nfmbj97wz1r3s59t2);
  wire smlrsduaqesh4yg4au3gqaeqxrvw1hi  = (wbletfvgmj22tsfe41_moe80ay & uuvo0ter1b1y6j1xfc);
  wire p5cdr4hplss042ubzgyi34btkaz6g78   = (wmeyhl03a273zu2s7qupf5h & cd4v4c_rw906kt5 & hv4wuttuo9jk_cqa8sxqwt);
  wire mh2wtnrxhqy03pbrrjvuw15hhr6sj2   = (wmeyhl03a273zu2s7qupf5h & idat72abxke4z9s & hv4wuttuo9jk_cqa8sxqwt);
  wire qa7h91vqmai0_6l67a0ohi23s7wh5qm8s   = (wmeyhl03a273zu2s7qupf5h & cd4v4c_rw906kt5 & ac8_dky9fhpbsxu0b9t88ag8);
  wire c9zdhvpduvc3sxet_rckpqh6raspp6m   = (wmeyhl03a273zu2s7qupf5h & idat72abxke4z9s & ac8_dky9fhpbsxu0b9t88ag8);
  wire ezo9aq6vqzzlj4mxue54 = xo1uoocz53uginn8n & evla4t4m7kx62w598l;
  wire kl75_su5ts4ncxua = xo1uoocz53uginn8n & oxberxo5xs4cqy454m0;

  wire hrjpps0u1el6sdpkvumeech9 = 
                     adi1tne59q4fj9gpvzopu1cjh9peva    
                   | rxvfzl0wv05oaumybran7wvqdf3ww0     
                   | bj2wyn7rse20tace3s37xhus8h0ppn_aq 
                   | jlva726ka65z9up1cmfrkh0wz38dvcv7;

  wire ypb4xehjnrzxssq3i3qzg75p15z9y = 
                     1'b0
                   | b08xw227fs65cv4t3ljg_650u5g5wn 
                   | smlrsduaqesh4yg4au3gqaeqxrvw1hi
                   ;


  wire blq8dmuhwtno2_o2glw38jo154fv = 
                     wh5ybgwfpmtfo57_js_ngl7k98u5elwp2
                   | zha0bsafnp8bvf2f0hpach3w54b41ix
                   | fds7hg2n4wmvmzq9ld13kq5gpv4t8k
                   | xgtje2gxllohikwc3j_ql2fchhhe3hl
                   ;

  wire ua77845ub9_kdh4dp3iap0etawtvqjpv44so = 
                     1'b0
                   | i0_i17y0yq11bismg5yaqrk1h4wi9iad9
                   | z0heerx232q93x2y8ewx75q0swerv
                   ;

  wire uti0ee1pemfxsobkm9837i3wizzzlw29mxa = 
                     1'b0
                   ;

  wire x62kevhmegzodop4ziik6er_k1z1j = 
                     p5cdr4hplss042ubzgyi34btkaz6g78   
                   | mh2wtnrxhqy03pbrrjvuw15hhr6sj2;

  wire b09b5lyi_s2bcv6vxim = (k6_34kl5n41c6xlwcq130vu4g3dp0mq_ | lewchw0ezo4jt8v22yrw8w56kl4bfb_);

  wire ioenbox_g6rd3jl1hjw_ = (p5cdr4hplss042ubzgyi34btkaz6g78 
                         |  qa7h91vqmai0_6l67a0ohi23s7wh5qm8s   
                         |  rxvfzl0wv05oaumybran7wvqdf3ww0
                         | wh5ybgwfpmtfo57_js_ngl7k98u5elwp2  
                         | fds7hg2n4wmvmzq9ld13kq5gpv4t8k  
                         );

  wire i33_fq2xr9qks17gti3r = (mh2wtnrxhqy03pbrrjvuw15hhr6sj2 
                          |  c9zdhvpduvc3sxet_rckpqh6raspp6m   
                          |  jlva726ka65z9up1cmfrkh0wz38dvcv7
                          |  hjysp7ahvean99t41k89pt       
                          | zha0bsafnp8bvf2f0hpach3w54b41ix  
                          | xgtje2gxllohikwc3j_ql2fchhhe3hl  
                          );

  wire l_wc20qa_jrwxs8im1c =  eqywl573zop4xk9qcqxsg8hofl60nlh31
                         ;
  wire iio4ar1e8jmmhmt = b08xw227fs65cv4t3ljg_650u5g5wn
                         |  i0_i17y0yq11bismg5yaqrk1h4wi9iad9  
                         ;
  wire b6ezo9ij_3xanedr = smlrsduaqesh4yg4au3gqaeqxrvw1hi
                          |  ggvuzlnuknlvg4a50n4hy7ok       
                          |  z0heerx232q93x2y8ewx75q0swerv
                          ;



  wire [64-1:0] hh49o83xz9_uu;
  assign hh49o83xz9_uu[64-1:10] = {(64-10){1'b0}};

  wire qd98gcnboxkmqcnqfei;
  assign {qd98gcnboxkmqcnqfei, hh49o83xz9_uu[9:0]}  = 
      mg31i1mqkc18cng71t81u4am419lz6 ?                       {~r4bs4k_53n5wp[0], 10'd0} 
    : b09b5lyi_s2bcv6vxim ?                                   {~r4bs4k_53n5wp[1], 10'd1} 
    : f1zgxm6uf8gjzesiiqgbeeey3j409  ?                        {~r4bs4k_53n5wp[2], 10'd2} 
    : (yyd7bchda2at_6ombe9lj_7yb | tg6dvyjbvr4lk8_esf1fjt) ? {~r4bs4k_53n5wp[3], 10'd3} 
    : adi1tne59q4fj9gpvzopu1cjh9peva ?                        {~r4bs4k_53n5wp[4], 10'd4} 
    : ioenbox_g6rd3jl1hjw_ ?                                    {~r4bs4k_53n5wp[5], 10'd5} 
    : bj2wyn7rse20tace3s37xhus8h0ppn_aq ?                     {~r4bs4k_53n5wp[6], 10'd6} 
    : i33_fq2xr9qks17gti3r ?                                   {~r4bs4k_53n5wp[7], 10'd7} 
    : (o5rg5rzrjydokq_ibohf3u3xc12 & (~aw82i964do) & (~y8_gkxsfle)) ?   {~r4bs4k_53n5wp[8], 10'd8} 
    : (o5rg5rzrjydokq_ibohf3u3xc12 & y8_gkxsfle) ?                  {~r4bs4k_53n5wp[9], 10'd9} 
    
    : (o5rg5rzrjydokq_ibohf3u3xc12 & aw82i964do) ?                  {~r4bs4k_53n5wp[11], 10'd11} 
    : l_wc20qa_jrwxs8im1c ?                                     {~r4bs4k_53n5wp[12], 10'd12} 
    : iio4ar1e8jmmhmt ?                                      {~r4bs4k_53n5wp[13], 10'd13} 
    : b6ezo9ij_3xanedr ?                                     {~r4bs4k_53n5wp[15], 10'd15} 
    : ezo9aq6vqzzlj4mxue54 ?                                     {1'b1, 10'd32}
    : kl75_su5ts4ncxua ?                                     {1'b1, 10'd33}
    : {1'b1, 10'h0};

  assign av15ikbsl_f = aw82i964do | qd98gcnboxkmqcnqfei;
  assign dbk9rh15g1 = ~av15ikbsl_f;               




  vx6hu6m3c9ub1xbqu6okmcqh6_ msz7p2tfzyrbv9t3fxmvsz_slae(
    .dn8riluj40uunvq5(dn8riluj40uunvq5), 
    .j2f1_e0en       (pydatzxqqi),
    .aw82i964do       (aw82i964do),
    .y8_gkxsfle       (y8_gkxsfle),
    .hh49o83xz9_uu   (5'b0),
    .g1fa4tixb       (l69ubuy_qz[9:0]),
  
    .lmu064oe20     (1'b0),
    .qemnpyvmwrt      (1'b1),
  
    .n6a0r_0zddzrme8   (n6a0r_0zddzrme8),
    .azll7rq5fab5ou   (azll7rq5fab5ou),
  
    .coeuovgdaw1  (efxi850xz4_6cjr),
    .o_gen1so7__xgr3pw2(sqv_vy58z6wkj_9z6) 
  );

  vx6hu6m3c9ub1xbqu6okmcqh6_ nyexm0e82y2lo03u6_i4ix63(
    .dn8riluj40uunvq5(1'b0), 
    .j2f1_e0en       (pydatzxqqi),
    .aw82i964do       (aw82i964do),
    .y8_gkxsfle       (y8_gkxsfle),
    .hh49o83xz9_uu   (hh49o83xz9_uu[4:0]),
    .g1fa4tixb       (10'b0),
  
    .lmu064oe20     (1'b1),
    .qemnpyvmwrt      (1'b0),
  
    .n6a0r_0zddzrme8   (n6a0r_0zddzrme8),
    .azll7rq5fab5ou   (azll7rq5fab5ou),
  
    .coeuovgdaw1  (dv16dpuz618c30za),
    .o_gen1so7__xgr3pw2(xnziswi3rasuzqr) 
  );






















  wire n8nhee4fy2dxtog_fbfv73 = cxij98yy3k4hy34_9o;

  wire stl2dyg;
  assign {stl2dyg,wtd_nuaeb_mpye} = 
               (x62kevhmegzodop4ziik6er_k1z1j) ? r_8f7p3tznijza5y03ko : 
               (yyd7bchda2at_6ombe9lj_7yb & zv3yqd89ktm50jultzaxa & vmkmkz3cm8cgbet959d4pw_0ti) ? {{64+1-64{1'b0}},n7orghfl8x_7wsaisuhpw9o} :   
               (yyd7bchda2at_6ombe9lj_7yb & zv3yqd89ktm50jultzaxa & zb322_7v29pmo4jvmvow3qi8) 
                                                                    ? {{64+1-64{1'b0}},wql66zm9cb_1pzbk} :   
               ( tg6dvyjbvr4lk8_esf1fjt) 
                                                                    ? {{64+1-64{1'b0}},uolend5_94trunxfp6p5} :   
               mg31i1mqkc18cng71t81u4am419lz6 ? {{64+1-64{1'b0}},wql66zm9cb_1pzbk} :
               (b09b5lyi_s2bcv6vxim & lewchw0ezo4jt8v22yrw8w56kl4bfb_) ? {{64+1-64{1'b0}},{lovkp0eqfnxtb7[64-1:3],3'b0}} :
               (b09b5lyi_s2bcv6vxim & k6_34kl5n41c6xlwcq130vu4g3dp0mq_) ? (

                                            {{64+1-64{1'b0}},{lovkp0eqfnxtb7[64-1:3],3'b0}}) :
               f1zgxm6uf8gjzesiiqgbeeey3j409 ? (fof2qu1zf51j1nid7vs4 ? {{64+1-32{1'b0}},skcwu9hiw7zl59wu} : {{64+1-16{1'b0}},skcwu9hiw7zl59wu[15:0]}) :
               hrjpps0u1el6sdpkvumeech9    ? {{64+1-64{1'b0}},n7orghfl8x_7wsaisuhpw9o} : 
               hjysp7ahvean99t41k89pt ? {{64+1-64{1'b0}}, lt3biawnyshgr5rw4q5chcg6u7rc} : 
               ggvuzlnuknlvg4a50n4hy7ok ? {{64+1-64{1'b0}}, lt3biawnyshgr5rw4q5chcg6u7rc} : 
               blq8dmuhwtno2_o2glw38jo154fv ? {{64+1-64{1'b0}},sq0y2gv0vwpq_6ckk9b89gybz} : 
               uti0ee1pemfxsobkm9837i3wizzzlw29mxa ? {{64+1-64{1'b0}},sq0y2gv0vwpq_6ckk9b89gybz} : 
               l_wc20qa_jrwxs8im1c ? {{64+1-64{1'b0}},{lovkp0eqfnxtb7[64-1:3],3'b0}} :
               ypb4xehjnrzxssq3i3qzg75p15z9y ? {{64+1-64{1'b0}},n7orghfl8x_7wsaisuhpw9o} : 
               ua77845ub9_kdh4dp3iap0etawtvqjpv44so ? {{64+1-64{1'b0}},sq0y2gv0vwpq_6ckk9b89gybz} : 
               {64+1{1'b0}};







  assign uolend5_94trunxfp6p5 = qwcb6hcmvfqmf032z ? cvvsn7xc8qg5uk : k84xk2u4clez; 
  assign elth4vimq_j = (oyiml9jn3w6vt88yja9asjx) ? wql66zm9cb_1pzbk : uolend5_94trunxfp6p5;




  assign xd66pm611ai1dg = r5sqfkv0bsgn5k6la ? hh49o83xz9_uu : l69ubuy_qz;




  assign xv08lot3vi9dag4vs0 = r9uxubpl2h2alj1q;

  assign ew08uu2kn2p9e11s[64-1:3] = {64-3{1'b0}};

  wire hhe88a661c3sax8g = sf0uuehfhfa & (
                          (b09b5lyi_s2bcv6vxim & 1'b0) | 
                          (ioenbox_g6rd3jl1hjw_ & 1'b0) |
                          (i33_fq2xr9qks17gti3r & 1'b0) 
                         ) 
                         ;

  wire j8zx4rgi5245pulk = sf0uuehfhfa & (
                          (b09b5lyi_s2bcv6vxim & lewchw0ezo4jt8v22yrw8w56kl4bfb_) | 
                          (ioenbox_g6rd3jl1hjw_ &  
                          (rxvfzl0wv05oaumybran7wvqdf3ww0 
                          | qa7h91vqmai0_6l67a0ohi23s7wh5qm8s
                          | fds7hg2n4wmvmzq9ld13kq5gpv4t8k
                                                     ))
                         | (i33_fq2xr9qks17gti3r & (jlva726ka65z9up1cmfrkh0wz38dvcv7 | c9zdhvpduvc3sxet_rckpqh6raspp6m
                            | xgtje2gxllohikwc3j_ql2fchhhe3hl  
                          ))
                        ) 
                      ;

  wire f3j12c67yn5ieysupy = sf0uuehfhfa & ( 
                          (b09b5lyi_s2bcv6vxim & k6_34kl5n41c6xlwcq130vu4g3dp0mq_ & (~lewchw0ezo4jt8v22yrw8w56kl4bfb_)) | 
                          (
                           ioenbox_g6rd3jl1hjw_ & 
                           ( 
                              ( p5cdr4hplss042ubzgyi34btkaz6g78
                              ) |
                              (wh5ybgwfpmtfo57_js_ngl7k98u5elwp2 & (~fds7hg2n4wmvmzq9ld13kq5gpv4t8k )) |
                              1'b0
                           )
                          ) |
                         (
                          i33_fq2xr9qks17gti3r & 
                          ( 
                             ( mh2wtnrxhqy03pbrrjvuw15hhr6sj2 
                              ) |
                             (zha0bsafnp8bvf2f0hpach3w54b41ix & (~xgtje2gxllohikwc3j_ql2fchhhe3hl )) | 
                              1'b0
                           )
                          )
                        ) 
                      ;


  wire a6cehuwu_3eui24c = sf0uuehfhfa & ( 
                          (b09b5lyi_s2bcv6vxim & 1'b0) | 
                          (ioenbox_g6rd3jl1hjw_ &  1'b0) |
                          (ioenbox_g6rd3jl1hjw_ &  1'b0) 
                         )
                         ;


  wire gcg_d8r4krsp1ebpm2mx = sf0uuehfhfa & ( 
                          (b09b5lyi_s2bcv6vxim & 1'b0) | 
                          (ioenbox_g6rd3jl1hjw_ &  1'b0) |
                          (b6ezo9ij_3xanedr   & ggvuzlnuknlvg4a50n4hy7ok) |
                          (i33_fq2xr9qks17gti3r & hjysp7ahvean99t41k89pt) 
                         )
                         ;


  wire ti4m6j9qpzikzczugji = sf0uuehfhfa & ( 
                          (l_wc20qa_jrwxs8im1c & eqywl573zop4xk9qcqxsg8hofl60nlh31)   | 
                          (iio4ar1e8jmmhmt  & b08xw227fs65cv4t3ljg_650u5g5wn)    |
                          (b6ezo9ij_3xanedr & smlrsduaqesh4yg4au3gqaeqxrvw1hi) |
                          (iio4ar1e8jmmhmt  & i0_i17y0yq11bismg5yaqrk1h4wi9iad9)   |
                          (b6ezo9ij_3xanedr & z0heerx232q93x2y8ewx75q0swerv)   |
                          (1'b0)                                                
                         )
                         ;


  wire lhfuupl5abhc7ovg = sf0uuehfhfa & ( 
                          (1'b0)                                                 
                         )
                         ;

  assign ew08uu2kn2p9e11s[3-1:0] = 
                     hhe88a661c3sax8g ? 3'd0 :
                     j8zx4rgi5245pulk ? 3'd1 :
                     f3j12c67yn5ieysupy ? 3'd2 :
                     a6cehuwu_3eui24c ? 3'd3 : 
                     gcg_d8r4krsp1ebpm2mx ? 3'd4 : 
                     ti4m6j9qpzikzczugji ? 3'd5 : 
                     lhfuupl5abhc7ovg ? 3'd6 : 
                                        3'd0 ;


  assign if5jz8qk0aqefy3v35o = 1'b0;

  assign mtc04rctrfyb[64-1:5] = {64-5{1'b0}};

  assign mtc04rctrfyb[5-1:0] = 5'b0
                                               | frfbo512g1_94ncrem_be859f
                                               ;




  assign jlud6jeuxe0espga     = (~pydatzxqqi) & (
                                (gxmbdujixw2_0t7d527dq & d7gc7q1qy89t05)  
                              | (r5sqfkv0bsgn5k6la & av15ikbsl_f )
                              | (z1ri4yxi78_p8hx8y  & gvvhhfwk9lgdcu  )
                          );
  assign sf0uuehfhfa   = r5sqfkv0bsgn5k6la;
  assign hvy2cpsp75f3    = gxmbdujixw2_0t7d527dq;
  assign z35xlcc6bt4    = z1ri4yxi78_p8hx8y;
  assign k3z202os   = vj6p6j6avq664060js8d_wit_7a;

  assign r9uxubpl2h2alj1q   = jlud6jeuxe0espga 
                             ;

  assign x7eg618xaszd4f21cl_g = jlud6jeuxe0espga & n8nhee4fy2dxtog_fbfv73;

  assign qeb3z0x5 =



               dbg_exc2dbg_req ? pldoasxyzlvx2
               : oyiml9jn3w6vt88yja9asjx ? wql66zm9cb_1pzbk : uolend5_94trunxfp6p5;
  assign ibhfuwrztbm8p4gg = dbg_entry_taken_ena;

  wire r6xevat8rjhff6rghc;


  assign b7g_vsn0zoewh6g1 = r6xevat8rjhff6rghc;
  assign onnv64ydiajl = aw82i964do ? 2'b11 : y8_gkxsfle  ? 2'b01 : 2'b00;       

  assign r6xevat8rjhff6rghc = dbg_entry_taken_ena;
  wire i80iwlprhf60uuod6v = jw4fsjecr0u919fr7;
  wire [2:0] gvnov11imobkfjf4 = 






                              aoanpm_v6evzqd4 ? 3'd5 : 
                              eq9_qziyj0kl7v  ? 3'd3 : 
                              ftbwgnjeq_iu ? 3'd4 :
                              fk4wnf38_vuoydu ? 3'd2 :
                              kkbon6pdajchuxp ? 3'd2 :
                              dbg_trig_req ? 3'd2 : 


                              (kz5i_8mxfpdjge1u | dbg_exc2dbg_req) ? 3'd1 : 
                                             3'd0;

  assign osv2437qj_3nuf = r6xevat8rjhff6rghc | i80iwlprhf60uuod6v;
  assign i8_5wt0vppx = r6xevat8rjhff6rghc ? gvnov11imobkfjf4 : 3'd0;


  assign d7gc7q1qy89t05 = (dn8riluj40uunvq5 ? jqsukc5b5drcc1e78 : s74_qw0a41imkgkdcsf0rdhta);
  assign xv76y4hz81uw_gu = (dn8riluj40uunvq5 ? gnn46rd7vvofruqij : tf2ird6le5az6cmue2y6_);
  assign z2g63deibg1b1quqr     = (~pydatzxqqi) & (
                                (gxmbdujixw2_0t7d527dq & (~d7gc7q1qy89t05) & xv76y4hz81uw_gu)  
                              | (r5sqfkv0bsgn5k6la & dbk9rh15g1 )
                              | (z1ri4yxi78_p8hx8y  & (~gvvhhfwk9lgdcu)  )
                          );
  assign p5jpgn4rvarpo = elth4vimq_j;
  assign dhjwho76fa8hqc   = z2g63deibg1b1quqr; 
  assign u25pqekq4df       = xd66pm611ai1dg; 
  assign icauf4l_12_c2xkj53lf  = dhjwho76fa8hqc;     
  assign xel6gw173w5x0      = ew08uu2kn2p9e11s;
  
  assign e_z6d7r9kxqg32te = 1'b0;     
  assign v8ydjtlz16x9tx     = mtc04rctrfyb;
  assign u_ufp_wg29ieoklxxz1 = z2g63deibg1b1quqr & n8nhee4fy2dxtog_fbfv73;
  assign tlgcdv86voe9     = wtd_nuaeb_mpye;









  assign o2qkf90r783 = a7_9q7k_ywckdao ? cxij98yy3k4hy34_9o : 1'b1;


  assign av1w8ld09cfofn = fh49u69v0he | cxij98yy3k4hy34_9o;


  assign im2b5l0h98avl6t4sj = r5sqfkv0bsgn5k6la | z1ri4yxi78_p8hx8y; 


  assign bw65wl7fvekfymd8vqx = gxmbdujixw2_0t7d527dq;


  assign pecbpcoa04vq = xd66pm611ai1dg;


  assign tb_snaxyfs = wtd_nuaeb_mpye;



  assign zc4mldgm25r = oyiml9jn3w6vt88yja9asjx ? wql66zm9cb_1pzbk : glime27x19feqrvvsa2nmeh5f ? uolend5_94trunxfp6p5 : wql66zm9cb_1pzbk;


  assign d23wb5yh1iyvf = skcwu9hiw7zl59wu;

  assign cy3nuhzm_v2p73mt = z2574r4ajgr7u7mtpb_wpetx;

  assign fvqwdz2hdbb = ij7ql6t124xbofcx;


  assign srim3bfnzhve = aw82i964do ? 2'b11 : y8_gkxsfle ? 2'b01 : 2'b00;


  assign e9u0rtvt8jrygyc8s = r2ovgzxgcrqk7dmnynz6j1zh_61qmz & (~se2buoxmq91dbic3y2m5hu); 



endmodule                                      






















module ybdbqemjrr2kv71i(
  input  rnx27onf2lbe,
  input  af5qc04tmn51e4u2h1z,

  
  
  
  
  input  mt0f3958vekbx9, 
  output x9a3z87q3adhgofd, 
  input  [4-1:0] lefkd05cxbpmfb,
  input  [64-1:0] wvg6yggd3_ngr,
  input  [64-1:0] fvamtne5n7,
  input  [64-1:0] w6fv3puuz49wu,

  input  [3-1:0] ahi4ptho3r9,
  input  tvy3ej4fztwicmyr,

  output i1517rq45m7oy8,

  
  
  
  output c0z4i4kyokyx7sug, 
  input  w2kcsfod60d_68, 
  output [64-1:0] ntu21o6bz2w2777k4u,
  output ffyib96xpww6adq,   
  output owq8xep05y1_39287n92,
  output ya8t4ev_aidf0t0x4or,

  
  
  
  output                         v657dksgaz1cki9,
  output                         qzz1jhwf_vd0r8g, 
  input                          dwn42a1uvd9x3myec, 
  input                          p5fn_ooo9rctbxkgm_jui, 
  output [4 -1:0] uiojikf9vcnz,
  output [64 -1:0] x1_k6oouttg7m3f,
  output [64 -1:0] fcvvhg9v3mx,
  output [64 -1:0] l_v5xmhbzqc,
  output [3-1:0] i7iq7ecm_d9pi6uw6,
  input  a5z_23_ryr_m29hhia_p ,

  input  gf33atgy,
  input  ru_wi
  );


   
 assign ffyib96xpww6adq  = 1'b1;
 assign ntu21o6bz2w2777k4u = 64'b0;

 wire la5tvybv3d6kerf8nnu;

 assign x9a3z87q3adhgofd = 
          (w2kcsfod60d_68)  
        & (la5tvybv3d6kerf8nnu); 

 wire bc32c336qlwlrfbul8b = mt0f3958vekbx9 & w2kcsfod60d_68;
 assign c0z4i4kyokyx7sug   = mt0f3958vekbx9 & la5tvybv3d6kerf8nnu;



  
  assign qzz1jhwf_vd0r8g   = (~rnx27onf2lbe) & bc32c336qlwlrfbul8b;
  assign la5tvybv3d6kerf8nnu = rnx27onf2lbe ? 1'b1 : dwn42a1uvd9x3myec;
    
    
  assign i1517rq45m7oy8 = p5fn_ooo9rctbxkgm_jui & (~rnx27onf2lbe) ;

  wire yax5elqurk7q5708omh_o = 1'b0;

  assign uiojikf9vcnz  = lefkd05cxbpmfb;
  assign x1_k6oouttg7m3f  = wvg6yggd3_ngr;
  assign fcvvhg9v3mx  = fvamtne5n7;
  assign l_v5xmhbzqc  = w6fv3puuz49wu;

  assign i7iq7ecm_d9pi6uw6  = ahi4ptho3r9;

  wire aiavj0qzm_f22ey;
  assign v657dksgaz1cki9  = mt0f3958vekbx9 & x9a3z87q3adhgofd & (~aiavj0qzm_f22ey);

  assign owq8xep05y1_39287n92 = a5z_23_ryr_m29hhia_p;

  assign aiavj0qzm_f22ey = owq8xep05y1_39287n92 | yax5elqurk7q5708omh_o;

      
  assign ya8t4ev_aidf0t0x4or = 
                          
                      af5qc04tmn51e4u2h1z & 
                          
                      qzz1jhwf_vd0r8g & 
                          
                      tvy3ej4fztwicmyr;


endmodule                                      





















module moqpszi6cm8qllh02c2ny2 (
  input                            jfb7utzuy3zdlp,


  input                            z4423w2ovxgs284, 
  output                           s9k46re7yyb4d9, 



  input                            l_clnlob7ji8v9527, 
  input                            pnc251fe9pp3tm, 
  input                            h4sfadnxw7z3wz14, 

  input [4-1:0]     cpi07x9cy64pn2, 
  input [4-1:0]     eyd9fc4vjxutcl, 
  input [4-1:0]     pyhxgdg6s29imj, 



  input                            a_rhsk184ulq9ofyz,
  input                            ovpwjtytlapia4s3cl,
  input                            uo331eh1sm8wclmxid,
  input                            aseeilkazdwwcb4raoo2,
  input                            d67xmgrcefvmtl4jvxtz,
  input                            kgrl1ycpn2xb_uhommxp,
  input                            dj75s2vvoi93lk6c1i,
  input [4-1:0]     radwr7skyhm3jqso5,
  input [4-1:0]     zdid44qi3bv7q4phl,
  input [4-1:0]     lgrrvklyk4mm3aai,
  input [4-1:0]     ijxk119_taxeoqx0n,
  input [4-1:0]     brw5ihk9eaoddaefi7,
  input [4-1:0]     spknpgo66_t6t3dm__y,
  input [4-1:0]     ql612i235fqhavkhdu,
  input                            gawf4cwltls4ro8y_u,
  input [4-1:0]     przse28gs3o6cuvfp21u,

  input                            rz544x9yj6wtz, 
  input [4-1:0]     nkffqtpacz_8,
  input                            ipht6ss_sh6h,

  output                           qomzw_wq7v_mblz0qrfi,
  output                           r3d0cws3w3xmt0koa6l6g5,
  output                           k9fd4y9sg2l8f8pi29mz,
  output                           llha0lc4h8ie3t0l8,
  output                           t9le19upn_tsza2pzh3zii,
  output                           hv33acidoo0f1j4kpbs,
  output                           vpst0pbni2odvl7nr,
  output                           f015ahr7wg2fbe5_c5ja8,
  output                           yzu_ab6e_rylfgno7k0o2,
  output                           jcs6ikpya0beppu6gdyf,
  output                           g97p2rs03luvt0no8_ksk,
  output                           ip8580r8cp1_26jkauyh1wb,
  output                           j1otk5cqg9j9l3e8ynv,
  output                           dd92276i_tlq259bo27zu,
  output [5-1:0]   g_sda8atgrsb3n64a1e,
  output [5-1:0]   ih20zj50pzg1yxubdakxiz,
  output [5-1:0]   jenm8icl2nmc7a1huf5,
  output [5-1:0]   mosdlr9l78vgfsp3tj1,
  output [5-1:0]   x1k7b9da53adlb0frcz,
  output [5-1:0]   ky4jzzww3o0e66ldnngw1p,
  output [5-1:0]   zv9jo3fw_4ik299ra2irk87,
  output                           e5fsovqfl70bx4m4ahb3o,
  output                           nlb0f26rp9onx17ui5yzy,
  output [5-1:0]   irsej5jxvp566dv071e6,
  output                           do0utstzhn7g1d7unzt,
  output                           zjz6klk8496qrc03ps2snhs,
  output                           xkeclsgck5wllhwobaopvb0,
  output                           alnssn8w7d9iksq1ou7y2u,


  output                           hh0mpxxw3c00cet,
  output                           k1rpfwk8imnpek5,
  output [5-1:0]   kayddlyy2ps8dzeq46a,
  output                           t7m_v9aew2ud1e0u,


  input                            lr9ry0wds3k88rvde7n,
  input  [4-1:0]    smjqotzwkn9j4hf2ev_,



  input                          gy5zhpbrnl ,
  input                          qv70a7n8p ,
  input                          yrmykp4o9t ,
  input                          ojbpo5z6urt ,
  input                          cp7yy8bv2o8n, 
  input                          ypmn53drey,
  input                          msz_o10r_pkr,
  input                          q7qac2db3cbk ,
  input  [5-1:0] cpt0qfwiz,
  input  [5-1:0] vf7a_1kae4zv5,
  input  [5-1:0] rqj15_sdahil,
  input  [5-1:0] fhhe7189lmum ,






  output [4-1:0]     zzxn5x18ahgk4, 




  output                            i0fdxue89ury  ,
  output                            z4ufug6cvdodh  ,
  output                            vt96ugjl7qf4rqnj3  ,
  output [4-1:0]     kbmj0dq2hvlwx78s,
  output [4-1:0]     rod5c8pxpam5dt9n9y,
  output [4-1:0]     xu91lmfwk_nbjrz_,

  output                            zuht4f9qjrazipld4u    , 
  output                            g4qik0dwtex1gpiep    ,
  output                            f__fcmmb1thlj    ,

  output skcjh3xhs73ucsbh77  ,
  output s9kw_2m8ozw73_mbk1o0o   ,
  output sbtst18g6wurw5m36lm8 ,

  input  gf33atgy,
  input  ru_wi
);








  wire liv3kpxviwkwcfkc, nn5raw48sfe11a86eqf;
  wire g_5fx95j72v067js = z4423w2ovxgs284 & (~jfb7utzuy3zdlp);


  wire [5-1:0]      mm5sy6fi9qx1ad [12-1:0];
  wire [12-1:0] wqiilg_f9y1crs  ;
  wire [12-1:0] jsxiwlj_4lv9d4u3  ;
  wire [12-1:0] q4_f3wrbzd212 ;


  wire iqc4v0fr9otqnffpgcw9 = l_clnlob7ji8v9527;
  wire mdngcm0w7zytwnd1l6aeb = pnc251fe9pp3tm;
  wire q5fjhs31lnwsutg6p = h4sfadnxw7z3wz14;

  wire jlcr8smh9my82ie = z4423w2ovxgs284; 
  wire bus0pdx9it = iqc4v0fr9otqnffpgcw9 & nn5raw48sfe11a86eqf;
  wire g682g4pw8 = mdngcm0w7zytwnd1l6aeb & nn5raw48sfe11a86eqf;
  wire nm9ybeixu76e4 = q5fjhs31lnwsutg6p & nn5raw48sfe11a86eqf;

  wire l0kqs5qujoo = (g_5fx95j72v067js & liv3kpxviwkwcfkc); 
  wire f8fvunfazuj5_ = (iqc4v0fr9otqnffpgcw9 | mdngcm0w7zytwnd1l6aeb | q5fjhs31lnwsutg6p) & nn5raw48sfe11a86eqf;

  wire kssxyu60f27py = l0kqs5qujoo | f8fvunfazuj5_; 

  wire [12-1:0] p0pxcm18ooy8xh6qvhdtw1v [12-1:0];
  wire [12-1:0] xrrl9u13vmnr_173cfqjvpsb [12-1:0];




  wire [12-1:0] bkx7il15h  = xrrl9u13vmnr_173cfqjvpsb[cpi07x9cy64pn2];



  assign sbtst18g6wurw5m36lm8 = (~(|(bkx7il15h & jsxiwlj_4lv9d4u3)));




  wire [12-1:0] rxwng869s4mbek63ri, fngc_uksja8pbqk4ta1uirnvq, qbr9sihg2b56 ;
  wire [4-1:0] ockieugshbpn1o  [12-1:0]; 
  reg  [4-1:0] s62g1g; 
  wire [12-1:0] tgy4_citrvtconuxe ;

  wire [12-1:0] o6525a3aqckh_xovy, u9eroqp1_tki_5_e, cf0elxuu8_dcnkrsbo, bwg8wh_quk17o3qy40;
  wire [12-1:0] ghm38wwp2amo365 ;

  wire [12-1:0] f7clubvlsg56y3;
  wire [12-1:0] go2bdvq4k26eal5iy;
  wire [5-1:0]      g6jc55yn0k72o  [12-1:0]; 
  wire [12-1:0] xmej2zok7a811;


  assign fngc_uksja8pbqk4ta1uirnvq = {rxwng869s4mbek63ri[12-2:0],1'b0};


  wire [12-1:0] fh6h3pamni4h3zwy = ~jsxiwlj_4lv9d4u3 & ~tgy4_citrvtconuxe;
  genvar eoq;
  generate
    for (eoq = 0; eoq < 12; eoq = eoq+1) begin:fg2r376f5d2cmecff

      assign wqiilg_f9y1crs  [eoq] = f7clubvlsg56y3[eoq];
      assign jsxiwlj_4lv9d4u3 [eoq] = go2bdvq4k26eal5iy[eoq];
      assign mm5sy6fi9qx1ad[eoq] = g6jc55yn0k72o[eoq];
      assign q4_f3wrbzd212[eoq] = xmej2zok7a811[eoq];
      assign tgy4_citrvtconuxe[eoq] = lr9ry0wds3k88rvde7n & (smjqotzwkn9j4hf2ev_ == eoq[4-1:0]);


      assign rxwng869s4mbek63ri [eoq] = |fh6h3pamni4h3zwy[eoq:0]; 
      assign qbr9sihg2b56[eoq] = ({rxwng869s4mbek63ri[eoq],fngc_uksja8pbqk4ta1uirnvq[eoq]} == 2'b10) & l0kqs5qujoo;

      assign ghm38wwp2amo365 [eoq] = (l_clnlob7ji8v9527 & (cpi07x9cy64pn2 == eoq[4-1:0])) 
                               | (pnc251fe9pp3tm & (eyd9fc4vjxutcl == eoq[4-1:0])) 
                               | (h4sfadnxw7z3wz14 & (pyhxgdg6s29imj == eoq[4-1:0])) 
                               | (h4sfadnxw7z3wz14 & p0pxcm18ooy8xh6qvhdtw1v[pyhxgdg6s29imj][eoq]) 
                               ;

      assign o6525a3aqckh_xovy [eoq] = qbr9sihg2b56[eoq];
      assign u9eroqp1_tki_5_e [eoq] = go2bdvq4k26eal5iy[eoq] & ghm38wwp2amo365 [eoq]; 
      assign bwg8wh_quk17o3qy40 [eoq] = o6525a3aqckh_xovy [eoq] | u9eroqp1_tki_5_e [eoq]; 
      assign cf0elxuu8_dcnkrsbo [eoq] = o6525a3aqckh_xovy [eoq] ; 

      ux607_gnrl_dfflr #(1) ywcrpheyx3_dsfcvgbo4  (bwg8wh_quk17o3qy40 [eoq], cf0elxuu8_dcnkrsbo [eoq], go2bdvq4k26eal5iy[eoq], gf33atgy, ru_wi);


      ux607_gnrl_dfflr #(1                ) ktlux66gjbgb0pm_4th    (o6525a3aqckh_xovy [eoq], q7qac2db3cbk, f7clubvlsg56y3[eoq], gf33atgy, ru_wi);
      ux607_gnrl_dfflr #(1                ) c_1xy3c72gp25ox55pe    (o6525a3aqckh_xovy [eoq], ojbpo5z6urt, xmej2zok7a811[eoq], gf33atgy, ru_wi);
      ux607_gnrl_dfflr #(5) mi1jpp3frklv4iaqz    (o6525a3aqckh_xovy [eoq], fhhe7189lmum, g6jc55yn0k72o[eoq], gf33atgy, ru_wi);


      assign ockieugshbpn1o[eoq] = {4{qbr9sihg2b56[eoq]}} & eoq[4-1:0];

    end
  endgenerate

  integer qwj30yt;
  always @* begin: lrsp687zubjg1sb
    s62g1g=4'b0;

    for (qwj30yt = 0; qwj30yt < 12; qwj30yt = qwj30yt + 1) begin: gtxt_jgs23g66tlc
      s62g1g = s62g1g | (ockieugshbpn1o[qwj30yt]);

    end
  end
  assign zzxn5x18ahgk4 = s62g1g;
  assign skcjh3xhs73ucsbh77 = ~(|jsxiwlj_4lv9d4u3); 
  assign s9kw_2m8ozw73_mbk1o0o  = (&jsxiwlj_4lv9d4u3);
  assign liv3kpxviwkwcfkc = ~s9kw_2m8ozw73_mbk1o0o;
  assign nn5raw48sfe11a86eqf = ~skcjh3xhs73ucsbh77;

  assign s9k46re7yyb4d9 = ~(&(jsxiwlj_4lv9d4u3 | tgy4_citrvtconuxe)); 




  wire [4-1:0] zduqs6z3y59gw95y61[12-1:0];
  wire [4-1:0] a9bzkwa5l11zdhsid[12-1:0];
  wire [4-1:0] oo6jvtdsdx1i7k[12-1:0];
  wire [12-1:0] mv1xo_5em6tdfbey5, ywnps_v2dcmvt8m5i, egf66zgj9t_5;
  wire [12-1:0] vxioz_sstf9ilmrm, je0mdjs97sgnsb16qz, b5z1nh2r4a_4vypazh;
  wire [12-1:0] g2hb5wy7305zra, f49iz19fhxzbyfxlp, do_6ywq83oxjzjnc01;
  wire [12-1:0] od2labe2838d, nb3g7kcdyt7bwtvq, u4vwxxdwlql;
  wire [12-1:0] nl72agtv59k8jxctx, nr4t304uw_0bwlhie, rvu8dfiq2f7agq48_9f;
  reg [4-1:0] ofxcqyaipegys, jyp69_3c6ce00h7e, e8fbphi7t5pf39a9p;


  assign g2hb5wy7305zra = mv1xo_5em6tdfbey5 & vxioz_sstf9ilmrm;
  assign f49iz19fhxzbyfxlp = ywnps_v2dcmvt8m5i & je0mdjs97sgnsb16qz;
  assign do_6ywq83oxjzjnc01 = egf66zgj9t_5 & b5z1nh2r4a_4vypazh;
  assign nl72agtv59k8jxctx = od2labe2838d & g2hb5wy7305zra;
  assign nr4t304uw_0bwlhie = nb3g7kcdyt7bwtvq & f49iz19fhxzbyfxlp;
  assign rvu8dfiq2f7agq48_9f = u4vwxxdwlql & do_6ywq83oxjzjnc01;
  genvar wbrnq;
  generate
    for (wbrnq = 0; wbrnq < 12; wbrnq = wbrnq+1) begin:kx2bi7fhakvtge6b
      assign mv1xo_5em6tdfbey5[wbrnq] = ( ((cpt0qfwiz == mm5sy6fi9qx1ad[wbrnq]  ) & (q4_f3wrbzd212[wbrnq] & gy5zhpbrnl))
                                      ) & (!(wqiilg_f9y1crs[wbrnq] ^ cp7yy8bv2o8n)) & jsxiwlj_4lv9d4u3[wbrnq];
      assign ywnps_v2dcmvt8m5i[wbrnq] = ( ((vf7a_1kae4zv5 == mm5sy6fi9qx1ad[wbrnq]  ) & (q4_f3wrbzd212[wbrnq] & qv70a7n8p))
                                      ) & (!(wqiilg_f9y1crs[wbrnq] ^ ypmn53drey)) & jsxiwlj_4lv9d4u3[wbrnq];

      assign egf66zgj9t_5[wbrnq] = (rqj15_sdahil == mm5sy6fi9qx1ad[wbrnq]) & (q4_f3wrbzd212[wbrnq] & yrmykp4o9t) & (!(wqiilg_f9y1crs[wbrnq] ^ msz_o10r_pkr)) & jsxiwlj_4lv9d4u3[wbrnq];

      assign od2labe2838d [wbrnq] =  1'b0;
      assign nb3g7kcdyt7bwtvq [wbrnq] =  1'b0;
      assign u4vwxxdwlql [wbrnq] =  1'b0;


      assign vxioz_sstf9ilmrm [wbrnq] = ~(|(mv1xo_5em6tdfbey5 & (p0pxcm18ooy8xh6qvhdtw1v[wbrnq])));
      assign je0mdjs97sgnsb16qz [wbrnq] = ~(|(ywnps_v2dcmvt8m5i & (p0pxcm18ooy8xh6qvhdtw1v[wbrnq])));
      assign b5z1nh2r4a_4vypazh [wbrnq] = ~(|(egf66zgj9t_5 & (p0pxcm18ooy8xh6qvhdtw1v[wbrnq])));

      assign zduqs6z3y59gw95y61[wbrnq] = wbrnq[4-1:0] & {4{g2hb5wy7305zra[wbrnq]}} ;
      assign a9bzkwa5l11zdhsid[wbrnq] = wbrnq[4-1:0] & {4{f49iz19fhxzbyfxlp[wbrnq]}} ;
      assign oo6jvtdsdx1i7k[wbrnq] = wbrnq[4-1:0] & {4{do_6ywq83oxjzjnc01[wbrnq]}} ;

    end
  endgenerate

  integer vle3;
  always @* begin: wsczerl4_t
    ofxcqyaipegys =4'b0;
    jyp69_3c6ce00h7e =4'b0;
    e8fbphi7t5pf39a9p =4'b0;

    for (vle3 = 0; vle3 < 12; vle3 = vle3 + 1) begin: gtxt_jgs23g66tlc
      ofxcqyaipegys = ofxcqyaipegys | (zduqs6z3y59gw95y61[vle3]);
      jyp69_3c6ce00h7e = jyp69_3c6ce00h7e | (a9bzkwa5l11zdhsid[vle3]);
      e8fbphi7t5pf39a9p = e8fbphi7t5pf39a9p | (oo6jvtdsdx1i7k[vle3]);

    end
  end
  assign i0fdxue89ury   = |mv1xo_5em6tdfbey5;  
  assign z4ufug6cvdodh   = |ywnps_v2dcmvt8m5i;  
  assign vt96ugjl7qf4rqnj3   = |egf66zgj9t_5;  
  assign kbmj0dq2hvlwx78s = ofxcqyaipegys ; 
  assign rod5c8pxpam5dt9n9y = jyp69_3c6ce00h7e ; 
  assign xu91lmfwk_nbjrz_ = e8fbphi7t5pf39a9p ; 
  assign zuht4f9qjrazipld4u   = |nl72agtv59k8jxctx;  
  assign g4qik0dwtex1gpiep   = |nr4t304uw_0bwlhie;  
  assign f__fcmmb1thlj   = |rvu8dfiq2f7agq48_9f;  





  wire [12-1:0] wc7c8o96y4if0z[12-1:0];
  wire [12-1:0] iqfgc9z_el9q6hz8[12-1:0];
  wire [12-1:0] sumastwf7034[12-1:0];
  wire [12-1:0] sld2qsgbvj;
  wire sn83ikwu_h3kkcf,ocmg1tojp4vb,gukp8go0eh0,df2wahbunonfn,vu3mus3flydr,i67o2cy5f4zugi,rybjy8izve53rn,pizbltrm54mpt2r;
  wire [5-1:0] viptn9weuzus6poy    = mm5sy6fi9qx1ad[radwr7skyhm3jqso5];
  wire [5-1:0] kg23oj7fdhorkrfx    = mm5sy6fi9qx1ad[zdid44qi3bv7q4phl];
  wire [5-1:0] x_0tfxmh71jnn1kg    = mm5sy6fi9qx1ad[lgrrvklyk4mm3aai];
  wire [5-1:0] rzkr84024ft6vf    = mm5sy6fi9qx1ad[ijxk119_taxeoqx0n];
  wire [5-1:0] x6hnyaqye0kpk    = mm5sy6fi9qx1ad[brw5ihk9eaoddaefi7];
  wire [5-1:0] vpz0v76shajcj    = mm5sy6fi9qx1ad[spknpgo66_t6t3dm__y];
  wire [5-1:0] os4i213avqe2r    = mm5sy6fi9qx1ad[ql612i235fqhavkhdu];
  wire                         e11620qkl5r3wou    = q4_f3wrbzd212[radwr7skyhm3jqso5];
  wire                         x9ex8h_2i7f6yvw57    = q4_f3wrbzd212[zdid44qi3bv7q4phl];
  wire                         sl87f0dgmnav    = q4_f3wrbzd212[lgrrvklyk4mm3aai];
  wire                         yix6t6qzaoz7x9    = q4_f3wrbzd212[ijxk119_taxeoqx0n];
  wire                         h5l26ewme9wv15gs    = q4_f3wrbzd212[brw5ihk9eaoddaefi7];
  wire                         awew6umngjkye5q    = q4_f3wrbzd212[spknpgo66_t6t3dm__y];
  wire                         xerlkdd2n7s41    = q4_f3wrbzd212[ql612i235fqhavkhdu];

  wire [5-1:0] a9k4377giahx1vqnvx   = mm5sy6fi9qx1ad[nkffqtpacz_8     ];
  wire                         rqsvtowc6b3kjcb   = q4_f3wrbzd212[nkffqtpacz_8     ];
  wire                         wtsc7hwkdv9x3l3zq   = wqiilg_f9y1crs  [nkffqtpacz_8     ];
  wire [5-1:0] oxa30f1dcoe39    = mm5sy6fi9qx1ad[przse28gs3o6cuvfp21u];
  wire                         j6zegjwzp7jk1w8    = q4_f3wrbzd212[przse28gs3o6cuvfp21u];

  wire                         ffmrjo6p37h5kuzq4  = wqiilg_f9y1crs[lgrrvklyk4mm3aai];
  wire                         ps9w3vnj4poqw8md  = wqiilg_f9y1crs[brw5ihk9eaoddaefi7];
  wire                         nlq2ovp6x9pg  = wqiilg_f9y1crs[spknpgo66_t6t3dm__y];
  wire                         ikzxx6j5_176t  = wqiilg_f9y1crs[ql612i235fqhavkhdu];

  genvar siq,k4p2;
  generate
    for (k4p2 = 0; k4p2 < 12; k4p2 = k4p2+1) begin:u4q1p2sur234niw2w
      for (siq = 0; siq < 12; siq = siq+1) begin:g4r8u2e3llgggvg2v3uo

        if (k4p2 < siq) begin:p1ubj_kf6wfz7ho4um4qga

          assign iqfgc9z_el9q6hz8[k4p2][siq] = ( ((mm5sy6fi9qx1ad[k4p2] == mm5sy6fi9qx1ad[siq]) & (q4_f3wrbzd212[k4p2] & q4_f3wrbzd212[siq])) 
                                        )  & ((~wqiilg_f9y1crs[k4p2] & ~wqiilg_f9y1crs[siq])) & (jsxiwlj_4lv9d4u3[k4p2] & jsxiwlj_4lv9d4u3[siq]) ;

          assign sumastwf7034[k4p2][siq] = wqiilg_f9y1crs[k4p2] & wqiilg_f9y1crs[siq] & jsxiwlj_4lv9d4u3[k4p2] & jsxiwlj_4lv9d4u3[siq];
          assign wc7c8o96y4if0z[k4p2][siq] =  iqfgc9z_el9q6hz8[k4p2][siq] | sumastwf7034[k4p2][siq];
        end else if (k4p2 > siq) begin:dotuksoasi2kkgzk2qarh
          assign iqfgc9z_el9q6hz8[k4p2][siq] = 1'b0;
          assign sumastwf7034[k4p2][siq] = 1'b0;
          assign wc7c8o96y4if0z[k4p2][siq] = wc7c8o96y4if0z[siq][k4p2]; 
        end else begin:cwlesy7oyn4
          assign iqfgc9z_el9q6hz8[k4p2][siq] = 1'b0;
          assign sumastwf7034[k4p2][siq] = 1'b0;
          assign wc7c8o96y4if0z[k4p2][siq] = 1'b0; 
        end 
      end
      assign sld2qsgbvj[k4p2] = |(wc7c8o96y4if0z[k4p2] & xrrl9u13vmnr_173cfqjvpsb[k4p2]);
    end
  endgenerate

  assign sn83ikwu_h3kkcf  = |(sld2qsgbvj[radwr7skyhm3jqso5]);
  assign ocmg1tojp4vb  = |(sld2qsgbvj[zdid44qi3bv7q4phl]);
  assign gukp8go0eh0  = |(sld2qsgbvj[lgrrvklyk4mm3aai]);
  assign df2wahbunonfn  = |(sld2qsgbvj[ijxk119_taxeoqx0n]);
  assign vu3mus3flydr  = |(sld2qsgbvj[brw5ihk9eaoddaefi7]);
  assign i67o2cy5f4zugi  = |(sld2qsgbvj[spknpgo66_t6t3dm__y]);
  assign rybjy8izve53rn  = |(sld2qsgbvj[ql612i235fqhavkhdu]);
  wire   yqym8e314ri5a5_  = |(sld2qsgbvj[przse28gs3o6cuvfp21u]);
  assign pizbltrm54mpt2r = |(sld2qsgbvj[nkffqtpacz_8     ]);


  assign qomzw_wq7v_mblz0qrfi = ~sn83ikwu_h3kkcf  ;
  assign r3d0cws3w3xmt0koa6l6g5 = ~ocmg1tojp4vb  ;
  assign k9fd4y9sg2l8f8pi29mz = ~gukp8go0eh0  ;
  assign llha0lc4h8ie3t0l8 = ~df2wahbunonfn  ;
  assign t9le19upn_tsza2pzh3zii = ~vu3mus3flydr  ;
  assign hv33acidoo0f1j4kpbs = ~i67o2cy5f4zugi  ;
  assign vpst0pbni2odvl7nr = ~rybjy8izve53rn  ;

  assign f015ahr7wg2fbe5_c5ja8 = e11620qkl5r3wou ;
  assign yzu_ab6e_rylfgno7k0o2 = x9ex8h_2i7f6yvw57 ;
  assign jcs6ikpya0beppu6gdyf = sl87f0dgmnav ;
  assign g97p2rs03luvt0no8_ksk = yix6t6qzaoz7x9 ;
  assign ip8580r8cp1_26jkauyh1wb = h5l26ewme9wv15gs ;
  assign j1otk5cqg9j9l3e8ynv = awew6umngjkye5q ;
  assign dd92276i_tlq259bo27zu = xerlkdd2n7s41 ;

  assign e5fsovqfl70bx4m4ahb3o   = ~yqym8e314ri5a5_  ;
  assign nlb0f26rp9onx17ui5yzy = j6zegjwzp7jk1w8 ;
  assign irsej5jxvp566dv071e6 = oxa30f1dcoe39 ;



  assign g_sda8atgrsb3n64a1e = viptn9weuzus6poy ;
  assign ih20zj50pzg1yxubdakxiz = kg23oj7fdhorkrfx ;
  assign jenm8icl2nmc7a1huf5 = x_0tfxmh71jnn1kg ;
  assign mosdlr9l78vgfsp3tj1 = rzkr84024ft6vf ;
  assign x1k7b9da53adlb0frcz = x6hnyaqye0kpk ;
  assign ky4jzzww3o0e66ldnngw1p = vpz0v76shajcj ;
  assign zv9jo3fw_4ik299ra2irk87 = os4i213avqe2r ;



  assign hh0mpxxw3c00cet        = ~pizbltrm54mpt2r ;
  assign k1rpfwk8imnpek5      = rqsvtowc6b3kjcb;
  assign kayddlyy2ps8dzeq46a      = a9k4377giahx1vqnvx;
  assign t7m_v9aew2ud1e0u      = wtsc7hwkdv9x3l3zq;

  assign do0utstzhn7g1d7unzt = ffmrjo6p37h5kuzq4 ;
  assign zjz6klk8496qrc03ps2snhs = ps9w3vnj4poqw8md ;
  assign xkeclsgck5wllhwobaopvb0 = nlq2ovp6x9pg ;
  assign alnssn8w7d9iksq1ou7y2u = ikzxx6j5_176t ;



  wire [12*12-1:0]  egekc6m62wqwt_hqe7nfhk;
  p_nv4xk50a2bh9h4mr5fv #(.o10eaknnnv(12))
     cvaxldgq7wiycs4xz2tjupu9 (
      .h1zifc6wetrm6wm (qbr9sihg2b56),
      .oybz4sq2nhg8_26o(egekc6m62wqwt_hqe7nfhk),

      .gf33atgy  (gf33atgy  ),
      .ru_wi(ru_wi)

  );
  genvar gmw1b,jgaeu52;
  generate
    for (gmw1b = 0; gmw1b < 12; gmw1b = gmw1b+1) begin:lhk_iy
      for (jgaeu52 = 0; jgaeu52 < 12; jgaeu52 = jgaeu52+1) begin:dfswcsxay



        if (gmw1b < jgaeu52) begin:fstpedp5s67a0fp 
          assign p0pxcm18ooy8xh6qvhdtw1v[gmw1b][jgaeu52] = ~egekc6m62wqwt_hqe7nfhk[gmw1b*12+jgaeu52];
        end
        else begin :a7o0gf5dl9wm9_t2
          assign p0pxcm18ooy8xh6qvhdtw1v[gmw1b][jgaeu52] = egekc6m62wqwt_hqe7nfhk[jgaeu52*12+gmw1b];

        end
        if (gmw1b <= jgaeu52) begin:a854ydgl64zv 
          assign xrrl9u13vmnr_173cfqjvpsb[gmw1b][jgaeu52] = egekc6m62wqwt_hqe7nfhk[gmw1b*12+jgaeu52];
        end
        else begin:ada_5kch5qcf9kcn7 
          assign xrrl9u13vmnr_173cfqjvpsb[gmw1b][jgaeu52] = ~egekc6m62wqwt_hqe7nfhk[jgaeu52*12+gmw1b];
        end
      end
    end
  endgenerate 

endmodule





















module uh_y21ipql6al1c4qkqfokr_0yd(



  input                          r25vjm_g303hv5mr__oydfc50s_6, 
  output                         q3nebxbyx8x_n2wgt90jxx5ppnlbuzt, 
  input  [64-1:0]        l9uyi_93i_vkb6davalokxbus3edyu ,
  input  [4 -1:0] kptoalwjf0vnjxpubirzzg8r1l0_hk7 ,
  input                          qd2ehv6u5ipjg2sd3swjn38uuab  , 

  input                          x0wwmbj55rz1_gzemtenuutvu4f5gtbr, 
  output                         tjf2j_x0_19wvbnushzloo4vpibe0q, 
  input  [64-1:0]        jcur3i2c0we7b6x5ms3vw9himw35v ,
  input  [4 -1:0] vmujqgbzxn6hqc5j49ufmtewa7 ,
  input                          x74i2xb96e9fui_1revcqt088tm0hf  , 


  input                          wqlni2o6ysdnyxmiesc2c9nx1nhsidr, 
  output                         bx1s0daa65s6eao0yo05dgpi6o_6e7, 
  input  [64-1:0]        cefmw490fob0947fn0zxl51_fkeb ,
  input  [4 -1:0] csw73tw17ceolm9eifmbhd887zfa ,
  input                          fu2trk07aq8pgduthe_h3zskathrh  , 
  input  [4:0]                   p5laf3iz7k000k42fpww1tjw97c514pj,

  input                          kq64hafe_jmlm63rt4w15_qnftr01,
  input                          en8f11yeo7j9u54v7agnvuncx9kha,
  input                          pqeyh89bzfwni86npwrcnmz1fjtb2dhfj,
  input                          os5_rc90_7gawcz0efrilvhb5wo74r9,
  input [64 -1:0]   zllz_u37t659z507dtl4d906nsg35,
  input [64 -1:0]     i5m1rrdydixypqcxzmalcomh  ,
  input                          laifryt4bl834uov7isyxe_4uk3_d  ,
  input                          yvw2qnvbiajkt2mcxp4j4xqiucb8  ,





  input                          obli6e3v4_8bjrltqdv6v18stt0fev4 , 
  output                         tb6a57t86vwitea0x8780ksclx8d4 , 
  input  [64-1:0]        jomr8wem988b32tidmg2zkgiqgl6  ,
  input  [4 -1:0] boxfq4ncnb8czlmq7p4msay3wg7o4  ,
  input                          k98w6098j0wekfd9wjqjkmtslxo   , 
  input  [4:0]                   jz83wrre56m2b7vf1dnwnnu8lme , 
  input                          vo9o42ohfekmv2b390b9ovdxs7hswv , 
  output                         xvr_92a8rcvf2quyrmigj7fzuftq , 
  input  [64-1:0]        yhqkr966fkfranbq6mys4_itfdsz8  ,
  input  [4 -1:0] ktpgkhezvy18ox4t8b5xhresqcnvqp6  ,
  input                          jqaxpjo0j1mrf8casph8bqvmhaf   , 
  input  [4:0]                   d4xh57em8iunsz9w5_jruofpuezsh , 
  input                          z0p5c0vl91tsjk1lmt8kxat0kig3dlom , 
  output                         kqhgic2ez1gu2b308vr7gayeops , 
  input  [64-1:0]        or2q_8b_zdv2o7h7ol6rtfs9p7sqzx9  ,
  input  [4 -1:0] zo0u9kjy8fmzeh_qnut3gcckfj_  ,
  input                          emdo9xkvazh0e830c3tezq85cr   , 
  input  [4:0]                   c90btjrwqlw7w7j9o1twzgjt43njm3wg , 
  input                          wqn_diiyx7s7t037qfg_nkqdnix, 
  output                         aeqpr5hrp251jp0yxm1vcqjoftohs, 
  input  [64-1:0]        vqzbvg_jyxunlaurqlpwhp34u_jx0 ,
  input  [4 -1:0] t1tkrihuzsa8iq9pywbo4a3ktie7wn4 ,
  input                          ytkv6_mmnisydnwtk48igroblctc  , 



  output                          gqat5ctwgmxi8n_5z03tivvpgqx6j5kb, 
  input                           n0cmggtax9qzrd4qsy1cdbik144lmx, 
  output  [64-1:0]        y4aoa0ok7ylngx_33gfqr0g1md0g8dj ,
  output  [4 -1:0] zmotzlbzlmuf2isjtqn2h8beel09 ,
  output                          vo2fj15n058l2wpxbodnsdqxwkdn08  , 

  output                          vi7663z7hxlc4ngkh1_yfoxfpvbiq, 
  input                           rhwm1lw0wyhvdhss4f3p_v5zkroo, 
  output  [64-1:0]        vsgctu8mzjw91ryb865p9r7s8fp ,
  output  [4 -1:0] ql2r_7apgocbap5k7ucf5a673x7v ,
  output                          sei0me3z77b60zu8tfykejc6_w  , 


  output                          bm0yhprev2rfpkaztktaxtnq7f8q0bp, 
  input                           f_7j356ybgmsh86n3umtlmih2ee8c5, 
  output  [64-1:0]        ktwrzuv2gg846pksncc26g4y0pe1h,
  output  [4 -1:0] i2kgxrwehfoyscnln10tc70_omph,
  output                          xp4xfk612_1jfargldlbq2rjb , 
  output  [4:0]                   lrojclgmk96728ugf1xss07x7gzfgls,

  output                           rdsej_3e3o2bh3ld92ygwf707k988,
  output                           eitel8xkigdj96m3f89nsi2w_71pvf,
  output                           eovnqir46kp7wnkzr0btiuicjboull,
  output                           qc6yp7yoe_bjq2am96mg0sizkq7os,
  output [64 -1:0]    lo4an3qbdgmg6hqsqosvvk8dwctnn1wy6c,
  output [64 -1:0]      xedi2t9w7jc8_rstzke961dl4l7  ,
  output                           az7mzc_81tib2dpb5d3a70_wdp73f  ,
  output                           oopk92ymqbivd2dxs85nt1ly5ccn  ,




  output                          gkb40bm903wc32_2zjmb0l25g21p7 , 
  input                           j0l8i3eed1ek492qjzm9uejf41sz , 
  output [64-1:0]         yyasjan35_68l3cq8a3ioaew9bbhr  ,
  output [4 -1:0]  yu_1foait_ukyv14b73xepo_1mj31mu  ,
  output                          pdkr3e96qk7jfuv5c8967qald7p   , 
  output  [4:0]                   xfz4lyb4bxla1gb3kuqf0gcek1_r8yz , 
  output                          scom2gns1t5jrniqayb84g_h2a1zaxbv , 
  input                           jzh4duikrv004mprz7zksk2dh9ty72 , 
  output [64-1:0]         geun5etyjtjsnydbal2egw52gf34  ,
  output [4 -1:0]  xpvibysxiip4tytx5_ry26i78ce4j4  ,
  output                          kng9rvszc8o8ob5v1_ak0ipg9lgbku   , 
  output  [4:0]                   avrbak7i2ou0is2fulrxcpx4b8qjfwus , 
  output                          ky7mnv5l4jl0v17ox278fwktul3qti , 
  input                           wt906274r_7subjpzosffvtc_8lbfu , 
  output [64-1:0]         fsr9hzh57oj6r29w8_fdfss2962  ,
  output [4 -1:0]  a9_1a439ejmx35qe2g8yihj84g5  ,
  output                          n412jv5dj1tvgdf8jls7u2bjvh   , 
  output  [4:0]                   ke2zqim9rdwj_bmursxrbh8ga08qo , 
  output                          rhx_hd60cwxftbqnr_uhlcmbab17eeue, 
  input                           gm94l7jeucs5_57r7b1ghqbrvubvg, 
  output  [64-1:0]        wtj2dgdc6vyaj4ptn464rhnsgz1 ,
  output  [4 -1:0] l_w88r7i0zq6u0xtcywbwzu__s ,
  output                          om2j1tmzbckjwmzuoudwijwh6gh_ig  , 


  input  gf33atgy,
  input  ru_wi
  );



  localparam aafrtcd422sh = 64 + 4 + 1;
  localparam jdklkkziw = 64 + 4 + 1;
  localparam ng5xxjooywsar = 64 
                       + 4 
                       + 1 
                       + 5
                       + 1 
                       + 1 
                       + 64 
                       + 64 
                       + 1  
                       + 1  
                       ; 
  localparam x7rgtpkxfa2t = 64 + 4 + 1+5;
  localparam tg_f7qr4nitb = 64 + 4 + 1+5;
  localparam p3emkgj9cw3k = 64 + 4 + 1+5;
  localparam srzgl2bpw5p0 = 64 
                       + 4 
                       + 1 
                       ;


  wire [aafrtcd422sh-1:0] hb34z7utpsm4t6sckxq0uxkb7o9dn = {
                                          l9uyi_93i_vkb6davalokxbus3edyu,
                                          kptoalwjf0vnjxpubirzzg8r1l0_hk7,   
                                          qd2ehv6u5ipjg2sd3swjn38uuab
                                        };   
  wire [aafrtcd422sh-1:0] dtw_j2_uf00leoaryr6b9g0a5b; 
  ux607_gnrl_bypbuf # (
    .DP(1),
    .DW(aafrtcd422sh) 
  ) e4xtcpqqz2ghklwcaerhx(
      .i_vld   (r25vjm_g303hv5mr__oydfc50s_6),
      .i_rdy   (q3nebxbyx8x_n2wgt90jxx5ppnlbuzt),

      .o_vld   (gqat5ctwgmxi8n_5z03tivvpgqx6j5kb),
      .o_rdy   (n0cmggtax9qzrd4qsy1cdbik144lmx),

      .i_dat   (hb34z7utpsm4t6sckxq0uxkb7o9dn),
      .o_dat   (dtw_j2_uf00leoaryr6b9g0a5b),

      .clk     (gf33atgy  ),
      .rst_n   (ru_wi)
  );
  assign { y4aoa0ok7ylngx_33gfqr0g1md0g8dj,
           zmotzlbzlmuf2isjtqn2h8beel09,   
           vo2fj15n058l2wpxbodnsdqxwkdn08
         } = dtw_j2_uf00leoaryr6b9g0a5b;



  wire [jdklkkziw-1:0] boakmkz1yknw7bmmvfhxb22gtu1 = {
                                          jcur3i2c0we7b6x5ms3vw9himw35v,
                                          vmujqgbzxn6hqc5j49ufmtewa7,   
                                          x74i2xb96e9fui_1revcqt088tm0hf
                                        };   
  wire [jdklkkziw-1:0] ezo7zt9b0s8ikxclqpvflwpusg; 
  ux607_gnrl_bypbuf # (
    .DP(1),
    .DW(jdklkkziw) 
  ) b3edcpig75a5bhzpn2f1hxa_g(
      .i_vld   (x0wwmbj55rz1_gzemtenuutvu4f5gtbr),
      .i_rdy   (tjf2j_x0_19wvbnushzloo4vpibe0q),

      .o_vld   (vi7663z7hxlc4ngkh1_yfoxfpvbiq),
      .o_rdy   (rhwm1lw0wyhvdhss4f3p_v5zkroo),

      .i_dat   (boakmkz1yknw7bmmvfhxb22gtu1),
      .o_dat   (ezo7zt9b0s8ikxclqpvflwpusg),

      .clk     (gf33atgy  ),
      .rst_n   (ru_wi)
  );
  assign { vsgctu8mzjw91ryb865p9r7s8fp,
           ql2r_7apgocbap5k7ucf5a673x7v,   
           sei0me3z77b60zu8tfykejc6_w
         } = ezo7zt9b0s8ikxclqpvflwpusg;



  wire [ng5xxjooywsar-1:0] v0unl2jq4xn1a6e7hn5g2loh3cc = {
                                 cefmw490fob0947fn0zxl51_fkeb,
                                 csw73tw17ceolm9eifmbhd887zfa,   
                                 fu2trk07aq8pgduthe_h3zskathrh,
                                 p5laf3iz7k000k42fpww1tjw97c514pj,

                                 kq64hafe_jmlm63rt4w15_qnftr01,
                                 en8f11yeo7j9u54v7agnvuncx9kha,
                                 zllz_u37t659z507dtl4d906nsg35,
                                 i5m1rrdydixypqcxzmalcomh  ,
                                 laifryt4bl834uov7isyxe_4uk3_d  ,
                                 yvw2qnvbiajkt2mcxp4j4xqiucb8   
                                        };   
  wire [ng5xxjooywsar-1:0] zbjsb7att7lfx3drs9t_zcph9r1ns02; 
  ux607_gnrl_bypbuf # (
    .DP(1),
    .DW(ng5xxjooywsar) 
  ) lm9v8zkuahz5wc66rhyt2(
      .i_vld   (wqlni2o6ysdnyxmiesc2c9nx1nhsidr),
      .i_rdy   (bx1s0daa65s6eao0yo05dgpi6o_6e7),

      .o_vld   (bm0yhprev2rfpkaztktaxtnq7f8q0bp),
      .o_rdy   (f_7j356ybgmsh86n3umtlmih2ee8c5),

      .i_dat   (v0unl2jq4xn1a6e7hn5g2loh3cc),
      .o_dat   (zbjsb7att7lfx3drs9t_zcph9r1ns02),

      .clk     (gf33atgy  ),
      .rst_n   (ru_wi)
  );
  assign { ktwrzuv2gg846pksncc26g4y0pe1h,
           i2kgxrwehfoyscnln10tc70_omph,   
           xp4xfk612_1jfargldlbq2rjb,
           lrojclgmk96728ugf1xss07x7gzfgls,
           rdsej_3e3o2bh3ld92ygwf707k988,
           eitel8xkigdj96m3f89nsi2w_71pvf,
           lo4an3qbdgmg6hqsqosvvk8dwctnn1wy6c,
           xedi2t9w7jc8_rstzke961dl4l7  ,
           az7mzc_81tib2dpb5d3a70_wdp73f  ,
           oopk92ymqbivd2dxs85nt1ly5ccn   

         } = zbjsb7att7lfx3drs9t_zcph9r1ns02;

assign  eovnqir46kp7wnkzr0btiuicjboull = 1'b0;
assign  qc6yp7yoe_bjq2am96mg0sizkq7os = 1'b0;








  wire [x7rgtpkxfa2t-1:0] oodnj3adhupvq1jpog_yxwp45j = {
                                          jomr8wem988b32tidmg2zkgiqgl6,
                                          boxfq4ncnb8czlmq7p4msay3wg7o4,   
                                          k98w6098j0wekfd9wjqjkmtslxo ,
                                          jz83wrre56m2b7vf1dnwnnu8lme   
                                        };   
  wire [x7rgtpkxfa2t-1:0] vdmdz2ogqpfn53rs6bdik1haf4kj857; 
  ux607_gnrl_bypbuf # (
    .DP(1),
    .DW(x7rgtpkxfa2t) 
  ) gi02bel2tob4p7ejgxjt(
      .i_vld   (obli6e3v4_8bjrltqdv6v18stt0fev4),
      .i_rdy   (tb6a57t86vwitea0x8780ksclx8d4),

      .o_vld   (gkb40bm903wc32_2zjmb0l25g21p7),
      .o_rdy   (j0l8i3eed1ek492qjzm9uejf41sz),

      .i_dat   (oodnj3adhupvq1jpog_yxwp45j),
      .o_dat   (vdmdz2ogqpfn53rs6bdik1haf4kj857),
  
      .clk     (gf33atgy  ),
      .rst_n   (ru_wi)
  );
  assign { yyasjan35_68l3cq8a3ioaew9bbhr,
           yu_1foait_ukyv14b73xepo_1mj31mu,   
           pdkr3e96qk7jfuv5c8967qald7p,
           xfz4lyb4bxla1gb3kuqf0gcek1_r8yz   
         } = vdmdz2ogqpfn53rs6bdik1haf4kj857;



  
  wire [tg_f7qr4nitb-1:0] hzlbzw3p7enjdx8zwc1s8fmgzr = {
                                          yhqkr966fkfranbq6mys4_itfdsz8,
                                          ktpgkhezvy18ox4t8b5xhresqcnvqp6,   
                                          jqaxpjo0j1mrf8casph8bqvmhaf,
                                          d4xh57em8iunsz9w5_jruofpuezsh   
                                        };   
  wire [tg_f7qr4nitb-1:0] qmjwor1dm2mnp2c5ec79mulcijdn; 
  ux607_gnrl_bypbuf # (
    .DP(1),
    .DW(tg_f7qr4nitb) 
  ) pfktstdzqxenrcpy2j2z8y2(
      .i_vld   (vo9o42ohfekmv2b390b9ovdxs7hswv),
      .i_rdy   (xvr_92a8rcvf2quyrmigj7fzuftq),

      .o_vld   (scom2gns1t5jrniqayb84g_h2a1zaxbv),
      .o_rdy   (jzh4duikrv004mprz7zksk2dh9ty72),

      .i_dat   (hzlbzw3p7enjdx8zwc1s8fmgzr),
      .o_dat   (qmjwor1dm2mnp2c5ec79mulcijdn),
  
      .clk     (gf33atgy  ),
      .rst_n   (ru_wi)
  );
  assign { geun5etyjtjsnydbal2egw52gf34,
           xpvibysxiip4tytx5_ry26i78ce4j4,   
           kng9rvszc8o8ob5v1_ak0ipg9lgbku,
           avrbak7i2ou0is2fulrxcpx4b8qjfwus   
         } = qmjwor1dm2mnp2c5ec79mulcijdn;


  
  wire [p3emkgj9cw3k-1:0] kjhdhrc8ggehzmh0wb4f5p81kix = {
                                          or2q_8b_zdv2o7h7ol6rtfs9p7sqzx9,
                                          zo0u9kjy8fmzeh_qnut3gcckfj_,   
                                          emdo9xkvazh0e830c3tezq85cr,
                                          c90btjrwqlw7w7j9o1twzgjt43njm3wg   
                                        };   
  wire [p3emkgj9cw3k-1:0] wbyta_rfxghemhgn5ozdn_glswiqvyu; 
  ux607_gnrl_bypbuf # (
    .DP(1),
    .DW(p3emkgj9cw3k) 
  ) h_dcqamkig9o7t27qj0e4u(
      .i_vld   (z0p5c0vl91tsjk1lmt8kxat0kig3dlom),
      .i_rdy   (kqhgic2ez1gu2b308vr7gayeops),

      .o_vld   (ky7mnv5l4jl0v17ox278fwktul3qti),
      .o_rdy   (wt906274r_7subjpzosffvtc_8lbfu),

      .i_dat   (kjhdhrc8ggehzmh0wb4f5p81kix),
      .o_dat   (wbyta_rfxghemhgn5ozdn_glswiqvyu),
  
      .clk     (gf33atgy  ),
      .rst_n   (ru_wi)
  );
  assign { fsr9hzh57oj6r29w8_fdfss2962,
           a9_1a439ejmx35qe2g8yihj84g5,   
           n412jv5dj1tvgdf8jls7u2bjvh,
           ke2zqim9rdwj_bmursxrbh8ga08qo   
         } = wbyta_rfxghemhgn5ozdn_glswiqvyu;






  wire [srzgl2bpw5p0-1:0] ildka6xii77uow6ottci71ayi997 = {
                                          vqzbvg_jyxunlaurqlpwhp34u_jx0,
                                          t1tkrihuzsa8iq9pywbo4a3ktie7wn4,   
                                          ytkv6_mmnisydnwtk48igroblctc 
                                        };   
  wire [srzgl2bpw5p0-1:0] nzik7bn1maqa35sfrrhvebxfpmqqp; 
  ux607_gnrl_pipe_stage # (
    .DP(2),
    .DW(srzgl2bpw5p0) 
  ) yufitvgtioha0e0m6fccedge(
      .i_vld   (wqn_diiyx7s7t037qfg_nkqdnix),
      .i_rdy   (aeqpr5hrp251jp0yxm1vcqjoftohs),

      .o_vld   (rhx_hd60cwxftbqnr_uhlcmbab17eeue),
      .o_rdy   (gm94l7jeucs5_57r7b1ghqbrvubvg),

      .i_dat   (ildka6xii77uow6ottci71ayi997),
      .o_dat   (nzik7bn1maqa35sfrrhvebxfpmqqp),
  
      .clk     (gf33atgy  ),
      .rst_n   (ru_wi)
  );
  assign { wtj2dgdc6vyaj4ptn464rhnsgz1,
           l_w88r7i0zq6u0xtcywbwzu__s,   
           om2j1tmzbckjwmzuoudwijwh6gh_ig
         } = nzik7bn1maqa35sfrrhvebxfpmqqp;



endmodule                                      


























module uv355zczoyyqi_qujlvi(



  input                         y40x_uwnqs6f   ,
  input                         qlykdb48c89hfbq5l3v ,
  input [5-1:0] ejlcmcywa2ghgwvj ,
  input                         fk7qm80i_py_6   ,
  input                         utfce4yxn08kh9t ,
  input [5-1:0] gof9x1lyu2n5rnf ,
  input                         f7t_bak0dfaq3   ,
  input                         oy1tzeyrsbr3bg7dr9u ,
  input                         rpnvo9xxx6nke515 , 
  input [5-1:0] v2fkznl9m7dtfymx ,
  input                         tdg7ccg5dltr5l9s, 
  input                         z5s1cielsyyeza34h, 
  input [5-1:0] ggpqgd6b8zuelz8, 


  input                           ll0_hbknv5bc_8mxvx5c,
  output                          qloskxsiztazdeq2ad95i,
  input [64-1:0]          px17v86p_7_1fdvm1w,
  input  [4-1:0]   jb9locwfccqzb06jjon,
  input                           a3g162j6o30b4qdpd_z,

  input                          q89zlvtwzxkjd6h5k, 
  input                          gjoru9khthrg8j6pfamu, 
  input                          vf6etunsloifr12azv4he6, 
  input [5-1:0]  f63hhh0gzajzsiyjd8cqb,
  input                          v7f1q1_fp5fc8b_u, 
  input                          mvneatl67xbzspkpyi1, 
  input                          ltzlg4gy4noc9555li, 
  input [5-1:0]  nfozodmnsmlv22fi3oe,
  input                          vmwegtj2c0zt7rilpw, 
  input                          szgl0r6i254qax8jkjr, 
  input                          bp90ffmjkj3u4__poo, 
  input [5-1:0]  nq8gzr65b3p_cdc52lshh,

  input                          ju3gksnn2mup5h81eh28, 
  output                         tymuflph4h7mej5umh86, 
  input  [64-1:0]        c5csn3nczo8zlvq621sy,
  input  [5-1:0]                 rd0rvbiicactt4sbf,
  input  [4 -1:0] g5gmidj6od8k58avl_h9y,
  input                          h5w2di84ketcahr4 , 

  input                          lanyt81iat_ws21fv, 
  output                         b1eabu9fa3jnjln5tc, 
  input  [64-1:0]        nt0ndhbk6x29ae8da95,
  input  [5-1:0]                 ri8f9g_paihffhz9_8qgu,
  input  [4 -1:0] u7vn3gjmd4owzsi7tk,
  input                          ik4ulvmx89l0u0ko ,

  input                          nz5iij5cadsnx4fokudqbo,
  output                         bz1hc72g_22hgoqs8,
  input  [64-1:0]        wctv6a1mmq6dtwsg9n,
  input  [5-1:0]                 onijw658b2__et8fr1has,
  input  [4 -1:0] zakjetcb_4mzmn_bchz,
  input                          ys8dsx5hx_injk9b ,





  input                         ipq0f4_yvmml7o06891, 
  output                        p4jgl36nmqe8ud7_g4i7, 
  input  [64-1:0]       wyhg5n7dklr59dxgm_bs,
  input                         cbr_upfu_0ywren54f,
  input  [4-1:0] ubk6j4rwgfrf5ryn1ibp,


  
  
  input  o9vvv_q4ikz_2yp0w, 
  output c1ilkc2r6es72c5h2vcc, 
  input  [64-1:0] l3sefagtx4ai4ljb,
  input  bjn5x3u7v4u3rm6d,
  input  [4-1:0] josyt39cvr3gignopao,



  input                          vacmjbyuw8jriztdg, 
  output                         dlogavn_28q56zummtut, 
  input  [64-1:0]        yhfc75p_gcdigu,
  input  [4 -1:0] zl0t249z3fcwyj4puu,
  input                          psylshnv8k3qqz5i , 
  input                          p_2daj_9kqsf0ekr101 ,
  input                          djb42mrmnunfufgxzh ,
  input  [64 -1:0]  vqldrx_4vk7av570m8fv,
  input  [64 -1:0]    zhwwio_mprrvjud04,
  input                          pxbhqh6yl6hotx, 
  input                          toib7p7z_deij2b, 
  input  [4:0]                   wk41j07s3anl9_t, 
  input                          p7ah58va5_2njbtv,
  input [64-1:0]         u981qrwkgi5h0e72b__gg19w,
  input                          p0i2i3v3j1tclelx51,



  output p1jdw9loxkz60taq_vkp_3, 
  input  ar7xgugq1a_pz7b82ds, 
  output [64-1:0] jwwku_el5h5h2lx6e0kyi,
  output [5-1:0] zt19omidnr_zyp2gc3bywfb,
  output [5 -1:0] vjhpkmep8g_u_cizhsw,
  output [4-1:0] eo5skx1ygvzuasbjgnyl,
  output v19st7vd9_bi485e6ak0,
  output gccap1c6hft7o1z7esm,




  output  z2qyay491938ppnlxuc,
  input   pbtolkl953sk14id0iy,
  output  zeseql2htbxpugyu5_j,
  output  al3t866kz4po45vfuyjy,
  output  xutsaulafh4onxtthm8n , 
  output  me7unt7fapqqhtc6epso , 
  output [64-1:0] m2as3qe7miuhj662j1zvt,







  output xd2ftroj1i79g4derw,
  output [4 -1:0] qoxd9f57dl083f6cm, 


  input  gf33atgy,
  input  ru_wi
  );

  wire mxa77etukhs8o_5z6962l19;
  wire vtv633e4nu9j19d_x9dbyga8du = (mxa77etukhs8o_5z6962l19 & (~z2qyay491938ppnlxuc)) 
                                  | p7ah58va5_2njbtv
                                  ; 

  localparam jwxxo5dwz741q1 = 64+4+1
                           ; 
  wire [jwxxo5dwz741q1-1:0] srufsypxvg1hqxwmw0y;
  wire [jwxxo5dwz741q1-1:0] yhopxd2wrapvsuiglom;


  ux607_gnrl_pipe_stage #(
  .CUT_READY(0),
  .DP(1),
  .DW(jwxxo5dwz741q1)
  ) ow_caaylzt9o9k0lbs(
    .i_vld      (vtv633e4nu9j19d_x9dbyga8du),
    .i_rdy      (),
    .i_dat      (srufsypxvg1hqxwmw0y),

    .o_vld      (z2qyay491938ppnlxuc),
    .o_rdy      (pbtolkl953sk14id0iy),
    .o_dat      (yhopxd2wrapvsuiglom),

    .clk        (gf33atgy),
    .rst_n      (ru_wi)
  );














  wire tj9rezp6j0u0mvddq;
  wire zl3w_sym4l3ca;

  wire bi2r_kikprjp537f   = vacmjbyuw8jriztdg
                    & (f7t_bak0dfaq3);




  wire gofb_xvfjsatvpae6l = (ipq0f4_yvmml7o06891 & fk7qm80i_py_6);
  assign tj9rezp6j0u0mvddq   =  gofb_xvfjsatvpae6l & (~bi2r_kikprjp537f);

  
  

  wire zx62ukmv5eyf3 = ipq0f4_yvmml7o06891 & p4jgl36nmqe8ud7_g4i7;

  wire  v47xf8kt__ckq6pm8ic = o9vvv_q4ikz_2yp0w & y40x_uwnqs6f;
  assign zl3w_sym4l3ca   = v47xf8kt__ckq6pm8ic  
                        & (~bi2r_kikprjp537f) & (~tj9rezp6j0u0mvddq) ;

  
  

  wire yopdnmqpounix9 = o9vvv_q4ikz_2yp0w & c1ilkc2r6es72c5h2vcc;



  wire f80c9kfaqm_llph13deg = ll0_hbknv5bc_8mxvx5c & tdg7ccg5dltr5l9s;
  wire zqdvxq2z9p52_   = f80c9kfaqm_llph13deg 
                        & (~bi2r_kikprjp537f) & (~zl3w_sym4l3ca) & (~tj9rezp6j0u0mvddq)  
                        ;

  

  wire   yukowgvwkyqgijo2fv3 = q89zlvtwzxkjd6h5k;
  wire qa7oqpph4a7i7xf6re   = ju3gksnn2mup5h81eh28 & yukowgvwkyqgijo2fv3 
                         & (~bi2r_kikprjp537f) & (~zl3w_sym4l3ca) & (~tj9rezp6j0u0mvddq) 
                         & (~zqdvxq2z9p52_)
                         ;

  wire   o8w0jo3q_y9x6ehb9 = v7f1q1_fp5fc8b_u;
  wire pyka5_r6eb9j1   = lanyt81iat_ws21fv & o8w0jo3q_y9x6ehb9 
                         & (~qa7oqpph4a7i7xf6re) & (~bi2r_kikprjp537f) & (~zl3w_sym4l3ca) & (~tj9rezp6j0u0mvddq) 
                         & (~zqdvxq2z9p52_)
                         ;

  wire   po7du4hib7cjmxyp = vmwegtj2c0zt7rilpw;
  wire ykowh_zywv6woag   = nz5iij5cadsnx4fokudqbo & po7du4hib7cjmxyp 
                         & (~pyka5_r6eb9j1) & (~qa7oqpph4a7i7xf6re) & (~bi2r_kikprjp537f) & (~zl3w_sym4l3ca) & (~tj9rezp6j0u0mvddq) 
                         & (~zqdvxq2z9p52_)
                         ;




  
  
  
  
  
  
  
  
  
  
  
  
  

  
  
  
  

  
  
  
  




 wire ehbp4qn2mf9zuvt;

  assign srufsypxvg1hqxwmw0y = 
             p7ah58va5_2njbtv ? 
              {
                p0i2i3v3j1tclelx51,
                (~p0i2i3v3j1tclelx51),
                1'b1,
                1'b0,
                u981qrwkgi5h0e72b__gg19w,
                1'b0
              } :
             ({jwxxo5dwz741q1{bi2r_kikprjp537f}} & 
              {
                pxbhqh6yl6hotx,
                toib7p7z_deij2b,
                p_2daj_9kqsf0ekr101,
                djb42mrmnunfufgxzh,
                vqldrx_4vk7av570m8fv,
                1'b0
              }) 

              ;

  assign {
         zeseql2htbxpugyu5_j   
        ,al3t866kz4po45vfuyjy  
        ,xutsaulafh4onxtthm8n
        ,me7unt7fapqqhtc6epso
        ,m2as3qe7miuhj662j1zvt
        ,ehbp4qn2mf9zuvt
        } = yhopxd2wrapvsuiglom;




  wire                         qzj6si9v4vdhaoi;
  wire                         gbay31fa2brf2;
  wire                         zhsv0cp6_4  ;
  wire                         yydetudxf41g;
  wire [64-1:0]        um__n7hbw6b;
  wire [5-1:0]                 vs4ta1kq798ck;
  wire [5-1:0] afgjc4gl7iktp1cf;
  wire                         gvycxr45os1jw;
  wire [4-1:0]  umd6fz93tap ;




  assign dlogavn_28q56zummtut = bi2r_kikprjp537f & gbay31fa2brf2 ;

  assign c1ilkc2r6es72c5h2vcc = zl3w_sym4l3ca & gbay31fa2brf2;
  
  assign p4jgl36nmqe8ud7_g4i7 = tj9rezp6j0u0mvddq & gbay31fa2brf2;
  assign qloskxsiztazdeq2ad95i = zqdvxq2z9p52_ & gbay31fa2brf2;
  assign tymuflph4h7mej5umh86 = qa7oqpph4a7i7xf6re & gbay31fa2brf2;
  assign b1eabu9fa3jnjln5tc = pyka5_r6eb9j1 & gbay31fa2brf2;
  assign bz1hc72g_22hgoqs8 = ykowh_zywv6woag & gbay31fa2brf2;

  assign qzj6si9v4vdhaoi = 
                        (bi2r_kikprjp537f  ) 
                      | (qa7oqpph4a7i7xf6re ) 
                      | (pyka5_r6eb9j1 ) 
                      | (ykowh_zywv6woag ) 
                      | (zl3w_sym4l3ca  ) 
                      | (tj9rezp6j0u0mvddq  ) 
                      | (zqdvxq2z9p52_)
                         ;

  wire [64-1:0] fiyi5b17rt4d4gp6yswwk = yhfc75p_gcdigu;
  wire [64-1:0] fs7rjgrwae0s323axaf7j = {{64-64{1'b0}},l3sefagtx4ai4ljb};
  wire [64-1:0] vf8up74ci1lxgxfzd_5p = {{64-64{1'b0}},wyhg5n7dklr59dxgm_bs};
  wire [64-1:0] timv678rmmwnyufgnbcz = {{64-64{1'b0}},px17v86p_7_1fdvm1w};

  assign um__n7hbw6b  = 

                        ({64{bi2r_kikprjp537f}} & fiyi5b17rt4d4gp6yswwk ) 
                      | ({64{qa7oqpph4a7i7xf6re}} & {{64-64{1'b0}},c5csn3nczo8zlvq621sy}) 
                      | ({64{pyka5_r6eb9j1}} & {{64-64{1'b0}},nt0ndhbk6x29ae8da95}) 
                      | ({64{ykowh_zywv6woag}} & {wctv6a1mmq6dtwsg9n}) 
                      
                      | ({64{zl3w_sym4l3ca}} & fs7rjgrwae0s323axaf7j) 
                      | ({64{tj9rezp6j0u0mvddq}} & vf8up74ci1lxgxfzd_5p) 
                      | ({64{zqdvxq2z9p52_}} & timv678rmmwnyufgnbcz) 
                         ;

  assign vs4ta1kq798ck  = 
                        ({5{bi2r_kikprjp537f}} & wk41j07s3anl9_t)
                      | ({5{qa7oqpph4a7i7xf6re}} & rd0rvbiicactt4sbf) 
                      | ({5{pyka5_r6eb9j1}} & ri8f9g_paihffhz9_8qgu) 
                      | ({5{ykowh_zywv6woag}} & onijw658b2__et8fr1has) 
                    ;
  assign zhsv0cp6_4   = 
                        (bi2r_kikprjp537f & psylshnv8k3qqz5i) 
                      | (qa7oqpph4a7i7xf6re & h5w2di84ketcahr4) 
                      | (pyka5_r6eb9j1 & ik4ulvmx89l0u0ko) 
                      | (ykowh_zywv6woag & ys8dsx5hx_injk9b) 
                      | (zl3w_sym4l3ca & bjn5x3u7v4u3rm6d) 
                      | (tj9rezp6j0u0mvddq & cbr_upfu_0ywren54f) 
                      | (zqdvxq2z9p52_ & a3g162j6o30b4qdpd_z) 
                         ;

  assign afgjc4gl7iktp1cf = 

                        ({5{bi2r_kikprjp537f}} & v2fkznl9m7dtfymx) 
                      | ({5{qa7oqpph4a7i7xf6re}} & f63hhh0gzajzsiyjd8cqb) 
                      | ({5{pyka5_r6eb9j1}} & nfozodmnsmlv22fi3oe) 
                      | ({5{ykowh_zywv6woag}} & nq8gzr65b3p_cdc52lshh) 
                      | ({5{zl3w_sym4l3ca}} & ejlcmcywa2ghgwvj) 
                      | ({5{tj9rezp6j0u0mvddq}} & gof9x1lyu2n5rnf) 
                      | ({5{zqdvxq2z9p52_}} & ggpqgd6b8zuelz8) 
                         ;


  assign gvycxr45os1jw = 

                        (bi2r_kikprjp537f & oy1tzeyrsbr3bg7dr9u)
                      | (qa7oqpph4a7i7xf6re & vf6etunsloifr12azv4he6 & !h5w2di84ketcahr4) 
                      | (pyka5_r6eb9j1 & ltzlg4gy4noc9555li & !ik4ulvmx89l0u0ko) 
                      | (ykowh_zywv6woag & bp90ffmjkj3u4__poo & !ys8dsx5hx_injk9b) 
                      | (zl3w_sym4l3ca & qlykdb48c89hfbq5l3v & !bjn5x3u7v4u3rm6d) 
                      | (tj9rezp6j0u0mvddq & utfce4yxn08kh9t & !cbr_upfu_0ywren54f) 
                      | (zqdvxq2z9p52_ & z5s1cielsyyeza34h & !a3g162j6o30b4qdpd_z) 
                         ;
  assign umd6fz93tap = 

                        ({4{bi2r_kikprjp537f}} & zl0t249z3fcwyj4puu) 
                      | ({4{qa7oqpph4a7i7xf6re}} & g5gmidj6od8k58avl_h9y) 
                      | ({4{pyka5_r6eb9j1}} & u7vn3gjmd4owzsi7tk) 
                      | ({4{ykowh_zywv6woag}} & zakjetcb_4mzmn_bchz) 
                      | ({4{zl3w_sym4l3ca}} & josyt39cvr3gignopao) 
                      | ({4{tj9rezp6j0u0mvddq}} & ubk6j4rwgfrf5ryn1ibp) 
                      | ({4{zqdvxq2z9p52_}} & jb9locwfccqzb06jjon) 
                         ;




  assign yydetudxf41g = 1'b0
                         | (bi2r_kikprjp537f  & rpnvo9xxx6nke515) 
                         | (qa7oqpph4a7i7xf6re & gjoru9khthrg8j6pfamu) 
                         | (pyka5_r6eb9j1 & mvneatl67xbzspkpyi1) 
                         | (ykowh_zywv6woag & szgl0r6i254qax8jkjr) 
                      ;





  wire mc19e3318 = gvycxr45os1jw;



  wire iezr51kzroh = zhsv0cp6_4;







  assign gbay31fa2brf2 = 
       (mc19e3318 ? ar7xgugq1a_pz7b82ds : 1'b1)

       ;





  wire xywba85npeg96 = gbay31fa2brf2 & qzj6si9v4vdhaoi & (
                        (zl3w_sym4l3ca )
                      | (tj9rezp6j0u0mvddq )
                      | (bi2r_kikprjp537f )
                      | (zqdvxq2z9p52_ )
                     );
  assign p1jdw9loxkz60taq_vkp_3 = mc19e3318 & qzj6si9v4vdhaoi;

  assign jwwku_el5h5h2lx6e0kyi  = um__n7hbw6b ;
  assign zt19omidnr_zyp2gc3bywfb = vs4ta1kq798ck;
  assign v19st7vd9_bi485e6ak0 = yydetudxf41g;
  assign gccap1c6hft7o1z7esm   = gvycxr45os1jw;
  assign vjhpkmep8g_u_cizhsw = afgjc4gl7iktp1cf;




  assign eo5skx1ygvzuasbjgnyl = umd6fz93tap;


  assign mxa77etukhs8o_5z6962l19 = iezr51kzroh & xywba85npeg96;

  assign xd2ftroj1i79g4derw = qzj6si9v4vdhaoi & gbay31fa2brf2;
  assign qoxd9f57dl083f6cm  = umd6fz93tap;

endmodule                                      
























module sdt_3ftsvyvhysb2f7uduiazuiu(



  input                         y40x_uwnqs6f   ,
  input                         fk7qm80i_py_6   ,
  input                         f7t_bak0dfaq3   ,

  input                         qlykdb48c89hfbq5l3v ,
  input                         utfce4yxn08kh9t ,
  input                         oy1tzeyrsbr3bg7dr9u ,
  input                         rpnvo9xxx6nke515 ,
  input                         tdg7ccg5dltr5l9s,
  input                         z5s1cielsyyeza34h,

  input [5-1:0] ejlcmcywa2ghgwvj ,
  input [5-1:0] gof9x1lyu2n5rnf ,
  input [5-1:0] v2fkznl9m7dtfymx ,
  input [5-1:0] ggpqgd6b8zuelz8,

  input                          ll0_hbknv5bc_8mxvx5c, 
  output                         qloskxsiztazdeq2ad95i, 
  input  [64-1:0]        px17v86p_7_1fdvm1w,
  input  [4 -1:0] jb9locwfccqzb06jjon,
  input                          a3g162j6o30b4qdpd_z , 

  input                          q89zlvtwzxkjd6h5k, 
  input                          gjoru9khthrg8j6pfamu, 
  input                          vf6etunsloifr12azv4he6, 
  input [5-1:0]  f63hhh0gzajzsiyjd8cqb,
  input                          v7f1q1_fp5fc8b_u, 
  input                          mvneatl67xbzspkpyi1, 
  input                          ltzlg4gy4noc9555li, 
  input [5-1:0]  nfozodmnsmlv22fi3oe,
  input                          vmwegtj2c0zt7rilpw, 
  input                          szgl0r6i254qax8jkjr, 
  input                          bp90ffmjkj3u4__poo, 
  input [5-1:0]  nq8gzr65b3p_cdc52lshh,

  input                          ju3gksnn2mup5h81eh28, 
  output                         tymuflph4h7mej5umh86, 
  input  [64-1:0]        c5csn3nczo8zlvq621sy ,
  input  [5-1:0]                 rd0rvbiicactt4sbf,
  input  [4 -1:0] g5gmidj6od8k58avl_h9y ,
  input                          h5w2di84ketcahr4  , 

  input                          lanyt81iat_ws21fv, 
  output                         b1eabu9fa3jnjln5tc, 
  input  [64-1:0]        nt0ndhbk6x29ae8da95,
  input  [5-1:0]                 ri8f9g_paihffhz9_8qgu,
  input  [4 -1:0] u7vn3gjmd4owzsi7tk,
  input                          ik4ulvmx89l0u0ko ,

  input                          nz5iij5cadsnx4fokudqbo,
  output                         bz1hc72g_22hgoqs8,
  input  [64-1:0]        wctv6a1mmq6dtwsg9n,
  input  [5-1:0]                 onijw658b2__et8fr1has,
  input  [4 -1:0] zakjetcb_4mzmn_bchz,
  input                          ys8dsx5hx_injk9b ,





  input                         ipq0f4_yvmml7o06891, 
  output                        p4jgl36nmqe8ud7_g4i7, 
  input  [64-1:0]       wyhg5n7dklr59dxgm_bs,
  input                         cbr_upfu_0ywren54f,
  input  [4-1:0] ubk6j4rwgfrf5ryn1ibp,


  
  
  input                         o9vvv_q4ikz_2yp0w, 
  output                        c1ilkc2r6es72c5h2vcc, 
  input  [64-1:0]       l3sefagtx4ai4ljb,
  input                         bjn5x3u7v4u3rm6d,
  input  [4-1:0] josyt39cvr3gignopao,




  input                          ret9emt0e4v60a6cwap10, 
  output                         l5447rrn286zsq9mt6k, 
  input  [64-1:0]        fg4h6qs_th28xw7il0,
  input  [4 -1:0] q7ns1l4tc_kuf5az3u,
  input                          h_ld26vo8tpdty , 
  input                          p_2daj_9kqsf0ekr101 ,
  input                          djb42mrmnunfufgxzh ,
  input  [64 -1:0]  vqldrx_4vk7av570m8fv,
  input  [64 -1:0]    zhwwio_mprrvjud04     ,
  input                          pxbhqh6yl6hotx     , 
  input                          toib7p7z_deij2b     , 
  input  [4:0]                   dufpf9uw3i8khwmvb2h,
  input                          p7ah58va5_2njbtv,
  input [64-1:0]    u981qrwkgi5h0e72b__gg19w,
  input                          p0i2i3v3j1tclelx51,




  output p1jdw9loxkz60taq_vkp_3, 
  input  ar7xgugq1a_pz7b82ds, 
  output [64-1:0] jwwku_el5h5h2lx6e0kyi,
  output [5-1:0] zt19omidnr_zyp2gc3bywfb,
  output [5 -1:0] vjhpkmep8g_u_cizhsw,
  output [4-1:0] eo5skx1ygvzuasbjgnyl,
  output v19st7vd9_bi485e6ak0,
  output gccap1c6hft7o1z7esm,






  output                          gqat5ctwgmxi8n_5z03tivvpgqx6j5kb, 
  output  [4 -1:0] zmotzlbzlmuf2isjtqn2h8beel09 ,

  output                          vi7663z7hxlc4ngkh1_yfoxfpvbiq, 
  output  [4 -1:0] ql2r_7apgocbap5k7ucf5a673x7v ,


  output                          bm0yhprev2rfpkaztktaxtnq7f8q0bp, 
  output  [4 -1:0] i2kgxrwehfoyscnln10tc70_omph,


  output                          gkb40bm903wc32_2zjmb0l25g21p7, 
  output  [4 -1:0] yu_1foait_ukyv14b73xepo_1mj31mu,
  output                          scom2gns1t5jrniqayb84g_h2a1zaxbv, 
  output  [4 -1:0] xpvibysxiip4tytx5_ry26i78ce4j4,
  output                          ky7mnv5l4jl0v17ox278fwktul3qti, 
  output  [4 -1:0] a9_1a439ejmx35qe2g8yihj84g5,
  output                          rhx_hd60cwxftbqnr_uhlcmbab17eeue, 
  output  [4 -1:0] l_w88r7i0zq6u0xtcywbwzu__s,


  output  z2qyay491938ppnlxuc,
  input   pbtolkl953sk14id0iy,
  output  zeseql2htbxpugyu5_j,
  output  al3t866kz4po45vfuyjy,
  output  xutsaulafh4onxtthm8n , 
  output  me7unt7fapqqhtc6epso , 
  output [64-1:0] m2as3qe7miuhj662j1zvt,



  output czyvvnzs3y3orktdmdfec8yla_1y,
  output [4 -1:0] o_tztjh1zql5hzdma85okucmgxh, 


  input  gf33atgy,
  input  ru_wi
  );


  wire                        cuzanreq1u8ev47iova; 
  wire                        pg0v_24f5gtcbo20w; 
  wire[64-1:0]        vuy4dkld2kpsy45c ; 
  wire [4-1:0] kbqrg_4bxmxn7b7up8 ; 
  wire                        mj86rmgsgeu75euwgxk2  ; 

  wire                        wgcdhfocgyd9bovps; 
  wire                        bpgjhz125ozfoh_yq_cze; 
  wire[64-1:0]        d7w4y25gmfw83aoc9 ; 
  wire [4-1:0] ppz9xrdau3m7w60f ; 
  wire                        zonryv578qcpvne  ; 

  wire                        noee4sp5nj0yu67gse95w7; 
  wire                        mk4t4nfrjj6kszdmlvx; 
  wire[64-1:0]        dmle1ahfbwbgdsus3urzc ; 
  wire [4-1:0] w8y2hbgpdiw40ue7 ; 
  wire                        uhlmwyl5pyhbili8  ; 


  wire                          zsgxtf4008xy__uvhtb ;
  wire                          s82s_18977u8wf_m03xle ;
  wire                          vo1wq92xi41ixlir3ymlrb6;
  wire                          tw0q0kvd274notuz0datc8 ;
  wire  [64 -1:0]  iqbltqegpktkmdbk_wp4o;
  wire  [64 -1:0]    w5aw4cypvoskbhpdkq     ;
  wire                          wp0j2jfw1xi0w3ty     ; 
  wire                          f9l2d7z_qipj5cefpi     ; 
  wire  [4:0]                   y_4zkek_lck4fr6cpsm  ;






  wire                        qcz2i1lzeluodju99g0; 
  wire                        vruj1aci16ru7rc5dr; 
  wire[64-1:0]        t4z031uv53p1rqo1lm9 ; 
  wire [4-1:0] mazfnbz00ya1f7wlojtz ; 
  wire                        fuhx6ea_0i4biqppt  ; 

  wire                        ahjuy_x5m5qihqghx7hpw; 
  wire                        u4pj98i_6_wxhdnzq; 
  wire[64-1:0]        hxhsc9xkvilz_l3_1nn ; 
  wire [4-1:0] zh2qii8n5s7pyqavvlc ; 
  wire                        i8n5vfo_dfg36lk7h  ; 
  wire [4:0]                  edx95k3p7jv9r96kacf; 
  wire                        jwn0vy3w73wvchqf2e_; 
  wire                        cumuievj81yzsmwme5vnb; 
  wire[64-1:0]        q9c69qv2eiojvdikkie ; 
  wire [4-1:0] tgrf16ko9nguy1ze ; 
  wire                        t50b3x1hdgvvw_k  ; 
  wire [4:0]                  t52jbjpudt9o21r24qxlx; 
  wire                        sg49_hmdhls607ljc1mz; 
  wire                        y9vl_d4wtjr06n0dyt; 
  wire[64-1:0]        g8ezms55j8q3tkse3igad ; 
  wire [4-1:0] uwu0k4ysqaaf7cq1 ; 
  wire                        l23pvox21yl49eb  ; 
  wire [4:0]                  apng_vbetdgo_5t3dis; 


  assign gqat5ctwgmxi8n_5z03tivvpgqx6j5kb = cuzanreq1u8ev47iova; 
  assign zmotzlbzlmuf2isjtqn2h8beel09  = kbqrg_4bxmxn7b7up8 ;
  assign vi7663z7hxlc4ngkh1_yfoxfpvbiq = wgcdhfocgyd9bovps; 
  assign ql2r_7apgocbap5k7ucf5a673x7v  = ppz9xrdau3m7w60f ;
  assign bm0yhprev2rfpkaztktaxtnq7f8q0bp = noee4sp5nj0yu67gse95w7; 
  assign i2kgxrwehfoyscnln10tc70_omph  = w8y2hbgpdiw40ue7 ;
  assign gkb40bm903wc32_2zjmb0l25g21p7 = ahjuy_x5m5qihqghx7hpw; 
  assign yu_1foait_ukyv14b73xepo_1mj31mu  = zh2qii8n5s7pyqavvlc ;
  assign scom2gns1t5jrniqayb84g_h2a1zaxbv = jwn0vy3w73wvchqf2e_; 
  assign xpvibysxiip4tytx5_ry26i78ce4j4  = tgrf16ko9nguy1ze ;
  assign ky7mnv5l4jl0v17ox278fwktul3qti = sg49_hmdhls607ljc1mz; 
  assign a9_1a439ejmx35qe2g8yihj84g5  = uwu0k4ysqaaf7cq1 ;
  assign rhx_hd60cwxftbqnr_uhlcmbab17eeue = qcz2i1lzeluodju99g0; 
  assign l_w88r7i0zq6u0xtcywbwzu__s  = mazfnbz00ya1f7wlojtz ;



uh_y21ipql6al1c4qkqfokr_0yd zwh9pl8_718zr38rl_h3ehienjcobl74(



  .r25vjm_g303hv5mr__oydfc50s_6(ipq0f4_yvmml7o06891), 
  .q3nebxbyx8x_n2wgt90jxx5ppnlbuzt(p4jgl36nmqe8ud7_g4i7), 
  .l9uyi_93i_vkb6davalokxbus3edyu (wyhg5n7dklr59dxgm_bs ),
  .kptoalwjf0vnjxpubirzzg8r1l0_hk7 (ubk6j4rwgfrf5ryn1ibp ),
  .qd2ehv6u5ipjg2sd3swjn38uuab  (cbr_upfu_0ywren54f  ), 

  .x0wwmbj55rz1_gzemtenuutvu4f5gtbr(o9vvv_q4ikz_2yp0w), 
  .tjf2j_x0_19wvbnushzloo4vpibe0q(c1ilkc2r6es72c5h2vcc), 
  .jcur3i2c0we7b6x5ms3vw9himw35v (l3sefagtx4ai4ljb ),
  .vmujqgbzxn6hqc5j49ufmtewa7 (josyt39cvr3gignopao ),
  .x74i2xb96e9fui_1revcqt088tm0hf  (bjn5x3u7v4u3rm6d  ), 


  .wqlni2o6ysdnyxmiesc2c9nx1nhsidr(ret9emt0e4v60a6cwap10), 
  .bx1s0daa65s6eao0yo05dgpi6o_6e7(l5447rrn286zsq9mt6k), 
  .cefmw490fob0947fn0zxl51_fkeb (fg4h6qs_th28xw7il0 ),
  .csw73tw17ceolm9eifmbhd887zfa (q7ns1l4tc_kuf5az3u ),
  .fu2trk07aq8pgduthe_h3zskathrh  (h_ld26vo8tpdty  ), 
  .p5laf3iz7k000k42fpww1tjw97c514pj(dufpf9uw3i8khwmvb2h),

  .kq64hafe_jmlm63rt4w15_qnftr01(p_2daj_9kqsf0ekr101),
  .en8f11yeo7j9u54v7agnvuncx9kha(djb42mrmnunfufgxzh),
  .pqeyh89bzfwni86npwrcnmz1fjtb2dhfj(1'b0),
  .os5_rc90_7gawcz0efrilvhb5wo74r9(1'b0),
  .zllz_u37t659z507dtl4d906nsg35(vqldrx_4vk7av570m8fv),
  .i5m1rrdydixypqcxzmalcomh     (zhwwio_mprrvjud04     ),
  .laifryt4bl834uov7isyxe_4uk3_d     (pxbhqh6yl6hotx     ),
  .yvw2qnvbiajkt2mcxp4j4xqiucb8     (toib7p7z_deij2b     ),



  .obli6e3v4_8bjrltqdv6v18stt0fev4(ju3gksnn2mup5h81eh28), 
  .tb6a57t86vwitea0x8780ksclx8d4(tymuflph4h7mej5umh86), 
  .jomr8wem988b32tidmg2zkgiqgl6 (c5csn3nczo8zlvq621sy ),
  .boxfq4ncnb8czlmq7p4msay3wg7o4 (g5gmidj6od8k58avl_h9y ),
  .k98w6098j0wekfd9wjqjkmtslxo  (h5w2di84ketcahr4  ), 
  .jz83wrre56m2b7vf1dnwnnu8lme(rd0rvbiicactt4sbf), 
  .vo9o42ohfekmv2b390b9ovdxs7hswv(lanyt81iat_ws21fv), 
  .xvr_92a8rcvf2quyrmigj7fzuftq(b1eabu9fa3jnjln5tc), 
  .yhqkr966fkfranbq6mys4_itfdsz8 (nt0ndhbk6x29ae8da95 ),
  .ktpgkhezvy18ox4t8b5xhresqcnvqp6 (u7vn3gjmd4owzsi7tk ),
  .jqaxpjo0j1mrf8casph8bqvmhaf  (ik4ulvmx89l0u0ko  ), 
  .d4xh57em8iunsz9w5_jruofpuezsh(ri8f9g_paihffhz9_8qgu), 
  .z0p5c0vl91tsjk1lmt8kxat0kig3dlom(nz5iij5cadsnx4fokudqbo), 
  .kqhgic2ez1gu2b308vr7gayeops(bz1hc72g_22hgoqs8), 
  .or2q_8b_zdv2o7h7ol6rtfs9p7sqzx9 (wctv6a1mmq6dtwsg9n ),
  .zo0u9kjy8fmzeh_qnut3gcckfj_ (zakjetcb_4mzmn_bchz ),
  .emdo9xkvazh0e830c3tezq85cr  (ys8dsx5hx_injk9b  ), 
  .c90btjrwqlw7w7j9o1twzgjt43njm3wg(onijw658b2__et8fr1has), 
  .wqn_diiyx7s7t037qfg_nkqdnix(ll0_hbknv5bc_8mxvx5c), 
  .aeqpr5hrp251jp0yxm1vcqjoftohs(qloskxsiztazdeq2ad95i), 
  .vqzbvg_jyxunlaurqlpwhp34u_jx0 (px17v86p_7_1fdvm1w ),
  .t1tkrihuzsa8iq9pywbo4a3ktie7wn4 (jb9locwfccqzb06jjon ),
  .ytkv6_mmnisydnwtk48igroblctc  (a3g162j6o30b4qdpd_z  ), 




  .gqat5ctwgmxi8n_5z03tivvpgqx6j5kb(cuzanreq1u8ev47iova), 
  .n0cmggtax9qzrd4qsy1cdbik144lmx(pg0v_24f5gtcbo20w), 
  .y4aoa0ok7ylngx_33gfqr0g1md0g8dj (vuy4dkld2kpsy45c ),
  .zmotzlbzlmuf2isjtqn2h8beel09 (kbqrg_4bxmxn7b7up8 ),
  .vo2fj15n058l2wpxbodnsdqxwkdn08  (mj86rmgsgeu75euwgxk2  ), 

  .vi7663z7hxlc4ngkh1_yfoxfpvbiq(wgcdhfocgyd9bovps), 
  .rhwm1lw0wyhvdhss4f3p_v5zkroo(bpgjhz125ozfoh_yq_cze), 
  .vsgctu8mzjw91ryb865p9r7s8fp (d7w4y25gmfw83aoc9 ),
  .ql2r_7apgocbap5k7ucf5a673x7v (ppz9xrdau3m7w60f ),
  .sei0me3z77b60zu8tfykejc6_w  (zonryv578qcpvne  ), 


  .bm0yhprev2rfpkaztktaxtnq7f8q0bp(noee4sp5nj0yu67gse95w7), 
  .f_7j356ybgmsh86n3umtlmih2ee8c5(mk4t4nfrjj6kszdmlvx), 
  .ktwrzuv2gg846pksncc26g4y0pe1h (dmle1ahfbwbgdsus3urzc ),
  .i2kgxrwehfoyscnln10tc70_omph (w8y2hbgpdiw40ue7 ),
  .xp4xfk612_1jfargldlbq2rjb  (uhlmwyl5pyhbili8  ), 
  .lrojclgmk96728ugf1xss07x7gzfgls(y_4zkek_lck4fr6cpsm),
  .rdsej_3e3o2bh3ld92ygwf707k988       (zsgxtf4008xy__uvhtb),
  .eitel8xkigdj96m3f89nsi2w_71pvf       (s82s_18977u8wf_m03xle),
  .eovnqir46kp7wnkzr0btiuicjboull      (vo1wq92xi41ixlir3ymlrb6),
  .qc6yp7yoe_bjq2am96mg0sizkq7os       (tw0q0kvd274notuz0datc8),
  .lo4an3qbdgmg6hqsqosvvk8dwctnn1wy6c      (iqbltqegpktkmdbk_wp4o),
  .xedi2t9w7jc8_rstzke961dl4l7           (w5aw4cypvoskbhpdkq     ),
  .az7mzc_81tib2dpb5d3a70_wdp73f           (wp0j2jfw1xi0w3ty     ),
  .oopk92ymqbivd2dxs85nt1ly5ccn           (f9l2d7z_qipj5cefpi     ),


  .gkb40bm903wc32_2zjmb0l25g21p7(ahjuy_x5m5qihqghx7hpw), 
  .j0l8i3eed1ek492qjzm9uejf41sz(u4pj98i_6_wxhdnzq), 
  .yyasjan35_68l3cq8a3ioaew9bbhr (hxhsc9xkvilz_l3_1nn ),
  .yu_1foait_ukyv14b73xepo_1mj31mu (zh2qii8n5s7pyqavvlc ),
  .pdkr3e96qk7jfuv5c8967qald7p  (i8n5vfo_dfg36lk7h  ), 
  .xfz4lyb4bxla1gb3kuqf0gcek1_r8yz(edx95k3p7jv9r96kacf), 
  .scom2gns1t5jrniqayb84g_h2a1zaxbv(jwn0vy3w73wvchqf2e_), 
  .jzh4duikrv004mprz7zksk2dh9ty72(cumuievj81yzsmwme5vnb), 
  .geun5etyjtjsnydbal2egw52gf34 (q9c69qv2eiojvdikkie ),
  .xpvibysxiip4tytx5_ry26i78ce4j4 (tgrf16ko9nguy1ze ),
  .kng9rvszc8o8ob5v1_ak0ipg9lgbku  (t50b3x1hdgvvw_k  ), 
  .avrbak7i2ou0is2fulrxcpx4b8qjfwus(t52jbjpudt9o21r24qxlx), 
  .ky7mnv5l4jl0v17ox278fwktul3qti(sg49_hmdhls607ljc1mz), 
  .wt906274r_7subjpzosffvtc_8lbfu(y9vl_d4wtjr06n0dyt), 
  .fsr9hzh57oj6r29w8_fdfss2962 (g8ezms55j8q3tkse3igad ),
  .a9_1a439ejmx35qe2g8yihj84g5 (uwu0k4ysqaaf7cq1 ),
  .n412jv5dj1tvgdf8jls7u2bjvh  (l23pvox21yl49eb  ), 
  .ke2zqim9rdwj_bmursxrbh8ga08qo(apng_vbetdgo_5t3dis), 
  .rhx_hd60cwxftbqnr_uhlcmbab17eeue(qcz2i1lzeluodju99g0), 
  .gm94l7jeucs5_57r7b1ghqbrvubvg(vruj1aci16ru7rc5dr), 
  .wtj2dgdc6vyaj4ptn464rhnsgz1 (t4z031uv53p1rqo1lm9 ),
  .l_w88r7i0zq6u0xtcywbwzu__s (mazfnbz00ya1f7wlojtz ),
  .om2j1tmzbckjwmzuoudwijwh6gh_ig  (fuhx6ea_0i4biqppt  ), 



  .gf33atgy  (gf33atgy  ),
  .ru_wi(ru_wi)
  );




  uv355zczoyyqi_qujlvi a7loowtd3371ybmyeuxfzj(

    .vacmjbyuw8jriztdg    (noee4sp5nj0yu67gse95w7 ),
    .dlogavn_28q56zummtut    (mk4t4nfrjj6kszdmlvx ),
    .yhfc75p_gcdigu     (dmle1ahfbwbgdsus3urzc  ),
    .zl0t249z3fcwyj4puu     (w8y2hbgpdiw40ue7  ),
    .psylshnv8k3qqz5i      (uhlmwyl5pyhbili8   ),
    .pxbhqh6yl6hotx       (wp0j2jfw1xi0w3ty     ),
    .toib7p7z_deij2b       (f9l2d7z_qipj5cefpi     ),
    .vqldrx_4vk7av570m8fv  (iqbltqegpktkmdbk_wp4o ),
    .zhwwio_mprrvjud04       (w5aw4cypvoskbhpdkq      ),
    .p_2daj_9kqsf0ekr101   (zsgxtf4008xy__uvhtb  ),
    .djb42mrmnunfufgxzh   (s82s_18977u8wf_m03xle  ),
    .wk41j07s3anl9_t    (y_4zkek_lck4fr6cpsm  ),
    .p7ah58va5_2njbtv      (p7ah58va5_2njbtv     ), 
    .u981qrwkgi5h0e72b__gg19w (u981qrwkgi5h0e72b__gg19w), 
    .p0i2i3v3j1tclelx51     (p0i2i3v3j1tclelx51    ), 
    .y40x_uwnqs6f         (y40x_uwnqs6f       ),
    .qlykdb48c89hfbq5l3v       (qlykdb48c89hfbq5l3v     ),
    .ejlcmcywa2ghgwvj       (ejlcmcywa2ghgwvj     ),
    .fk7qm80i_py_6         (fk7qm80i_py_6       ),
    .utfce4yxn08kh9t       (utfce4yxn08kh9t     ),
    .gof9x1lyu2n5rnf       (gof9x1lyu2n5rnf     ),
    .f7t_bak0dfaq3         (f7t_bak0dfaq3       ),
    .oy1tzeyrsbr3bg7dr9u       (oy1tzeyrsbr3bg7dr9u     ),
    .rpnvo9xxx6nke515       (rpnvo9xxx6nke515     ),
    .v2fkznl9m7dtfymx       (v2fkznl9m7dtfymx     ),
    .tdg7ccg5dltr5l9s      (tdg7ccg5dltr5l9s  ),
    .ggpqgd6b8zuelz8    (ggpqgd6b8zuelz8),
    .z5s1cielsyyeza34h    (z5s1cielsyyeza34h),


    .q89zlvtwzxkjd6h5k   (q89zlvtwzxkjd6h5k   ), 
    .gjoru9khthrg8j6pfamu (gjoru9khthrg8j6pfamu ), 
    .vf6etunsloifr12azv4he6 (vf6etunsloifr12azv4he6 ), 
    .f63hhh0gzajzsiyjd8cqb (f63hhh0gzajzsiyjd8cqb ),
    .v7f1q1_fp5fc8b_u   (v7f1q1_fp5fc8b_u   ), 
    .mvneatl67xbzspkpyi1 (mvneatl67xbzspkpyi1 ), 
    .ltzlg4gy4noc9555li (ltzlg4gy4noc9555li ), 
    .nfozodmnsmlv22fi3oe (nfozodmnsmlv22fi3oe ),
    .vmwegtj2c0zt7rilpw   (vmwegtj2c0zt7rilpw   ), 
    .szgl0r6i254qax8jkjr (szgl0r6i254qax8jkjr ), 
    .bp90ffmjkj3u4__poo (bp90ffmjkj3u4__poo ), 
    .nq8gzr65b3p_cdc52lshh (nq8gzr65b3p_cdc52lshh ),

    .ju3gksnn2mup5h81eh28   (ahjuy_x5m5qihqghx7hpw), 
    .tymuflph4h7mej5umh86   (u4pj98i_6_wxhdnzq), 
    .c5csn3nczo8zlvq621sy    (hxhsc9xkvilz_l3_1nn ),
    .g5gmidj6od8k58avl_h9y    (zh2qii8n5s7pyqavvlc ),
    .h5w2di84ketcahr4     (i8n5vfo_dfg36lk7h  ), 
    .rd0rvbiicactt4sbf   (edx95k3p7jv9r96kacf), 

    .lanyt81iat_ws21fv   (jwn0vy3w73wvchqf2e_), 
    .b1eabu9fa3jnjln5tc   (cumuievj81yzsmwme5vnb), 
    .nt0ndhbk6x29ae8da95    (q9c69qv2eiojvdikkie ),
    .u7vn3gjmd4owzsi7tk    (tgrf16ko9nguy1ze ),
    .ik4ulvmx89l0u0ko     (t50b3x1hdgvvw_k  ), 
    .ri8f9g_paihffhz9_8qgu   (t52jbjpudt9o21r24qxlx), 
                         
    .nz5iij5cadsnx4fokudqbo   (sg49_hmdhls607ljc1mz),
    .bz1hc72g_22hgoqs8   (y9vl_d4wtjr06n0dyt),
    .wctv6a1mmq6dtwsg9n    (g8ezms55j8q3tkse3igad ),
    .zakjetcb_4mzmn_bchz    (uwu0k4ysqaaf7cq1 ),
    .ys8dsx5hx_injk9b     (l23pvox21yl49eb  ),
    .onijw658b2__et8fr1has   (apng_vbetdgo_5t3dis), 

    .o9vvv_q4ikz_2yp0w    (wgcdhfocgyd9bovps), 
    .c1ilkc2r6es72c5h2vcc    (bpgjhz125ozfoh_yq_cze),
    .l3sefagtx4ai4ljb     (d7w4y25gmfw83aoc9 ),
    .josyt39cvr3gignopao     (ppz9xrdau3m7w60f ),
    .bjn5x3u7v4u3rm6d      (zonryv578qcpvne  ), 

    .ipq0f4_yvmml7o06891    (cuzanreq1u8ev47iova), 
    .p4jgl36nmqe8ud7_g4i7    (pg0v_24f5gtcbo20w),
    .wyhg5n7dklr59dxgm_bs     (vuy4dkld2kpsy45c ),
    .ubk6j4rwgfrf5ryn1ibp     (kbqrg_4bxmxn7b7up8 ),
    .cbr_upfu_0ywren54f      (mj86rmgsgeu75euwgxk2  ), 



    .ll0_hbknv5bc_8mxvx5c    (qcz2i1lzeluodju99g0), 
    .qloskxsiztazdeq2ad95i    (vruj1aci16ru7rc5dr),
    .px17v86p_7_1fdvm1w     (t4z031uv53p1rqo1lm9 ),
    .jb9locwfccqzb06jjon     (mazfnbz00ya1f7wlojtz ),
    .a3g162j6o30b4qdpd_z      (fuhx6ea_0i4biqppt  ), 

    .p1jdw9loxkz60taq_vkp_3   (p1jdw9loxkz60taq_vkp_3 ), 
    .ar7xgugq1a_pz7b82ds   (ar7xgugq1a_pz7b82ds ),
    .jwwku_el5h5h2lx6e0kyi    (jwwku_el5h5h2lx6e0kyi  ),
    .vjhpkmep8g_u_cizhsw   (vjhpkmep8g_u_cizhsw ),
    .v19st7vd9_bi485e6ak0   (v19st7vd9_bi485e6ak0 ),
    .zt19omidnr_zyp2gc3bywfb   (zt19omidnr_zyp2gc3bywfb ),
    .gccap1c6hft7o1z7esm     (gccap1c6hft7o1z7esm   ), 
    .eo5skx1ygvzuasbjgnyl    (eo5skx1ygvzuasbjgnyl  ), 

    .pbtolkl953sk14id0iy   (pbtolkl953sk14id0iy  ),
    .z2qyay491938ppnlxuc   (z2qyay491938ppnlxuc  ),
    .zeseql2htbxpugyu5_j      (zeseql2htbxpugyu5_j     ),
    .al3t866kz4po45vfuyjy      (al3t866kz4po45vfuyjy     ),
    .xutsaulafh4onxtthm8n  (xutsaulafh4onxtthm8n ),
    .me7unt7fapqqhtc6epso  (me7unt7fapqqhtc6epso ),
    .m2as3qe7miuhj662j1zvt (m2as3qe7miuhj662j1zvt),



    .xd2ftroj1i79g4derw(czyvvnzs3y3orktdmdfec8yla_1y),
    .qoxd9f57dl083f6cm (o_tztjh1zql5hzdma85okucmgxh ), 



    .gf33atgy                 (gf33atgy          ),
    .ru_wi               (ru_wi        ) 
  );


endmodule                                      














































module vnidphqictr3gtptdwbgr(

  
  
  
  
  input  bwvpn4pm5q2m2, 
  output e79c5kbq9c5f, 

  input  [64-1:0] loc9a4t09i4,
  input  [64-1:0] k2jxyry72hc9nl,
  input  [64-1:0] xtlt33xlczy37q,
  input  [19-1:0] uzxs4linfwcrjy,
  input  [4-1:0] t86na4x45h4ficw,

  output ah6dvj4hwj480v,

  
  
  
  output i_swuedh0b3s, 
  input  qvhs4kakyng1sk, 



  
  
  output baeb5atyeipjmjtwdx66m, 
  input  zf3zgw37xlcc2o5eprc5k, 
  output [64-1:0] a9rvmf7a9nbie6nd923,
  output gzyfsm1lj5vk008,   
  output [4-1:0] w6xoq8do9qo8kitx8e,
  


  input  gf33atgy,
  input  ru_wi
  );

  wire opddptxe1    = uzxs4linfwcrjy[5:5   ];
  wire rm85kx   = uzxs4linfwcrjy[6:6  ];
  wire xt2jzmuzqs = uzxs4linfwcrjy[7:7];
  wire w_wyjws0ma  = uzxs4linfwcrjy[8:8 ];
  wire bu2stjoruwb   = uzxs4linfwcrjy[14:14  ];

          
  
  
  wire tehfiaojgjrpfp_3 = (w_wyjws0ma)            ? 1'b0 : loc9a4t09i4[64-1];
  wire jxdck9cps1z8 = (xt2jzmuzqs | w_wyjws0ma) ? 1'b0 : k2jxyry72hc9nl[64-1];
  wire [64:0] uuxezgs = 
                        {tehfiaojgjrpfp_3, loc9a4t09i4};
  wire [64:0] ajmvhu65z = 
                        {jxdck9cps1z8, k2jxyry72hc9nl};
  
  
  

  
  assign gzyfsm1lj5vk008 = 1'b0;

  
  assign ah6dvj4hwj480v = 1'b0;

  
  
  
  
  
  
  
  
  
  
  
  






  
    wire [2:0] adtau ={ajmvhu65z[1:0],1'b0};
    wire [2:0] f49g58 = ajmvhu65z[3:1];
    wire [2:0] rhgpt = ajmvhu65z[5:3];
    wire [2:0] ollg7 = ajmvhu65z[7:5];
    wire [2:0] xw = ajmvhu65z[9:7];
    wire [2:0] qfmfb5 = ajmvhu65z[11:9];
    wire [2:0] q1z9nzm = ajmvhu65z[13:11];
    wire [2:0] cf6_ = ajmvhu65z[15:13];
    wire [2:0] zq5iq = ajmvhu65z[17:15];
    wire [2:0] ksc = ajmvhu65z[19:17];
    wire [2:0] llw = ajmvhu65z[21:19];
    wire [2:0] hcm2g84 = ajmvhu65z[23:21];
    wire [2:0] rsq0n = ajmvhu65z[25:23];
    wire [2:0] gdrdah = ajmvhu65z[27:25];
    wire [2:0] ys7m = ajmvhu65z[29:27];
    wire [2:0] aa8b73lt = ajmvhu65z[31:29];
    wire [2:0] kzib = ajmvhu65z[33:31];
    wire [2:0] mbigdy = ajmvhu65z[35:33];
    wire [2:0] lf_yup = ajmvhu65z[37:35];
    wire [2:0] j2tdf6cz = ajmvhu65z[39:37];
    wire [2:0] si7g9wy1 = ajmvhu65z[41:39];
    wire [2:0] afy6p = ajmvhu65z[43:41];
    wire [2:0] p6aa8 = ajmvhu65z[45:43];
    wire [2:0] cj9rozp4 = ajmvhu65z[47:45];
    wire [2:0] a4c = ajmvhu65z[49:47];
    wire [2:0] uno = ajmvhu65z[51:49];
    wire [2:0] g904q85c = ajmvhu65z[53:51];
    wire [2:0] egvo = ajmvhu65z[55:53];
    wire [2:0] rk8z = ajmvhu65z[57:55];
    wire [2:0] y3voy9l = ajmvhu65z[59:57];
    wire [2:0] c_sbw3x9 = ajmvhu65z[61:59];
    wire [2:0] kut = ajmvhu65z[63:61];
    wire [2:0] vh6vv44u ={ajmvhu65z[64],ajmvhu65z[64:63]};

    wire [65:0] uhou4275;
    wire [65:0] so6;
    wire [65:0] r28ro5n;
    wire [65:0] wn19654e;
    wire [65:0] ujn4hcqy;
    wire [65:0] bk3frbro;
    wire [65:0] kvm58ey6;
    wire [65:0] m7wg3wdw;
    wire [65:0] gvdlb;
    wire [65:0] j6qw;
    wire [65:0] de2yw;
    wire [65:0] lqr6n54ds;
    wire [65:0] flkp4gvn4;
    wire [65:0] aa4a26a;
    wire [65:0] w_2qgra2;
    wire [65:0] sdxfgz;
    wire [65:0] ski6a;
    wire [65:0] n0rxyxxr;
    wire [65:0] ho9l9u21;
    wire [65:0] zuqqb4;
    wire [65:0] snpg9b;
    wire [65:0] y_6xawz;
    wire [65:0] gsm_x9kx;
    wire [65:0] vksr23hyn;
    wire [65:0] o7myx;
    wire [65:0] odvgzr;
    wire [65:0] i2eoxni0c;
    wire [65:0] u4s5xf2f;
    wire [65:0] tr8s9f;
    wire [65:0] rb1s7rjun;
    wire [65:0] t9xi9g;
    wire [65:0] z4ivp;
    wire [65:0] mhyyf;

    wire [32:0] lit3d5utbsdp3j;


    sneku_08a9mn2xq1ql88_9w6 #(65) e58jpvxqu0kk9u32rpl(.x(adtau), .y(uuxezgs), .iyeq5(uhou4275), .ugjvcvd2l_(lit3d5utbsdp3j[0]));
    sneku_08a9mn2xq1ql88_9w6 #(65) d6_tcp0iskkm_4k8k50_ry(.x(f49g58), .y(uuxezgs), .iyeq5(so6), .ugjvcvd2l_(lit3d5utbsdp3j[1]));
    sneku_08a9mn2xq1ql88_9w6 #(65) m8k9q9gcxlymou7lqq(.x(rhgpt), .y(uuxezgs), .iyeq5(r28ro5n), .ugjvcvd2l_(lit3d5utbsdp3j[2]));
    sneku_08a9mn2xq1ql88_9w6 #(65) syszuxfv6yh7vq66w5d(.x(ollg7), .y(uuxezgs), .iyeq5(wn19654e), .ugjvcvd2l_(lit3d5utbsdp3j[3]));
    sneku_08a9mn2xq1ql88_9w6 #(65) byh9gd6rwzs33_jv73(.x(xw), .y(uuxezgs), .iyeq5(ujn4hcqy), .ugjvcvd2l_(lit3d5utbsdp3j[4]));
    sneku_08a9mn2xq1ql88_9w6 #(65) lyleih1mgwr2qur7qu7wh6(.x(qfmfb5), .y(uuxezgs), .iyeq5(bk3frbro), .ugjvcvd2l_(lit3d5utbsdp3j[5]));
    sneku_08a9mn2xq1ql88_9w6 #(65) jvgf9r0n4vqufegzv(.x(q1z9nzm), .y(uuxezgs), .iyeq5(kvm58ey6), .ugjvcvd2l_(lit3d5utbsdp3j[6]));
    sneku_08a9mn2xq1ql88_9w6 #(65) k7rhcug2ddfzpmvnct5(.x(cf6_), .y(uuxezgs), .iyeq5(m7wg3wdw), .ugjvcvd2l_(lit3d5utbsdp3j[7]));
    sneku_08a9mn2xq1ql88_9w6 #(65) bdwuap8ckn5wsjvioyf65(.x(zq5iq), .y(uuxezgs), .iyeq5(gvdlb), .ugjvcvd2l_(lit3d5utbsdp3j[8]));
    sneku_08a9mn2xq1ql88_9w6 #(65) zw3_o4opyxmw6jb5fx7(.x(ksc), .y(uuxezgs), .iyeq5(j6qw), .ugjvcvd2l_(lit3d5utbsdp3j[9]));
    sneku_08a9mn2xq1ql88_9w6 #(65) vego3pvr7mjmlbb_znega(.x(llw), .y(uuxezgs), .iyeq5(de2yw), .ugjvcvd2l_(lit3d5utbsdp3j[10]));
    sneku_08a9mn2xq1ql88_9w6 #(65) ral_rgv5g17f4c_fu1(.x(hcm2g84), .y(uuxezgs), .iyeq5(lqr6n54ds), .ugjvcvd2l_(lit3d5utbsdp3j[11]));
    sneku_08a9mn2xq1ql88_9w6 #(65) fhlg2fx_64t2x9q29zlfo(.x(rsq0n), .y(uuxezgs), .iyeq5(flkp4gvn4), .ugjvcvd2l_(lit3d5utbsdp3j[12]));
    sneku_08a9mn2xq1ql88_9w6 #(65) zej7_jv9af2sahk9nq2y8tk(.x(gdrdah), .y(uuxezgs), .iyeq5(aa4a26a), .ugjvcvd2l_(lit3d5utbsdp3j[13]));
    sneku_08a9mn2xq1ql88_9w6 #(65) gxcgtfmgrte2p9krl_(.x(ys7m), .y(uuxezgs), .iyeq5(w_2qgra2), .ugjvcvd2l_(lit3d5utbsdp3j[14]));
    sneku_08a9mn2xq1ql88_9w6 #(65) uoakmrlbtd171bu7n_(.x(aa8b73lt), .y(uuxezgs), .iyeq5(sdxfgz), .ugjvcvd2l_(lit3d5utbsdp3j[15]));
    sneku_08a9mn2xq1ql88_9w6 #(65) l55iu_cp84v6lqj7ctfbk(.x(kzib), .y(uuxezgs), .iyeq5(ski6a), .ugjvcvd2l_(lit3d5utbsdp3j[16]));
    sneku_08a9mn2xq1ql88_9w6 #(65) gsyymdli_05eb6v9ty(.x(mbigdy), .y(uuxezgs), .iyeq5(n0rxyxxr), .ugjvcvd2l_(lit3d5utbsdp3j[17]));
    sneku_08a9mn2xq1ql88_9w6 #(65) lb33cboqbahew6zjpt(.x(lf_yup), .y(uuxezgs), .iyeq5(ho9l9u21), .ugjvcvd2l_(lit3d5utbsdp3j[18]));
    sneku_08a9mn2xq1ql88_9w6 #(65) fzkg41m4mpm5tb0a9ghmv(.x(j2tdf6cz), .y(uuxezgs), .iyeq5(zuqqb4), .ugjvcvd2l_(lit3d5utbsdp3j[19]));
    sneku_08a9mn2xq1ql88_9w6 #(65) lpenzlq8yk_fzi81hr6t(.x(si7g9wy1), .y(uuxezgs), .iyeq5(snpg9b), .ugjvcvd2l_(lit3d5utbsdp3j[20]));
    sneku_08a9mn2xq1ql88_9w6 #(65) vpx0k6k006t22_vvkrorxt2(.x(afy6p), .y(uuxezgs), .iyeq5(y_6xawz), .ugjvcvd2l_(lit3d5utbsdp3j[21]));
    sneku_08a9mn2xq1ql88_9w6 #(65) x84u2zqpsk9tmt21d6wk(.x(p6aa8), .y(uuxezgs), .iyeq5(gsm_x9kx), .ugjvcvd2l_(lit3d5utbsdp3j[22]));
    sneku_08a9mn2xq1ql88_9w6 #(65) rhp737jtvnseui1zhn8x(.x(cj9rozp4), .y(uuxezgs), .iyeq5(vksr23hyn), .ugjvcvd2l_(lit3d5utbsdp3j[23]));
    sneku_08a9mn2xq1ql88_9w6 #(65) m08qxjo4aocbvjthog(.x(a4c), .y(uuxezgs), .iyeq5(o7myx), .ugjvcvd2l_(lit3d5utbsdp3j[24]));
    sneku_08a9mn2xq1ql88_9w6 #(65) teqycch9pc9cogqr8zgv7(.x(uno), .y(uuxezgs), .iyeq5(odvgzr), .ugjvcvd2l_(lit3d5utbsdp3j[25]));
    sneku_08a9mn2xq1ql88_9w6 #(65) eo7gou3wc1v2xh1059(.x(g904q85c), .y(uuxezgs), .iyeq5(i2eoxni0c), .ugjvcvd2l_(lit3d5utbsdp3j[26]));
    sneku_08a9mn2xq1ql88_9w6 #(65) ous5ov0eacow957uq9p73we(.x(egvo), .y(uuxezgs), .iyeq5(u4s5xf2f), .ugjvcvd2l_(lit3d5utbsdp3j[27]));
    sneku_08a9mn2xq1ql88_9w6 #(65) tpsw99c3emvib01f38pw(.x(rk8z), .y(uuxezgs), .iyeq5(tr8s9f), .ugjvcvd2l_(lit3d5utbsdp3j[28]));
    sneku_08a9mn2xq1ql88_9w6 #(65) wli6tw5y_d_zo3k9473_6vn(.x(y3voy9l), .y(uuxezgs), .iyeq5(rb1s7rjun), .ugjvcvd2l_(lit3d5utbsdp3j[29]));
    sneku_08a9mn2xq1ql88_9w6 #(65) jflpq4r00ftlk0ve4es(.x(c_sbw3x9), .y(uuxezgs), .iyeq5(t9xi9g), .ugjvcvd2l_(lit3d5utbsdp3j[30]));
    sneku_08a9mn2xq1ql88_9w6 #(65) dswbsd1sq26p0d6ufwwi7x(.x(kut), .y(uuxezgs), .iyeq5(z4ivp), .ugjvcvd2l_(lit3d5utbsdp3j[31]));
    sneku_08a9mn2xq1ql88_9w6 #(65) dgpa9zk_papsg0wxp3ocf(.x(vh6vv44u), .y(uuxezgs), .iyeq5(mhyyf), .ugjvcvd2l_(lit3d5utbsdp3j[32]));




    wire [72:0] artseaok2bnfqwpe1nu2s0 = {{7{uhou4275[65]}},uhou4275}      ;
    wire [72:0] bogyj9x3h4yf8db1pv2te = {{5{so6[65]}},so6,1'b0,lit3d5utbsdp3j[0]} ;
    wire [72:0] l7xt4f3ihc86nn75xya_4 = {{3{r28ro5n[65]}},r28ro5n,1'b0,lit3d5utbsdp3j[1],2'b0} ;
    wire [72:0] aw1hm_tzj_htzy2ocwl0c1 = {wn19654e[65],wn19654e,1'b0,lit3d5utbsdp3j[2],4'b0}      ;
    wire [72:0] b0mo4gs12av2s7rwyv;
    wire [72:0] a1idx6s5tyjkkhg7wtdnd0e;



    mm88fxnds62ofbh80 #(73) v88bm9jhfx6l9ajqjp2( 
                                            .frgfco(artseaok2bnfqwpe1nu2s0),
                                            .ii(bogyj9x3h4yf8db1pv2te),
                                            .fij51v(l7xt4f3ihc86nn75xya_4),
                                            .cuzhl9(aw1hm_tzj_htzy2ocwl0c1),
                                            .c (b0mo4gs12av2s7rwyv),
                                            .s (a1idx6s5tyjkkhg7wtdnd0e)
                                            );


    wire [74:0] vv9yhc5u7uflv9en_eml0f = {{7{ujn4hcqy[65]}},ujn4hcqy,1'b0,lit3d5utbsdp3j[3]}      ;
    wire [74:0] v0eck3vsxjz_wothijmjuirg = {{5{bk3frbro[65]}},bk3frbro,1'b0,lit3d5utbsdp3j[4],2'b0} ;
    wire [74:0] k2o9gmrco6jh5af84h6l1fby = {{3{kvm58ey6[65]}},kvm58ey6,1'b0,lit3d5utbsdp3j[5],4'b0} ;
    wire [74:0] xha1rgvfmkdf2yhmqpb7 = {m7wg3wdw[65],m7wg3wdw,1'b0,lit3d5utbsdp3j[6],6'b0}      ;
    wire [74:0] tuh_9eul1k6smbwhh_rbxg;
    wire [74:0] dy3xtimz9e6_hzbnuu1rk;
    wire [74:0] l_jt4wq5z723fg_93uh5a99du = {{7{gvdlb[65]}},gvdlb,1'b0,lit3d5utbsdp3j[7]}      ;
    wire [74:0] oysbgf5usuf7t8amildgu = {{5{j6qw[65]}},j6qw,1'b0,lit3d5utbsdp3j[8],2'b0} ;
    wire [74:0] i4h_vig7m_4cz8uptt24gmil3 = {{3{de2yw[65]}},de2yw,1'b0,lit3d5utbsdp3j[9],4'b0} ;
    wire [74:0] fj4rz9lp13qngi1wm4wm = {lqr6n54ds[65],lqr6n54ds,1'b0,lit3d5utbsdp3j[10],6'b0}      ;
    wire [74:0] gmwwb1oy9iuj9ksid24o_8bk;
    wire [74:0] rgfjcrpkp7kldkm752d4ti1;
    wire [74:0] qprncc5t6t7cedz428_2ru2ep = {{7{flkp4gvn4[65]}},flkp4gvn4,1'b0,lit3d5utbsdp3j[11]}      ;
    wire [74:0] ex4n9ov6sh9eu5isjcdwqb11lg = {{5{aa4a26a[65]}},aa4a26a,1'b0,lit3d5utbsdp3j[12],2'b0} ;
    wire [74:0] wbehy1mlinq6mmeop_mhj2805w = {{3{w_2qgra2[65]}},w_2qgra2,1'b0,lit3d5utbsdp3j[13],4'b0} ;
    wire [74:0] fubh867zwdatmf4vcdg7t7ex7 = {sdxfgz[65],sdxfgz,1'b0,lit3d5utbsdp3j[14],6'b0}      ;
    wire [74:0] wwp3992ul88cguj4nzkb5eu;
    wire [74:0] jhq8kol0mc7qgwbrxamz;
    wire [74:0] aroan00ywfn4mbk2wgu438f5u = {{7{ski6a[65]}},ski6a,1'b0,lit3d5utbsdp3j[15]}      ;
    wire [74:0] lmc13yfnhtkd88ng6vg25dq = {{5{n0rxyxxr[65]}},n0rxyxxr,1'b0,lit3d5utbsdp3j[16],2'b0} ;
    wire [74:0] zarhesuwa8rzfrdb1rjpr_kevp = {{3{ho9l9u21[65]}},ho9l9u21,1'b0,lit3d5utbsdp3j[17],4'b0} ;
    wire [74:0] mosd6jwym_rjlij4gu_xu47 = {zuqqb4[65],zuqqb4,1'b0,lit3d5utbsdp3j[18],6'b0}      ;
    wire [74:0] cog31c8vbugu6ll4xcqdxxmnp;
    wire [74:0] whrlys_hu8bedrjn3i03hvk;
    wire [74:0] zftvswl45hkmm09dmmuwken = {{7{snpg9b[65]}},snpg9b,1'b0,lit3d5utbsdp3j[19]}      ;
    wire [74:0] ftehnvh5_7c5e1ms9d70dcu = {{5{y_6xawz[65]}},y_6xawz,1'b0,lit3d5utbsdp3j[20],2'b0} ;
    wire [74:0] wfqhmju69ql45bm1mqlh9 = {{3{gsm_x9kx[65]}},gsm_x9kx,1'b0,lit3d5utbsdp3j[21],4'b0} ;
    wire [74:0] w19xw0yb9ti4kwb2k_nltwz8 = {vksr23hyn[65],vksr23hyn,1'b0,lit3d5utbsdp3j[22],6'b0}      ;
    wire [74:0] tiyhmxq22wuwlcs7nbsvr;
    wire [74:0] o8oyg3oy5vqfs5znl0wvf1a1v;
    wire [74:0] oes8dinyxo993z_24jinv = {{7{o7myx[65]}},o7myx,1'b0,lit3d5utbsdp3j[23]}      ;
    wire [74:0] j3w01y5tbh7hqth9l86wf77hp = {{5{odvgzr[65]}},odvgzr,1'b0,lit3d5utbsdp3j[24],2'b0} ;
    wire [74:0] yv8kdk6y63u_tpaxnprrzcgi6r = {{3{i2eoxni0c[65]}},i2eoxni0c,1'b0,lit3d5utbsdp3j[25],4'b0} ;
    wire [74:0] iuqbg94t5907efuons8s00 = {u4s5xf2f[65],u4s5xf2f,1'b0,lit3d5utbsdp3j[26],6'b0}      ;
    wire [74:0] hqhnq414f4jzb0fwgb6r75e8;
    wire [74:0] ko9ada4o4fzcrfgxynewslr;
    wire [74:0] x_nvsu_6a565nja94h9e0ust4 = {{7{tr8s9f[65]}},tr8s9f,1'b0,lit3d5utbsdp3j[27]}      ;
    wire [74:0] bhiv7dibelh14du6_51l165 = {{5{rb1s7rjun[65]}},rb1s7rjun,1'b0,lit3d5utbsdp3j[28],2'b0} ;
    wire [74:0] ut9dukgypfd0ttlw6qz6z5 = {{3{t9xi9g[65]}},t9xi9g,1'b0,lit3d5utbsdp3j[29],4'b0} ;
    wire [74:0] g18slisntfvg8r52921qtqv = {z4ivp[65],z4ivp,1'b0,lit3d5utbsdp3j[30],6'b0}      ;
    wire [74:0] x9j2dvl4azif8cf7hreff;
    wire [74:0] nzhrp3j69rcvgvs2fd5f4xfm7;



    mm88fxnds62ofbh80 #(75) vqcbz4sb8i45a5vx( 
                                            .frgfco(vv9yhc5u7uflv9en_eml0f),
                                            .ii(v0eck3vsxjz_wothijmjuirg),
                                            .fij51v(k2o9gmrco6jh5af84h6l1fby),
                                            .cuzhl9(xha1rgvfmkdf2yhmqpb7),
                                            .c (tuh_9eul1k6smbwhh_rbxg),
                                            .s (dy3xtimz9e6_hzbnuu1rk)
                                            );

    mm88fxnds62ofbh80 #(75) ql_mzujlocx22g731( 
                                            .frgfco(l_jt4wq5z723fg_93uh5a99du),
                                            .ii(oysbgf5usuf7t8amildgu),
                                            .fij51v(i4h_vig7m_4cz8uptt24gmil3),
                                            .cuzhl9(fj4rz9lp13qngi1wm4wm),
                                            .c (gmwwb1oy9iuj9ksid24o_8bk),
                                            .s (rgfjcrpkp7kldkm752d4ti1)
                                            );

    mm88fxnds62ofbh80 #(75) aa5zhqctw02eowglai61xud( 
                                            .frgfco(qprncc5t6t7cedz428_2ru2ep),
                                            .ii(ex4n9ov6sh9eu5isjcdwqb11lg),
                                            .fij51v(wbehy1mlinq6mmeop_mhj2805w),
                                            .cuzhl9(fubh867zwdatmf4vcdg7t7ex7),
                                            .c (wwp3992ul88cguj4nzkb5eu),
                                            .s (jhq8kol0mc7qgwbrxamz)
                                            );

    mm88fxnds62ofbh80 #(75) xrdl77vy1ipordwf70t2d( 
                                            .frgfco(aroan00ywfn4mbk2wgu438f5u),
                                            .ii(lmc13yfnhtkd88ng6vg25dq),
                                            .fij51v(zarhesuwa8rzfrdb1rjpr_kevp),
                                            .cuzhl9(mosd6jwym_rjlij4gu_xu47),
                                            .c (cog31c8vbugu6ll4xcqdxxmnp),
                                            .s (whrlys_hu8bedrjn3i03hvk)
                                            );

    mm88fxnds62ofbh80 #(75) ku7rgyql9d7tjz2rhfac( 
                                            .frgfco(zftvswl45hkmm09dmmuwken),
                                            .ii(ftehnvh5_7c5e1ms9d70dcu),
                                            .fij51v(wfqhmju69ql45bm1mqlh9),
                                            .cuzhl9(w19xw0yb9ti4kwb2k_nltwz8),
                                            .c (tiyhmxq22wuwlcs7nbsvr),
                                            .s (o8oyg3oy5vqfs5znl0wvf1a1v)
                                            );

    mm88fxnds62ofbh80 #(75) bx07iwm4hk47m1th5ukm( 
                                            .frgfco(oes8dinyxo993z_24jinv),
                                            .ii(j3w01y5tbh7hqth9l86wf77hp),
                                            .fij51v(yv8kdk6y63u_tpaxnprrzcgi6r),
                                            .cuzhl9(iuqbg94t5907efuons8s00),
                                            .c (hqhnq414f4jzb0fwgb6r75e8),
                                            .s (ko9ada4o4fzcrfgxynewslr)
                                            );

    mm88fxnds62ofbh80 #(75) kg22c62yfsw7qr4r6bann( 
                                            .frgfco(x_nvsu_6a565nja94h9e0ust4),
                                            .ii(bhiv7dibelh14du6_51l165),
                                            .fij51v(ut9dukgypfd0ttlw6qz6z5),
                                            .cuzhl9(g18slisntfvg8r52921qtqv),
                                            .c (x9j2dvl4azif8cf7hreff),
                                            .s (nzhrp3j69rcvgvs2fd5f4xfm7)
                                            );



    wire [81:0] qo_2neg6_gtug5n9q8kc = {{9{b0mo4gs12av2s7rwyv[72]}},b0mo4gs12av2s7rwyv}    ;
    wire [81:0] nv500uy_zrnl5dm4o3hq51j = {{9{a1idx6s5tyjkkhg7wtdnd0e[72]}},a1idx6s5tyjkkhg7wtdnd0e}    ;
    wire [81:0] j4yj5bjku_wvfy9m5x_ = {tuh_9eul1k6smbwhh_rbxg[74],tuh_9eul1k6smbwhh_rbxg,6'b0}  ;
    wire [81:0] d0htfqflvcnbx7bc_omv = {dy3xtimz9e6_hzbnuu1rk[74],dy3xtimz9e6_hzbnuu1rk,6'b0}  ;
    wire [81:0] lowiib1xy2c5vjzu652;
    wire [81:0] rjjzv5dt85m56wfinhltab;




    mm88fxnds62ofbh80 #(82) cgd4_uposvz_ybm2(
                                            .frgfco(qo_2neg6_gtug5n9q8kc),
                                            .ii(nv500uy_zrnl5dm4o3hq51j),
                                            .fij51v(j4yj5bjku_wvfy9m5x_),
                                            .cuzhl9(d0htfqflvcnbx7bc_omv),
                                            .c (lowiib1xy2c5vjzu652),
                                            .s (rjjzv5dt85m56wfinhltab)
                                            );





    wire [83:0] vwdxukzfhex2s_3rbcya4oaw = {{9{gmwwb1oy9iuj9ksid24o_8bk[74]}},gmwwb1oy9iuj9ksid24o_8bk}    ;
    wire [83:0] o0sc58hn5h05ldlgxwsxl1r3 = {{9{rgfjcrpkp7kldkm752d4ti1[74]}},rgfjcrpkp7kldkm752d4ti1}    ;
    wire [83:0] wuo00f94qhxx_xnbjf8axtj3 = {wwp3992ul88cguj4nzkb5eu[74],wwp3992ul88cguj4nzkb5eu,8'b0}  ;
    wire [83:0] vt_yoz_9gnj0qye_r45mf = {jhq8kol0mc7qgwbrxamz[74],jhq8kol0mc7qgwbrxamz,8'b0}  ;
    wire [83:0] reryysqv5uk8acg9tu_coses;
    wire [83:0] uqe_xa0mbvlcuhgw8t3hlmo;

    wire [83:0] zn2s_h6vhecr0bjvaarc4qms = {{9{cog31c8vbugu6ll4xcqdxxmnp[74]}},cog31c8vbugu6ll4xcqdxxmnp}    ;
    wire [83:0] cscgi3k5_aops7m_a0p_t = {{9{whrlys_hu8bedrjn3i03hvk[74]}},whrlys_hu8bedrjn3i03hvk}    ;
    wire [83:0] yp9aq9ox3bssrsg8b3g6dlb8 = {tiyhmxq22wuwlcs7nbsvr[74],tiyhmxq22wuwlcs7nbsvr,8'b0}  ;
    wire [83:0] o_mslaup_6wgykcoehb6ck = {o8oyg3oy5vqfs5znl0wvf1a1v[74],o8oyg3oy5vqfs5znl0wvf1a1v,8'b0}  ;
    wire [83:0] tejm0pqk6irgx5wnzb_xizf6k;
    wire [83:0] g7dfsj7xj2o1u66s8xs0n6si;

    wire [83:0] tfyrp8z_m8o5j9lmpot_e = {{9{hqhnq414f4jzb0fwgb6r75e8[74]}},hqhnq414f4jzb0fwgb6r75e8}    ;
    wire [83:0] vd75xxrhbbju_102av1u2 = {{9{ko9ada4o4fzcrfgxynewslr[74]}},ko9ada4o4fzcrfgxynewslr}    ;
    wire [83:0] jjdcpss2a_c54a30b6v6_ = {x9j2dvl4azif8cf7hreff[74],x9j2dvl4azif8cf7hreff,8'b0}  ;
    wire [83:0] r4kij6cuslp43loqddyqv8l = {nzhrp3j69rcvgvs2fd5f4xfm7[74],nzhrp3j69rcvgvs2fd5f4xfm7,8'b0}  ;
    wire [83:0] d7khfpdzothcf4ws20m1q;
    wire [83:0] j03byb664ak5qx4lmj6fnwf;




    mm88fxnds62ofbh80 #(84) ciu340o76n0mi6tnduv(
                                            .frgfco(vwdxukzfhex2s_3rbcya4oaw),
                                            .ii(o0sc58hn5h05ldlgxwsxl1r3),
                                            .fij51v(wuo00f94qhxx_xnbjf8axtj3),
                                            .cuzhl9(vt_yoz_9gnj0qye_r45mf),
                                            .c (reryysqv5uk8acg9tu_coses),
                                            .s (uqe_xa0mbvlcuhgw8t3hlmo)
                                            );



    mm88fxnds62ofbh80 #(84) z4b9shs6yv2ztpi2s68yv(
                                            .frgfco(zn2s_h6vhecr0bjvaarc4qms),
                                            .ii(cscgi3k5_aops7m_a0p_t),
                                            .fij51v(yp9aq9ox3bssrsg8b3g6dlb8),
                                            .cuzhl9(o_mslaup_6wgykcoehb6ck),
                                            .c (tejm0pqk6irgx5wnzb_xizf6k),
                                            .s (g7dfsj7xj2o1u66s8xs0n6si)
                                            );



    mm88fxnds62ofbh80 #(84) i2c21sw5v29urvz27t(
                                            .frgfco(tfyrp8z_m8o5j9lmpot_e),
                                            .ii(vd75xxrhbbju_102av1u2),
                                            .fij51v(jjdcpss2a_c54a30b6v6_),
                                            .cuzhl9(r4kij6cuslp43loqddyqv8l),
                                            .c (d7khfpdzothcf4ws20m1q),
                                            .s (j03byb664ak5qx4lmj6fnwf)
                                            );





    wire [98:0] dobz8mu1bx05if98iwxcbuii = {{17{lowiib1xy2c5vjzu652[81]}},lowiib1xy2c5vjzu652}   ;
    wire [98:0] ir4_disya8tp3mnqny4ge8mrb = {{17{rjjzv5dt85m56wfinhltab[81]}},rjjzv5dt85m56wfinhltab}   ;
    wire [98:0] q0a4irzufgr1i6h7xxstk0t = {reryysqv5uk8acg9tu_coses[83],reryysqv5uk8acg9tu_coses,14'b0} ;
    wire [98:0] v5o_eh92bqax8hw2nrism_o = {uqe_xa0mbvlcuhgw8t3hlmo[83],uqe_xa0mbvlcuhgw8t3hlmo,14'b0} ;
    wire [98:0] j979ctfnafqdzi10al133dcr;
    wire [98:0] q0orucfbnv92bvtgbi7;

    mm88fxnds62ofbh80 #(99) wwdj_pcz6za60lmlkj03l(
                                            .frgfco(dobz8mu1bx05if98iwxcbuii),
                                            .ii(ir4_disya8tp3mnqny4ge8mrb),
                                            .fij51v(q0a4irzufgr1i6h7xxstk0t),
                                            .cuzhl9(v5o_eh92bqax8hw2nrism_o),
                                            .c (j979ctfnafqdzi10al133dcr),
                                            .s (q0orucfbnv92bvtgbi7)
                                            );






    wire [100:0] ry7mv5r6r7decfuil1nvpddt6e = {{17{tejm0pqk6irgx5wnzb_xizf6k[83]}},tejm0pqk6irgx5wnzb_xizf6k}   ;
    wire [100:0] d92msahalq4xn211c5ld0tyq = {{17{g7dfsj7xj2o1u66s8xs0n6si[83]}},g7dfsj7xj2o1u66s8xs0n6si}   ;
    wire [100:0] ag8ycz6qg28vupccjabu4w1j3_ = {d7khfpdzothcf4ws20m1q[83],d7khfpdzothcf4ws20m1q,16'b0} ;
    wire [100:0] ifpofwz9u_w8om9vptvi6pf = {j03byb664ak5qx4lmj6fnwf[83],j03byb664ak5qx4lmj6fnwf,16'b0} ;
    wire [100:0] z6_frvzvzlu2901frkti4;
    wire [100:0] njxr0sukghngyiyis1_zy;

    mm88fxnds62ofbh80 #(101) l5o3wla5mq826jadk0t(
                                            .frgfco(ry7mv5r6r7decfuil1nvpddt6e),
                                            .ii(d92msahalq4xn211c5ld0tyq),
                                            .fij51v(ag8ycz6qg28vupccjabu4w1j3_),
                                            .cuzhl9(ifpofwz9u_w8om9vptvi6pf),
                                            .c (z6_frvzvzlu2901frkti4),
                                            .s (njxr0sukghngyiyis1_zy)
                                            );








    localparam eix5yfq_9smolgn22c = 99*2 + 101*2 + 66 + 2 + 5 + 4;

    wire [eix5yfq_9smolgn22c-1:0] p2m0vw0_2ox53 ={
                                        j979ctfnafqdzi10al133dcr,
                                        q0orucfbnv92bvtgbi7,
                                        z6_frvzvzlu2901frkti4,
                                        njxr0sukghngyiyis1_zy,
                                        mhyyf,
                                        lit3d5utbsdp3j[31],
                                        lit3d5utbsdp3j[32],
                                        opddptxe1, 
                                        rm85kx, 
                                        xt2jzmuzqs,
                                        w_wyjws0ma,
                                        bu2stjoruwb,
                                        t86na4x45h4ficw
                                        };
    wire [eix5yfq_9smolgn22c-1:0] rhs_t37ij54sv37;
    wire tzul_ch7haingdjl = bwvpn4pm5q2m2 & qvhs4kakyng1sk;
    wire u8tkz3vm0w0bfsaj3b;
    assign  e79c5kbq9c5f = qvhs4kakyng1sk & u8tkz3vm0w0bfsaj3b;
    assign  i_swuedh0b3s = bwvpn4pm5q2m2 & u8tkz3vm0w0bfsaj3b;
    
    wire u43jg7xrb7hnl, s81rsj8wxn777l;
    ux607_gnrl_pipe_stage # (
     .CUT_READY(0),
     .DP(1),
     .DW(eix5yfq_9smolgn22c)
    ) dfgyxcmvfdxo7mplbr (
      .i_vld(tzul_ch7haingdjl), 
      .i_rdy(u8tkz3vm0w0bfsaj3b), 
      .i_dat(p2m0vw0_2ox53 ),
      .o_vld(u43jg7xrb7hnl), 
      .o_rdy(s81rsj8wxn777l), 
      .o_dat(rhs_t37ij54sv37 ),

      .clk  (gf33atgy  ),
      .rst_n(ru_wi)  
     );

    wire f31k2irxac1h, n0ucnwblq5_p9w, fk6u20a6q_a768, cuufn57r8amwl9, lf75xcymewz9;
    wire [4-1:0] vceby3abadx5w3irv13;
    wire [98:0] b_qehkn641cgx7yckmh6pginjbd;
    wire [98:0] ra1m09r1vzetfg91ohotzdhql3ay;
    wire [100:0] zvo8y4p5t0kfttmgj2ss1bqs0o52to;
    wire [100:0] zmed7do3ajqsnse0xayni52l5kv;
    wire [65:0] ahv0qe18zj8a5;
    wire        s5wu2ztotq0n9oqn592zc;
    wire        vg1njuqyid4zobv1qk60c;
    assign {b_qehkn641cgx7yckmh6pginjbd,
            ra1m09r1vzetfg91ohotzdhql3ay,
            zvo8y4p5t0kfttmgj2ss1bqs0o52to,
            zmed7do3ajqsnse0xayni52l5kv,
            ahv0qe18zj8a5,
            s5wu2ztotq0n9oqn592zc,
            vg1njuqyid4zobv1qk60c,
            f31k2irxac1h,
            n0ucnwblq5_p9w,
            fk6u20a6q_a768,
            cuufn57r8amwl9,
            lf75xcymewz9,
            vceby3abadx5w3irv13
            } = rhs_t37ij54sv37;





    wire [131:0] heuc5j0phvwdztm2iw3bcliq = {{33{b_qehkn641cgx7yckmh6pginjbd[98]}},b_qehkn641cgx7yckmh6pginjbd}       ;
    wire [131:0] dh67xqurkx49gyno4s956xi4x = {{33{ra1m09r1vzetfg91ohotzdhql3ay[98]}},ra1m09r1vzetfg91ohotzdhql3ay}       ;
    wire [131:0] rn1q5v0q8f2jh05srf2h = {zvo8y4p5t0kfttmgj2ss1bqs0o52to[100],zvo8y4p5t0kfttmgj2ss1bqs0o52to,30'b0}   ;
    wire [131:0] dv4az7spmixb71lc5yb0udck = {zmed7do3ajqsnse0xayni52l5kv[100],zmed7do3ajqsnse0xayni52l5kv,30'b0}   ;
    wire [131:0] utepmmhq68fopal1qsolvm;
    wire [131:0] oxysblq2yv0mr2f8odruhbpt;

    mm88fxnds62ofbh80 #(132) hh670k73ixx3gw2a9(
                                            .frgfco(heuc5j0phvwdztm2iw3bcliq),
                                            .ii(dh67xqurkx49gyno4s956xi4x),
                                            .fij51v(rn1q5v0q8f2jh05srf2h),
                                            .cuzhl9(dv4az7spmixb71lc5yb0udck),
                                            .c (utepmmhq68fopal1qsolvm),
                                            .s (oxysblq2yv0mr2f8odruhbpt)
                                            );




    
    wire [130:0] nrii3wq28qbjn9u_ymmd40wy = utepmmhq68fopal1qsolvm[130:0];
    wire [130:0] itws_si6qiqjgj1p3rlj9g3a = oxysblq2yv0mr2f8odruhbpt[130:0];
    wire [130:0] qfczfkz30yn2o08mdacuwppy9 = {ahv0qe18zj8a5[65],ahv0qe18zj8a5,1'b0,s5wu2ztotq0n9oqn592zc,62'b0};
    wire [130:0] ep8lfw7qjnjts2_5zttu2vmj = {66'b0, vg1njuqyid4zobv1qk60c,64'b0};
    wire [130:0] b9r9xzkmfg7lr8hlgy7;
    wire [130:0] kxxd16j6b1japw7s0hn5k;

    mm88fxnds62ofbh80 #(131) c0p6xwtv8lvicjcauel2gh(
                                            .frgfco(nrii3wq28qbjn9u_ymmd40wy),
                                            .ii(itws_si6qiqjgj1p3rlj9g3a),
                                            .fij51v(qfczfkz30yn2o08mdacuwppy9),
                                            .cuzhl9(ep8lfw7qjnjts2_5zttu2vmj),
                                            .c (b9r9xzkmfg7lr8hlgy7),
                                            .s (kxxd16j6b1japw7s0hn5k)
                                            );


    localparam sdvetn3bnzz0_hpiyu = 4 * 64 + 5 + 4; 

    wire [sdvetn3bnzz0_hpiyu-1:0] i7r5kurxvcwo42 = { 
                                            b9r9xzkmfg7lr8hlgy7[2*64-1:0], 
                                            kxxd16j6b1japw7s0hn5k[2*64-1:0],
                                            f31k2irxac1h,
                                            n0ucnwblq5_p9w,
                                            fk6u20a6q_a768,
                                            cuufn57r8amwl9,
                                            lf75xcymewz9,
                                            vceby3abadx5w3irv13
                                            };
 
    
    wire [sdvetn3bnzz0_hpiyu-1:0] ixyuzhmi46_8;
    wire avfgzyfbb4mp4y;
    wire sums7_3xypuac33_6o;

    ux607_gnrl_pipe_stage # (
    .CUT_READY(0),
    .DP(0),
    .DW(sdvetn3bnzz0_hpiyu)
    ) mgjo0_fpra_wk_na6 (
        .i_vld(u43jg7xrb7hnl),
        .i_rdy(s81rsj8wxn777l),
        .i_dat(i7r5kurxvcwo42),
        .o_vld(avfgzyfbb4mp4y),
        .o_rdy(sums7_3xypuac33_6o),
        .o_dat(ixyuzhmi46_8),

        .clk   (gf33atgy),
        .rst_n (ru_wi)
    );
    
    wire e7dz9m7fya_a, utio9j3ajijhds, vj3rb70xb6pop_v, kj8c7zaqibye9m;
    wire h5vuk2dh4n;

    wire [4-1:0] vynxjbp4xjqmn4h3ul8;
    wire [2*64-1:0] z_ytubdlq72fq;
    wire [2*64-1:0] j64wathign93n;

    assign {z_ytubdlq72fq,
            j64wathign93n,
            e7dz9m7fya_a,
            utio9j3ajijhds,
            vj3rb70xb6pop_v,
            kj8c7zaqibye9m,
            h5vuk2dh4n,
            vynxjbp4xjqmn4h3ul8
            } = ixyuzhmi46_8;





    wire [2*64-1:0] wrcjvt7pl1j_ = z_ytubdlq72fq[2*64-1:0] + j64wathign93n[2*64-1:0];
    

    wire [64-1:0] k6vc5gb7qcv     = wrcjvt7pl1j_[64-1:0];
    wire [64-1:0] nsraxk6bxkv    = wrcjvt7pl1j_[2*64-1:64];
    wire [64-1:0] x1z_g1j61g  = wrcjvt7pl1j_[2*64-1:64];
    wire [64-1:0] lnvdkfx8skcfm   = wrcjvt7pl1j_[2*64-1:64];
    wire [63:0] ncu6_95gm7ck    = {{32{wrcjvt7pl1j_[31]}},wrcjvt7pl1j_[31:0]};

    assign baeb5atyeipjmjtwdx66m = avfgzyfbb4mp4y;
    assign sums7_3xypuac33_6o = zf3zgw37xlcc2o5eprc5k;
    assign a9rvmf7a9nbie6nd923 = 
           ({64{e7dz9m7fya_a   }} & k6vc5gb7qcv    )
         | ({64{utio9j3ajijhds  }} & nsraxk6bxkv   )
         | ({64{vj3rb70xb6pop_v}} & x1z_g1j61g )
         | ({64{kj8c7zaqibye9m }} & lnvdkfx8skcfm  )
         | ({64{h5vuk2dh4n  }} & ncu6_95gm7ck   )
         ;

    assign w6xoq8do9qo8kitx8e = vynxjbp4xjqmn4h3ul8;








































































endmodule                                      
























































module b0gv4gv3sqckul0vbemwxr #(
 parameter gdctpuyrfi_b        = 0,
 parameter l_7qc0w_2x6i        = 0,
 parameter f6daaph5or1       = 0,
 parameter t5462hhws9i6ynbxi    = 0 
)(

  input [4-1:0]        cu1owrury8wsed,
  input [4-1:0]        mt1z8r_sz,
  input [4-1:0]        uc9k3lw_iehx,
  input [4-1:0]        radwr7skyhm3jqso5,
  input [4-1:0]        zdid44qi3bv7q4phl,
  input [4-1:0]        x4owqbu74zh_xxr,

  input                            b43m7n67rav8he, 
  input                            qcutfgh43gov5u4urt,
  input                            s73raoa0ilom1wyi,
  input                            dnwb40nhmse7rcj0epzjo,
  input                            omeribg0gbgvpn78urilv_a,
  input                            jxogr1vy8jotyh8ivd2u,

  input [64-1:0]           kl8zh4diafqs , 
  input [64-1:0]           jiartjoiycj2 , 
  input [64-1:0]           dtypmpwq1q2j , 
  input                            uwl7jm0d1lv0xpo, 
  input                            u2l80pdclhyu1bl, 
  input                            uamf3ccv7ouhi18,  
  input [64-1:0]           pkw60eo867gghh , 
  input [64-1:0]           strg8286lgex8p4_0m , 
  input [64-1:0]           avpvrch0prpui67 , 


  input                            e7nqb0p7cffw4lrkd  ,


  input                            cvqaktep17ac   ,
  output                           h91pmjbyad1itr37   ,
  input [32-1:0]     nv33gk9s6_      ,
  input [64-1:0]        cyudxl51e      ,
  input [4-1:0]     z8xxe17sssy8tr8q219,
  input [64-1:0]           plk8ixck4wj7c    , 
  input                            u4k7uyzg9lp3zlf  ,
  input                            ej5tfrzf8ad7noezo8gdkb1xg4 ,
  input                            ekmvur7r4qz7ea7htd ,
  input                            ndvqmbwgzq08mbdaxnn4 ,
  input                            dorqi70cvs05s ,
  input                            pgfbjdj832ly_ ,
  input                            z0yti764_a15nwanb , 
  input                            k5yu5na0oo41y  ,
  input                            n8g2a10i7cbowtvjhc  ,
  input                            pzlsmt96uolwfb47  ,
  input [5-1:0]    uzn8ik3rkkwib6p  , 

  input [64-1:0]           kh00jq7wde_slaj , 
  input [64-1:0]           rezwnhzl7vmkg , 
  input [64-1:0]           nq_d1dxi6n86s , 

  input [64-1:0]        rx4zxlit4v_5k4fclu   ,
  input [64-1:0]        k_7iagb48feg9b3wj    ,
  input [4*8-1:0]    lot9xvzuqrd5jm0scdx5t,
  input [7:0]                      mn3tic51ckga0gc,
  input [2:0]                      k0be3wres3xocvs9tpkn4fu,  
  input                            akk0_n8kvb1w0wxrz,
  input                            cnp1c4afdljmpemgot3sa,
  input                            wsh7h1p7b0zifvs0kwabih,
  input                            qhk0gez3kmex8twzly7mxn,
  input [64-1:0]        rafwujb8lw59lcbn9vsz8o,
  input                            dqpwtmmizdh6bvzsx6,
  input                            cuxay1hemfm214cwu1513x,
  input                            s6in6vliinq9udhsofa,
  input [2-1:0]      ephp7dpea6ymyg0eucjv0,
  input [9-1:0]   w42z5c2wv916u4df79p,
  input                            vq3a19my9wldb5hug_nnbu0,

  input                            imj0glh0tzynz,
  input                            mn8sk0gr9oh54zn_o  ,
  input                            oetzq1g528ymdza0maph  ,
  input                            bwsazwvhtn9in7lpyjssdk  ,
  input                            aly0oms0x8r1kmmdgyob ,
  input                            vckb4tc8r10z7n621obxkju ,
  input                            f3lw5s13_0u5q6o4ep ,
  input    [4-1:0]     x11xtpe4e78unv1ahgzinz4n,
  input    [4-1:0]     ialrcyi5grz5o0hc0jyjuwv,
  input    [4-1:0]     wfpum3du8gc8hr_xuerx,

  input                            rtjejhmafpq7db,
  input                            vnc88f08k1s0obtnvb,
  input                            u5pfnkzvz6fsvmgw4,
  input                            zlk2yur1jgjwg,
  input                            ow91ik9ily4bugcc43pp,
  input                                bf8iyrsqp4a2s,
  input                                pu764metopn524rq4hg2c24,
  input [105-1:0]  j7l4qmkctu4k_1q6c,
  input [50-1:0] x6t2ufv1z2uufogo,
  input                              q5_q35rctah_,
  input                              hm3iwty3s1d4si2p4,
  input                              txcys7e9ezk6xikpy2hu987,
  input [48-1:0]    eph11j28sez0oftr7b,  
  input [64-1:0]             lq6932o27hlk9v4f1m,
  input                              sll07sleuwo2fkitj,
  input                              v2e4q5r07qxd6fxruqia3f,
  input                              e5nqx8gg2u3gxy0y4c,
  input                              ajka24wmafrwpta96cf2,
  input                              bod813pzaejozw9p1,

  input                              z1et08p41uxcl76,
  input [48-1:0]    jymdjzitd0hv0e9uhul,  
  input                            pwppbjb8emt8vd9_w,
  input [19-1:0]  z69pfny03ofcxvjyygmo6, 
  input [48-1:0]  juyjh9cdf4vvzhq,

  input                            vh0cb71_xnjsewqur3,
  input                            gbgabhg8e_ul0e24r6jq,
  input                            mtsy6_whdwum2fu   ,
  input                            k_igx5_oeq1ag3m   ,
  input                            th3snuy_v19o06eanj,
  input                            xxggjmznfu9b_    ,
  input  [64-1:0]          t9kvx890cyg     ,
  input  [64-1:0]          i984chc2gxtcivks ,
  input                            w37tf6nz0oty_z89xv1,
  input                            pfeci7n4c83yiwln58,
  input                            mzu7xfmjf4mwa0b ,
  input                            g3t8ql0mi58ddizau_8t3 ,
  input                            gg468ty1pm6_zgec ,
  input                            jtvucg9wp5nxn,
  input                            ofe8xctslv6q5w48ky,
  input                            axbsuznhe7w6rrd   ,
  input                            j49by1lxo4ie9_ho   ,
  input                            tv7ak8mtfqswt    ,
  input                            kr13pzf9ml9ic_vbl    ,
  input                            wkixlev_tj12x_lfp6p04t ,
  input                            jzx45r8bb79aj5ddz7h_565f,


  input                            rgip60bn9st8htirgmhnohyj    ,
  input                            duo6acmepph_0ahl_0ebyyjh  ,
  input                            mylxtynzir7dvcouvb5thi    ,
  input                            o5yttui8un64i2r3s3yxxxjc25iwv  ,

  input                            fxsynukaasxx8lt57bwdodyn3cem  ,
  input                            oel93f4rkl6esczbag9yld       ,
  input                            vmp6zvyj46lrfmg3bl_kecu59    ,
  input                            gj_lc7e2uh1cdx5b2bmynhvw   ,
  input                            b7ker79ak62g5qei_oa7kxdm0   ,
  input  [64-1:0]     i3rcr_tmnynzs9lr254bac9x2b  ,
  input                            ti5a3yv8_m3rzzigzeuzrt1 ,
  input                            cb86_62ddnv8i2whbc   ,

  input                            i_2lk2qupeba0sjgw6sdnbedc,
  input                            a46z1a4rlrucmwj5ju3o83orp8jx2e,
  input                            ti9h9knu4vrm6k3vqry9vfxbc4b,
  input                            p8zi9oi86dxmkaq4uqhu8j1hl0e,
  input                            plmzz80_s0_tb0kwjjgu5p7uktpi2,
  input  [64-1:0]     z_r1pp7wjooqw6n7rnoyv7nka81o,

  output                           akdv8vv97zk549v,   
  input                            k_wnu24cz94zwh8,   
  output [64-1:0]       zpdph1sve,      
  output [32-1:0]    o9d_zhwhmsph,      
  output [4-1:0]       dte0cay394mhjhkr,
  output [64-1:0]          v8zi5h4rj36jt    ,
  output [64-1:0]          livvja2ywo91o8v    ,
  output [64-1:0]          t5p9q190fm    ,

  output [64-1:0]          dckyl_qt92wqvghtw3    ,
  output [64-1:0]          vyug4w9rb9kj6bmwwu    ,
  output [64-1:0]          h40f1u8xaz57o3c    ,
  output [64-1:0]          bv8rdomgcr9w6r2z    ,
  output [64-1:0]          ujgn98iv8k5xidjk    ,

  output [64-1:0]          fw_dplmj46w6    ,
  output                           jdngc81st67hk8p  ,
  output                           u4t194j1c9najq  ,
  output                           gkzjw6iff1idxo   ,
  output [5-1:0]   jcj76rmi3pqujm3v  ,
  output                           ptu54kun7juh0 ,
  output                           tsns5phts_z2fnf ,
  output                           rsdyvyptjiksvewu ,
  output                           pysgbgu5mzucuewf1,   
  output                           g65q46nnz7gip0zyo,
  output                           zf1w750jg2mtdij,   
  output                           pw6i533r0oou6ub,   
  output                           getq71b86zu18ri7x,   
  output                           tp46wehs200pll2qi,   
  output                           iouqv7uynzgvde_v,    
  output                           hb36pq8e0n24raht15 ,
  output                           xphk4z06widyipxfcjr ,
  output                           xcu8n5tos13pfc6jhw22 ,
  output                           lbx9pnfl2z4is68kam,
  output                           hl9x8gmcd9k2ttm0hui2j,
  output                           ioka849821_gx48yl9gk,
  output [4-1:0]       j9fcegru44_r74xlm2sbp,
  output [4-1:0]       uw1jajj_fvu9278tlptmv_, 
  output [4-1:0]       tdwhghf609ku2jek72pn3, 
  output [64-1:0]          cc7_9__0hrnupts,     
  output [64-1:0]          pba2_zyealgm_jf64t, 

  output                           r26sxdceh7f2t6xroiyejiud7e,
  output [7:0]                     pcmvrs0wuwr_x06ql,
  output [2:0]                     du9lzthd93rvmfcw7rz0wap,  
  output [4*8-1:0]   nabilb10azux1hnithsys,
  output                           q2vmic6hc_08xqnvwhw,
  output                           v175vi3kjhjhl37_p,
  output                           vir1r5sxmryfghdpp_u82bq6,
  output                           soumhrmo71_bkr9v6s5,
  output [2-1:0]     fqx1jny69kgy_gimut,
  output [9-1:0]  sd2su0k2v13e1jhtkwj,
  output [64-1:0]       h_4gbwx46f8brur_wc    ,
  output [64-1:0]       ruzuip2lmd_5bjdch    ,
  output                           t7xboey2yuqaq15sxya1b5,
  output                           v4icsnfwb3y76_4utq,
  output [64-1:0]       u4560ic2z4t9ft8jb0rvw,
  output                           de7s4aih29brxnb18p,

  output                           vyis_kjmkr7org4mer  ,
  output                           n20czkexgpbptzj5w  ,
  output                           uvysjueb4qilrx7   ,
  output                           qd0yrkr028oru_36lsp9,
  output                           zkhg8302rekq3   ,
  output                           yjox8n6veh2dfp4   ,
  output                           xa_tll8bjyk6hu8 ,
  output                           r9098zakm9jc     ,
  output                           ye_x11o9y0je9god    ,
  output                           cmbn4qx1zcverw    ,
  output [48-1:0] fwpoqfymdxr45bq2,

  output                           rnub9co3myzraj2l,
  output                           azbeqtr4zo_xorty8,
  output                           fv_51fuukywshp7hm,
  output                           w20nxrvpdf716_,
  output                           x2ypwv3n6g8jsweuweebmhq,
  output                                dwvp6uc1acommla,
  output                                p8to9sivjjwpc0pn2bvf21se3,
  output [105-1:0]  x9t5ge71i97il9r8,
  output [50-1:0] n7fla3l_dqx9jnxul4,
  output                              vg7c1san7ef_,
  output                              umwzm3ilav51kmk7r,
  output                              c8l2f5n1fhxm76kt3vlu6jp,
  output [48-1:0]    hibevegtudxlh_nk6e8e,  
  output [64-1:0]             y6lolb8cmealsn6ev,
  output                              x2bck2rbbpoyqbz62ld0tg,
  output                              abkeecplc6ueo97vo24tg,
  output                              b_fk_j1filrux_uod,
  output                              oaedrllyjbu5y92f,
  output                              plgwduxqtms73miw0,
  output   [64-1:0]           mf_okovo5c__xpv1x,
  output   [64-1:0]           i1_2srs1sequ9t,
  output   [64-1:0]           a4aa8t_dofc7_82w,

  output                              q6sud8b_vapga5ru5c,
  output [48-1:0]    latkf6ie2l8fv5dg98qec,  
  output   [64-1:0]           azmawprujj_u7q6ofj,
  output   [64-1:0]           wigxwsu_39gcyutr_re,
  output   [64-1:0]           l0_j3191k35720flisiv,
  output   [64-1:0]           cf059q4pm79who8jb,


  output                           itofghyluwwiwmqnj_4imeao    ,
  output                           j47kiegbvv22z361yv9n5  ,
  output                           r75dlj23fr96kve4fzd8xpw2zn    ,
  output                           mx7juirxj661i6i9lns4hnnyw0ep  ,

  output                           pdns51exd9ffhf5pykv42sq ,
  output                           k09nslb_nkoy4r0t34xu6,
  output                           frehkmd0xqj4qeyqqodmp0onx7  ,
  output                           ms95k2pmbvtrb33p5oa2q       ,
  output                           r928tvy6d88uh6s9qun65udol2    ,
  output                           jtgchf8072p4v1h9xclp0t   ,
  output                           jekm9yqqqogc7_czwax0r6an_f   ,
  output [64-1:0]     vs9f2qtmvyxt6ycc5e_z47fnjr  ,
  output                           wvywyxp28r9wdwncg13zbc_6 ,
  output                           suaktr_howpmkqxx3p5j4   ,

  output                           ussyj508sxu9v0    ,

  output                           mnym6ha4fxtg2oqq9hlac5s1,
  output                           p6wfurur4eut85r8tktdi03zxb,
  output                           xxr9qx83ggzl9q98ig_ys5w60a,
  output                           lozr9fiy6p7y8rinc582m2bt2ha_xmf,
  output                           u78ade2idh660umk_1m66fdlksb9b,
  output [64-1:0]     z3j5lbdgqwmp5zmv4g_zn29fgvintdc,




  output                           p1kjflyurzeuxj,
  output                           yvjlu1e9eng5_5tme,
  output [4-1:0]    hh8nc68zrpki2m9r,

  output                           v8wv99vga5gkl8xhk7x9in,
  output                           ahfx5rs9jkdyw3b8ztscfx,
  output [4-1:0]    ts3_k4ergzh8upz7,
  output [64-1:0]          ktqya1x1mfi5j3q7,
  output                           z6njhanl_m_hv48x5i9y,
  output                           dvm_h24fnflt11prmyvme,
  output [4-1:0]    uvyubcp0tbk9yirhz,
  output [64-1:0]          ivoui15mvw3de5ds44,





  output                                   jm4ru1fdiqtw706w8,
  output [19-1:0]  j021ufdslrlb4m5c5h2,
  output [64-1:0]                  crr9jljkvi3gsixv1_v8,
  output [64-1:0]                  sca7p0942a6kocjqqvat,
  output [64-1:0]                  go_m73qp_w0p7abohs24,
  output                           pket_pq2m99ayix3fk5yps,
  output                           ty49bqt9pydf4fr50f89,

  input  gf33atgy,
  input  ru_wi
  );





  wire [64-1:0] nsph0, yk8g9nis;
  wire [64-1:0] ny6lnci;
  wire [64-1:0] frgsqzgn0;
  wire [64-1:0] ay1h7j45ex4sqr;
  wire [64-1:0] bihnkz;

  wire bgn0kteb_8_x8gy6;
  wire mprd8f9bcmzkm_m;
  wire ergtosintr_qu;
  wire wza0m_ubqdukti34;
  wire s1u27hydhjys;
  wire u13lvaym24h7;
  wire ijomb1x0;
  wire rdlfxqf8;
  wire ciaqg62qrzne;
  wire [4-1:0] c1suh2jqglqdt6, jprib8qcyar3osk6 , p2usgr1j2bdu2daclo8 ;
  wire [4-1:0] idmjx9akqjlxnru2v ;
  wire [64-1:0] zdyk61t1j,t8b69o0ss;
  wire [64-1:0]    qb3k8_95n0k5gblo;
  wire [32-1:0] cxea1bdq1t2;
  wire yegbnqo2n4,va2_bl8hseu5, mbdfs7v8w,r4r2y8p;
  wire i5w9n6x9c, ycw1qucy1, a7kf63mkflg, vmze27ob2cy;
  wire m18d45glia74ly;
  wire b129regxq_4_;
  wire [105-1:0]  u3ha2g0qwmeq4s;
  wire [50-1:0] kzjz3lqozt3dmzo;
  wire m4ym0905s8pyqg9bhvs;
  wire [64-1:0] ivik66aksp;
  wire [64-1:0] yfbph0f2bzthnh;
    wire [64-1:0]               oyd81my_twgbtz;

  wire                              zdykvgl_mc;
  wire                              k0ab90pinn8;
  wire                              cistktgs2yjqga_2e;
  wire [48-1:0]    tcd_45_gx4ssqq;  
  wire [64-1:0]             lk_h0xurtx;
  wire                              ax4ahtf316zoev;
  wire                              h7jd3bxg3vb5ki;
  wire                              mwxgcnv_5_jd;
  wire                              jqfj544dp2cb;
  wire                              xg4pg_p97h;
  wire [64-1:0]             h9_wdq7h6;
  wire [64-1:0]             k28peem24d9ts;
  wire [64-1:0]             y7eur82cjk9r; 

  wire                              cs5oy2n8k08rtw;
  wire [48-1:0]    ebpafsre29c1c;  
  wire [64-1:0]             u_x7t53qamy1ma_;
  wire [64-1:0]             lezhwkr_wxtgf;
  wire [64-1:0]             k8nsdxg9w21;
  wire [64-1:0]             w722m1qcnuznp;
  wire p428idthlk91;
  wire [19-1:0]  uiug3i4kuqimc;
  wire [64-1:0] bplid7_q2mwu6f9, xfmtyw53vycvz7ow, ylghhwm40190t;
  wire                      rj8vqubs4fbhoqdmdbutku;
  wire [64-1:0]  sl4ljoqdgrgf5xq   ;
  wire [64-1:0]  ltkf0drscru5nbk40   ;
  wire [48-1:0]  i5uwzakbdn;
  wire hw87q7y3ka1ce3cf;
  wire t34t4sxf0vge;
  wire xq7_8a4tmvq72qzi ;
  wire jvbb9wysosshvb9;
  wire e6scnj06m ,f5yetvw_f7,b3qg60ck8hbf;
  wire h2j202k2_h2;
  wire kr65vpwn31r279;
  wire fm4d1r6ip9d3;
  wire ujgkuoavh ;
  wire t7y6dm970g6nyutdm ;
  wire og5hyvaovkaj ;
  wire xvh8ja0ivjz ;
  wire ch9pg0w3st ;
  wire [4*8-1:0]      hxp04fxso6sgjraa5;
  wire [7:0]      jw77minock;
  wire [2:0]      a2mv_cpge41qs2p9lx;
  wire ng6l_wwjcq763yj;
  wire bidv0g7keket; 
  wire qj3kcyyo_mj4n4g;
  wire o93a_6syaiqzt83d7;
  wire wwq0ynqkhyyd88ysee;
  wire nhml4wi8atuicrq9;
  wire [64-1:0] ewn2ga5jg8g602f3;
  wire w0e45bp2c_69hv;
  wire suca9h8s7z2;
  wire [2-1:0] xx4eq74chgxf9;
  wire [9-1:0] yy98t18hg5sfal;


  wire   n5c5v69zesumwty    ;
  wire   dnyg2nba4qnttvpy_  ;
  wire   gcuafcqpbtm4jn4wl    ;
  wire   dsvgzb_ckrnd_7h3gwn52m  ;

  wire m1m8zl_robbyztr01mtvt73    ; 
  wire qi_vhihdg1g7krvsdp         ; 
  wire dr7shdz251oj346h      ; 
  wire d3um711skad08s3cghqj     ; 
  wire eqxz7pvl8qvj63dwx_nh     ; 
  wire [64-1:0] jf16idqnvj2k5c3jix    ; 
  wire n50a0572igbciguq5     ; 
  wire dd3aq4w2_otde7     ; 

  wire dt6w0zkcz72w6ctu_l     ; 
  wire foftuihyj2l66w_oto2_n  ; 
  wire er2z0hm5khvf9haqza4z6wxj ; 
  wire bi0ec7mchd7wzkb3_9begl ; 
  wire yjmz9fbw8j9ck09ty4j9k48f0j ; 
  wire [64-1:0] eljv84ctnizg2rl5rqnm23qboa_    ; 





  wire oy9al5d = cvqaktep17ac & h91pmjbyad1itr37;
  wire b7nkstim3k = oy9al5d ? hm3iwty3s1d4si2p4 : k0ab90pinn8; 
  wire cdlm5zrwv = oy9al5d ? z1et08p41uxcl76 : cs5oy2n8k08rtw; 
  wire wmdpf0pqd6_4 = oy9al5d ? (q5_q35rctah_ & vnc88f08k1s0obtnvb) : (zdykvgl_mc & ycw1qucy1); 
  wire w86hm036xqu9hguo = b7nkstim3k | cdlm5zrwv ;
  wire p_u7cog99yxpzfb7p9has = hm3iwty3s1d4si2p4 & (eph11j28sez0oftr7b[32:32] | eph11j28sez0oftr7b[33:33]);
  wire gy8nwlp18wmlu7lgswrw = k0ab90pinn8 & (tcd_45_gx4ssqq[32:32] | tcd_45_gx4ssqq[33:33]);
  wire qnim506cfe4egy7czi = oy9al5d ? p_u7cog99yxpzfb7p9has : gy8nwlp18wmlu7lgswrw; 

  wire mxn4wdlge = oy9al5d ? bf8iyrsqp4a2s : b129regxq_4_;


  wire s0aynip0upf = oy9al5d ? pwppbjb8emt8vd9_w : p428idthlk91;



  wire ei82smlw45m = !mxn4wdlge & !w86hm036xqu9hguo; 


  wire vumxz5fuj = (~e7nqb0p7cffw4lrkd) & oy9al5d; 
  wire cl1hpce = ei82smlw45m & vumxz5fuj; 
  wire amk_mv9we = mxn4wdlge & vumxz5fuj; 
  wire rrurxkl633 = w86hm036xqu9hguo & vumxz5fuj; 
  wire gy6ddml = akdv8vv97zk549v & k_wnu24cz94zwh8;
  wire [4-1:0] ofxcqyaipegys = oy9al5d ? x11xtpe4e78unv1ahgzinz4n : jprib8qcyar3osk6;
  wire [4-1:0] jyp69_3c6ce00h7e = oy9al5d ? ialrcyi5grz5o0hc0jyjuwv : p2usgr1j2bdu2daclo8;
  wire [4-1:0] e8fbphi7t5pf39a9p = oy9al5d ? wfpum3du8gc8hr_xuerx : idmjx9akqjlxnru2v;




  wire zu59zys2m8jihleqj7     = ((x11xtpe4e78unv1ahgzinz4n == cu1owrury8wsed      ) & b43m7n67rav8he & uwl7jm0d1lv0xpo);
  wire cb7hqu8c7d8syx3q92c5     = ((x11xtpe4e78unv1ahgzinz4n == mt1z8r_sz      ) & qcutfgh43gov5u4urt & u2l80pdclhyu1bl);
  wire ng1dz8t0x9rxyak2cuoh1     = ((x11xtpe4e78unv1ahgzinz4n == uc9k3lw_iehx      ) & s73raoa0ilom1wyi & uamf3ccv7ouhi18);
  wire hmq1zl_yqh54uolnv0_3ancr    = ((x11xtpe4e78unv1ahgzinz4n == radwr7skyhm3jqso5) & dnwb40nhmse7rcj0epzjo);
  wire cj9zgxzx7wnzpmqq124d9_3    = ((x11xtpe4e78unv1ahgzinz4n == zdid44qi3bv7q4phl) & omeribg0gbgvpn78urilv_a);
  wire yjhtq7j0ba644m7xvagubq   = ((x11xtpe4e78unv1ahgzinz4n == x4owqbu74zh_xxr    ) & jxogr1vy8jotyh8ivd2u);


  wire d_udvn_fhsozg79auof8s     = ((jprib8qcyar3osk6 == cu1owrury8wsed      ) & b43m7n67rav8he & uwl7jm0d1lv0xpo);
  wire eed38vcw6hq0srxd9ip82     = ((jprib8qcyar3osk6 == mt1z8r_sz      ) & qcutfgh43gov5u4urt & u2l80pdclhyu1bl);
  wire t2a8j16l8grlvqs7eu6mghk     = ((jprib8qcyar3osk6 == uc9k3lw_iehx      ) & s73raoa0ilom1wyi & uamf3ccv7ouhi18);
  wire z59arm4zrorwqg26_kh_    = ((jprib8qcyar3osk6 == radwr7skyhm3jqso5) & dnwb40nhmse7rcj0epzjo);
  wire g4zjt570w69eu_7omu9sz3id    = ((jprib8qcyar3osk6 == zdid44qi3bv7q4phl) & omeribg0gbgvpn78urilv_a);
  wire h2w2eu2td4ggopupheuyu4   = ((jprib8qcyar3osk6 == x4owqbu74zh_xxr    ) & jxogr1vy8jotyh8ivd2u);



  wire w8as4ber7dagal4e_g7     = ((ialrcyi5grz5o0hc0jyjuwv == cu1owrury8wsed      ) & b43m7n67rav8he & uwl7jm0d1lv0xpo);
  wire dpt_nw0clt5h3ktp95v9     = ((ialrcyi5grz5o0hc0jyjuwv == mt1z8r_sz      ) & qcutfgh43gov5u4urt & u2l80pdclhyu1bl);
  wire aqa4n9k_rlj0ymz0jk1     = ((ialrcyi5grz5o0hc0jyjuwv == uc9k3lw_iehx      ) & s73raoa0ilom1wyi & uamf3ccv7ouhi18);
  wire ahanzmie8jevvv7dc6ns    = ((ialrcyi5grz5o0hc0jyjuwv == radwr7skyhm3jqso5) & dnwb40nhmse7rcj0epzjo);
  wire jsj7wrauyipq88vo4729dxzg    = ((ialrcyi5grz5o0hc0jyjuwv == zdid44qi3bv7q4phl) & omeribg0gbgvpn78urilv_a);
  wire ba7jz59isnply2cgwqgh_yyts   = ((ialrcyi5grz5o0hc0jyjuwv == x4owqbu74zh_xxr    ) & jxogr1vy8jotyh8ivd2u);


  wire audnzsdj1_yzncr0q8vpu1m     = ((p2usgr1j2bdu2daclo8 == cu1owrury8wsed      ) & b43m7n67rav8he & uwl7jm0d1lv0xpo);
  wire cfld037px9t5ubeiaztk1c6     = ((p2usgr1j2bdu2daclo8 == mt1z8r_sz      ) & qcutfgh43gov5u4urt & u2l80pdclhyu1bl);
  wire g4lk01zbl21eovjceac     = ((p2usgr1j2bdu2daclo8 == uc9k3lw_iehx      ) & s73raoa0ilom1wyi & uamf3ccv7ouhi18);
  wire v3hx0p8qlgg1fxhefr8    = ((p2usgr1j2bdu2daclo8 == radwr7skyhm3jqso5) & dnwb40nhmse7rcj0epzjo);
  wire svxp1jfpzn7vh35v7gdg6jf    = ((p2usgr1j2bdu2daclo8 == zdid44qi3bv7q4phl) & omeribg0gbgvpn78urilv_a);
  wire j_f7voq6e5tbrpbsivfcn2x_4   = ((p2usgr1j2bdu2daclo8 == x4owqbu74zh_xxr    ) & jxogr1vy8jotyh8ivd2u);


  wire oc98mdlhakpty2xro5ube4o     = ((wfpum3du8gc8hr_xuerx == cu1owrury8wsed      ) & b43m7n67rav8he & uwl7jm0d1lv0xpo);
  wire pfv44wqws10yge4sybh     = ((wfpum3du8gc8hr_xuerx == mt1z8r_sz      ) & qcutfgh43gov5u4urt & u2l80pdclhyu1bl);
  wire jcckdr8jsrrek1l9g0uhc     = ((wfpum3du8gc8hr_xuerx == uc9k3lw_iehx      ) & s73raoa0ilom1wyi & uamf3ccv7ouhi18);
  wire ke9l3tx2o1y8h_6405bsg0yg    = ((wfpum3du8gc8hr_xuerx == radwr7skyhm3jqso5) & dnwb40nhmse7rcj0epzjo);
  wire c26lrzkz8chjwv1f9ajp7z    = ((wfpum3du8gc8hr_xuerx == zdid44qi3bv7q4phl) & omeribg0gbgvpn78urilv_a);
  wire uo2rtnhi0yk0zt59pz9t   = ((wfpum3du8gc8hr_xuerx == x4owqbu74zh_xxr    ) & jxogr1vy8jotyh8ivd2u);


  wire jdz8iwclaki25v4a_3qq5     = ((idmjx9akqjlxnru2v == cu1owrury8wsed      ) & b43m7n67rav8he & uwl7jm0d1lv0xpo);
  wire irc0gu8bhar5o492ipf8z     = ((idmjx9akqjlxnru2v == mt1z8r_sz      ) & qcutfgh43gov5u4urt & u2l80pdclhyu1bl);
  wire bd8q_o8t5950aeradu     = ((idmjx9akqjlxnru2v == uc9k3lw_iehx      ) & s73raoa0ilom1wyi & uamf3ccv7ouhi18);
  wire amk1gzymdqi1nmplv6j2kkb4    = ((idmjx9akqjlxnru2v == radwr7skyhm3jqso5) & dnwb40nhmse7rcj0epzjo);
  wire s6qbup8u3k_vhvfwxmwmhh8    = ((idmjx9akqjlxnru2v == zdid44qi3bv7q4phl) & omeribg0gbgvpn78urilv_a);
  wire rmuu4wlbib0jcamytbcy9l5   = ((idmjx9akqjlxnru2v == x4owqbu74zh_xxr    ) & jxogr1vy8jotyh8ivd2u);



  wire tzs42knj7_eryjzjtrz = zu59zys2m8jihleqj7 |cb7hqu8c7d8syx3q92c5 | ng1dz8t0x9rxyak2cuoh1 
                       | hmq1zl_yqh54uolnv0_3ancr|cj9zgxzx7wnzpmqq124d9_3|yjhtq7j0ba644m7xvagubq 
                       ;
  wire qlpxdzyu05l61708l = d_udvn_fhsozg79auof8s |eed38vcw6hq0srxd9ip82 | t2a8j16l8grlvqs7eu6mghk 
                       | z59arm4zrorwqg26_kh_|g4zjt570w69eu_7omu9sz3id|h2w2eu2td4ggopupheuyu4
                       ;   

  wire x2d2gww2ztt7jh5 = w8as4ber7dagal4e_g7 |dpt_nw0clt5h3ktp95v9 | aqa4n9k_rlj0ymz0jk1 
                       | ahanzmie8jevvv7dc6ns|jsj7wrauyipq88vo4729dxzg|ba7jz59isnply2cgwqgh_yyts  
                       ;
  wire tlunyp28yeovvupm = audnzsdj1_yzncr0q8vpu1m |cfld037px9t5ubeiaztk1c6 | g4lk01zbl21eovjceac 
                       | v3hx0p8qlgg1fxhefr8|svxp1jfpzn7vh35v7gdg6jf|j_f7voq6e5tbrpbsivfcn2x_4   
                       ;   

  wire gq8tvqe22letpz672jip = oc98mdlhakpty2xro5ube4o |pfv44wqws10yge4sybh | jcckdr8jsrrek1l9g0uhc 
                       | ke9l3tx2o1y8h_6405bsg0yg|c26lrzkz8chjwv1f9ajp7z|uo2rtnhi0yk0zt59pz9t  
                       ;
  wire ucox8xw5yglf0jr9 = jdz8iwclaki25v4a_3qq5 |irc0gu8bhar5o492ipf8z | bd8q_o8t5950aeradu 
                       | amk1gzymdqi1nmplv6j2kkb4|s6qbup8u3k_vhvfwxmwmhh8|rmuu4wlbib0jcamytbcy9l5
                       ;   


  wire [64-1:0] jfbrikll = kl8zh4diafqs;
  wire [64-1:0] nqoz3ir = jiartjoiycj2;
  wire [64-1:0] ot2kbo = dtypmpwq1q2j;
  wire [64-1:0] jujagfre4ih3ec = pkw60eo867gghh;
  wire [64-1:0] d2zp8wdrny5zn_p = strg8286lgex8p4_0m;
  wire [64-1:0] e_j8qusu0gzawi1a = avpvrch0prpui67;


  wire [64-1:0] y_pzu3lb8d8df = 
                ({64{zu59zys2m8jihleqj7 }} &        jfbrikll) 
              | ({64{cb7hqu8c7d8syx3q92c5 }} &        nqoz3ir) 
              | ({64{ng1dz8t0x9rxyak2cuoh1 }} &  ot2kbo)
              | ({64{hmq1zl_yqh54uolnv0_3ancr}} &  jujagfre4ih3ec) 
              | ({64{cj9zgxzx7wnzpmqq124d9_3}} &  d2zp8wdrny5zn_p) 
              | ({64{yjhtq7j0ba644m7xvagubq}} &  (e_j8qusu0gzawi1a)) 
              ;
  wire [64-1:0] d5pokq9kkxbp = 
                ({64{d_udvn_fhsozg79auof8s }} &        jfbrikll) 
              | ({64{eed38vcw6hq0srxd9ip82 }} &        nqoz3ir) 
              | ({64{t2a8j16l8grlvqs7eu6mghk }} &  (ot2kbo))
              | ({64{z59arm4zrorwqg26_kh_}} &  jujagfre4ih3ec) 
              | ({64{g4zjt570w69eu_7omu9sz3id}} &  d2zp8wdrny5zn_p) 
              | ({64{h2w2eu2td4ggopupheuyu4}} &  (e_j8qusu0gzawi1a)) 
              ;

  wire [64-1:0] xv5to55_4wd = 
                ({64{w8as4ber7dagal4e_g7 }} &        jfbrikll) 
              | ({64{dpt_nw0clt5h3ktp95v9 }} &        nqoz3ir) 
              | ({64{aqa4n9k_rlj0ymz0jk1 }} &  (ot2kbo))
              | ({64{ahanzmie8jevvv7dc6ns}} &  jujagfre4ih3ec) 
              | ({64{jsj7wrauyipq88vo4729dxzg}} &  d2zp8wdrny5zn_p) 
              | ({64{ba7jz59isnply2cgwqgh_yyts}} &  (e_j8qusu0gzawi1a)) 
              ;
  wire [64-1:0] e_bpogyelz0h = 
                ({64{audnzsdj1_yzncr0q8vpu1m }} &        jfbrikll) 
              | ({64{cfld037px9t5ubeiaztk1c6 }} &        nqoz3ir) 
              | ({64{g4lk01zbl21eovjceac }} &  (ot2kbo))
              | ({64{v3hx0p8qlgg1fxhefr8}} &  jujagfre4ih3ec) 
              | ({64{svxp1jfpzn7vh35v7gdg6jf}} &  d2zp8wdrny5zn_p) 
              | ({64{j_f7voq6e5tbrpbsivfcn2x_4}} &  (e_j8qusu0gzawi1a)) 
              ;

  wire [64-1:0] zdtbiubtnca3d7 = 
                ({64{oc98mdlhakpty2xro5ube4o }} &        jfbrikll) 
              | ({64{pfv44wqws10yge4sybh }} &        nqoz3ir) 
              | ({64{jcckdr8jsrrek1l9g0uhc }} &  (ot2kbo))
              | ({64{ke9l3tx2o1y8h_6405bsg0yg}} &  jujagfre4ih3ec) 
              | ({64{c26lrzkz8chjwv1f9ajp7z}} &  d2zp8wdrny5zn_p) 
              | ({64{uo2rtnhi0yk0zt59pz9t}} &  (e_j8qusu0gzawi1a)) 
              ;
  wire [64-1:0] rqnwqusf0x5gy = 
                ({64{jdz8iwclaki25v4a_3qq5 }} &        jfbrikll) 
              | ({64{irc0gu8bhar5o492ipf8z }} &        nqoz3ir) 
              | ({64{bd8q_o8t5950aeradu }} &  (ot2kbo))
              | ({64{amk1gzymdqi1nmplv6j2kkb4}} &  jujagfre4ih3ec) 
              | ({64{s6qbup8u3k_vhvfwxmwmhh8}} &  d2zp8wdrny5zn_p) 
              | ({64{rmuu4wlbib0jcamytbcy9l5}} &  (e_j8qusu0gzawi1a)) 
              ;


  wire [64-1:0] wbkfq64ah9 = mn8sk0gr9oh54zn_o ? y_pzu3lb8d8df : kh00jq7wde_slaj;
  wire [64-1:0] awpq068vos = oetzq1g528ymdza0maph ? xv5to55_4wd : rezwnhzl7vmkg;
  wire [64-1:0] qj5940g9m = bwsazwvhtn9in7lpyjssdk ? zdtbiubtnca3d7 : nq_d1dxi6n86s;
  wire [64-1:0] fez_yrwve3h = wza0m_ubqdukti34 ? d5pokq9kkxbp : nsph0;
  wire [64-1:0] k67tywvm9gpl = s1u27hydhjys ? e_bpogyelz0h : yk8g9nis;
  wire [64-1:0] bxmcxgi = u13lvaym24h7 ? rqnwqusf0x5gy  : ny6lnci;


  wire [64-1:0] d0vtqvwh6t2 = oy9al5d ? wbkfq64ah9 : fez_yrwve3h;
  wire [64-1:0] swbwo112tnd = oy9al5d ? awpq068vos : k67tywvm9gpl;
  wire [64-1:0] k9n6vqknux9 = oy9al5d ? qj5940g9m : bxmcxgi;

  wire iry8vuin9srt75m = (tzs42knj7_eryjzjtrz & mn8sk0gr9oh54zn_o) ; 
  wire w36v74h15xbskqsaro = (x2d2gww2ztt7jh5 & oetzq1g528ymdza0maph) ; 
  wire mhnhpspolpe_1g8_aa = (gq8tvqe22letpz672jip & bwsazwvhtn9in7lpyjssdk) ; 
  wire xvw8qq7frj_5t = (qlpxdzyu05l61708l & wza0m_ubqdukti34); 
  wire agtf8ysq1jyhkuqgf = (tlunyp28yeovvupm & s1u27hydhjys); 
  wire uujc0ia4q4lwgifdg1 = (ucox8xw5yglf0jr9 & u13lvaym24h7); 

  wire apzevf3rv_0a92m1 = oy9al5d ? iry8vuin9srt75m : xvw8qq7frj_5t;
  wire yy95v2lcrr0n8sm = oy9al5d ? w36v74h15xbskqsaro : agtf8ysq1jyhkuqgf;
  wire w9uw03y254ah = oy9al5d ? mhnhpspolpe_1g8_aa : uujc0ia4q4lwgifdg1;

  wire eumzg8wq90izxng_eu95oxm = (~iry8vuin9srt75m) & mn8sk0gr9oh54zn_o;
  wire i6ihojwqvaqothl9tnn = (~w36v74h15xbskqsaro) & oetzq1g528ymdza0maph;
  wire oj9p6ur5uz1rclr80yqsol = (~mhnhpspolpe_1g8_aa) & bwsazwvhtn9in7lpyjssdk;
  wire x4ob1mylgh7sk3ap27 = (~xvw8qq7frj_5t) & wza0m_ubqdukti34;
  wire y4yttfmw2lh009kvliv = (~agtf8ysq1jyhkuqgf) & s1u27hydhjys;
  wire e4uenegyxsfugkmm7gf = (~uujc0ia4q4lwgifdg1) & u13lvaym24h7;



  wire l3q8ztenzfi6x = gy6ddml & (~oy9al5d);


  wire rtxazwz =  (
           (oy9al5d & (~mn8sk0gr9oh54zn_o) & (dorqi70cvs05s | k5yu5na0oo41y)) 
           | (apzevf3rv_0a92m1 & (~l3q8ztenzfi6x)) 
           )
         ;

  wire n2e11ebegn = (
           (oy9al5d & (~oetzq1g528ymdza0maph) & (pgfbjdj832ly_ | n8g2a10i7cbowtvjhc)) 
           | (yy95v2lcrr0n8sm & (~l3q8ztenzfi6x)) 
           )
         ;
  wire y4rl0n0q = (
           (oy9al5d & (~bwsazwvhtn9in7lpyjssdk) & (z0yti764_a15nwanb )) 
           | (w9uw03y254ah & (~l3q8ztenzfi6x)) 
           )
         ;





        
        generate
        if (gdctpuyrfi_b == 0) begin: hffbvgnj42j9fgv3ujrsxmkc1
          ux607_gnrl_dfflr #(64) b0ij0hrcdv98c (rtxazwz, d0vtqvwh6t2  , nsph0, gf33atgy, ru_wi);
          ux607_gnrl_dfflr #(64) sbarltevx0u (n2e11ebegn, swbwo112tnd  , yk8g9nis, gf33atgy, ru_wi);
          ux607_gnrl_dfflr #(64) oeamlq7aubxt (y4rl0n0q, k9n6vqknux9  , ny6lnci, gf33atgy, ru_wi);

          assign frgsqzgn0 = nsph0; 
          assign ay1h7j45ex4sqr = yk8g9nis;    
          assign h9_wdq7h6 = {64{1'b0}}; 
          assign k28peem24d9ts = {64{1'b0}};    
          assign y7eur82cjk9r = {64{1'b0}};    
            assign ivik66aksp = {64{1'b0}}; 
            assign yfbph0f2bzthnh = {64{1'b0}};    
            assign oyd81my_twgbtz = {64{1'b0}};    
        end else begin: ovxrovwx61jsf8u23zjms
          
          wire ct7dah3_yijtngy = ei82smlw45m & rtxazwz;
          wire d88yulyt88_pw = ei82smlw45m & n2e11ebegn;
          ux607_gnrl_dfflr #(64) x7ui4zrydbedvt (ct7dah3_yijtngy, d0vtqvwh6t2  , frgsqzgn0, gf33atgy, ru_wi);
          ux607_gnrl_dfflr #(64) kcitljusc04fhvs (d88yulyt88_pw, swbwo112tnd  , ay1h7j45ex4sqr, gf33atgy, ru_wi);

          
            wire jstj89yvwkd5k = mxn4wdlge & rtxazwz;
            wire ryh8jrgxzp8c_ = mxn4wdlge & n2e11ebegn;
            wire a08p6dqzdkzs = mxn4wdlge & y4rl0n0q;
            ux607_gnrl_dfflr #(64) ct7hmntqiavmkbmzw (jstj89yvwkd5k, d0vtqvwh6t2  , ivik66aksp, gf33atgy, ru_wi);
            ux607_gnrl_dfflr #(64) xma96v9qmy6ydhv (ryh8jrgxzp8c_, swbwo112tnd  , yfbph0f2bzthnh, gf33atgy, ru_wi);
            ux607_gnrl_dfflr #(64) treldqnonrph2nr9iz (a08p6dqzdkzs , k9n6vqknux9 , oyd81my_twgbtz, gf33atgy, ru_wi);

          
          wire fbbuaw3s584 = w86hm036xqu9hguo & rtxazwz;
          wire dw7k2sxaw00k = w86hm036xqu9hguo & n2e11ebegn;
          wire tijezy01rmn = w86hm036xqu9hguo & y4rl0n0q;
          ux607_gnrl_dfflr #(64) ec29tacm9cspo6 (fbbuaw3s584, d0vtqvwh6t2, h9_wdq7h6, gf33atgy, ru_wi);
          ux607_gnrl_dfflr #(64) hohiv4mgwzr332sa1 (dw7k2sxaw00k, swbwo112tnd, k28peem24d9ts, gf33atgy, ru_wi);
          ux607_gnrl_dfflr #(64) my1pdp9r1tsbuxn (tijezy01rmn, k9n6vqknux9, y7eur82cjk9r, gf33atgy, ru_wi);
          assign nsph0 = {64{1'b0}}; 
          assign yk8g9nis = {64{1'b0}};    
          assign ny6lnci = {64{1'b0}};    
        end
        endgenerate
  

  wire mxpzil60c4_2b;
  wire am9icjqa;
  wire enabtauddm3i;
  wire [5-1:0] xkx07g_p;

  ux607_gnrl_dfflr #(1) n4jlllh2dp63m_ (vumxz5fuj, k5yu5na0oo41y , mxpzil60c4_2b, gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1) kwe7alledqas (vumxz5fuj, n8g2a10i7cbowtvjhc , am9icjqa, gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1) b2bpyamq9chp6ah (vumxz5fuj, pzlsmt96uolwfb47 , enabtauddm3i, gf33atgy, ru_wi);


  ux607_gnrl_dfflr #(1) d9a49ivs11qitj1phkpmj (vumxz5fuj, aly0oms0x8r1kmmdgyob , bgn0kteb_8_x8gy6, gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1) ttmzrwajq_oy8lrw9 (vumxz5fuj, vckb4tc8r10z7n621obxkju , mprd8f9bcmzkm_m, gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1) deeosj3o0gd_miqzmc6vkg (vumxz5fuj, f3lw5s13_0u5q6o4ep , ergtosintr_qu, gf33atgy, ru_wi);


  wire k6l5_unp2j5swq = (oy9al5d | apzevf3rv_0a92m1); 
  wire p9y5qthv_fd9v02 = (oy9al5d | yy95v2lcrr0n8sm); 
  wire gwifxqjlicaezim_n = (oy9al5d | w9uw03y254ah); 


  wire drve_jpu7nsbilsa = oy9al5d ? eumzg8wq90izxng_eu95oxm : x4ob1mylgh7sk3ap27;
  wire cy4nzm6_1ruro5f0 = oy9al5d ? i6ihojwqvaqothl9tnn : y4yttfmw2lh009kvliv;
  wire ae33sheg72571frji = oy9al5d ? oj9p6ur5uz1rclr80yqsol : e4uenegyxsfugkmm7gf;




  ux607_gnrl_dfflr #(1) nr2zldr1y63pelnlmsy37 (k6l5_unp2j5swq, drve_jpu7nsbilsa  , wza0m_ubqdukti34, gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1) hkc07ites1nqbtb9hnb9a (p9y5qthv_fd9v02, cy4nzm6_1ruro5f0  , s1u27hydhjys, gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1) wik1tsyd6pa4_oom (gwifxqjlicaezim_n, ae33sheg72571frji  , u13lvaym24h7, gf33atgy, ru_wi);





  ux607_gnrl_dfflr #(1                  ) d8wfrjrz_yern           (vumxz5fuj , xxggjmznfu9b_           , mbdfs7v8w        , gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1                  ) axo3z09prx8f          (vumxz5fuj , mtsy6_whdwum2fu          , r4r2y8p       , gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1                  ) r55u_ictydnpe2mc         (vumxz5fuj , dorqi70cvs05s         , ijomb1x0      , gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1                  ) c25k7hn_zso45         (vumxz5fuj , pgfbjdj832ly_         , rdlfxqf8      , gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1                  ) kmqyo94hc5oe         (vumxz5fuj , z0yti764_a15nwanb         , ciaqg62qrzne       , gf33atgy, ru_wi);

  ux607_gnrl_dfflr #(4      ) q4amg04c1bl7wxxiwehf   (vumxz5fuj , ofxcqyaipegys          , jprib8qcyar3osk6, gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(4      ) tvjcv06a71heaxup3yezt8k   (vumxz5fuj , jyp69_3c6ce00h7e          , p2usgr1j2bdu2daclo8, gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(4      ) txtfpf5l9oq1dcqih8ku9un   (vumxz5fuj , e8fbphi7t5pf39a9p           , idmjx9akqjlxnru2v , gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(64         ) hwb_1w9e4h7lnl            (vumxz5fuj , t9kvx890cyg            , zdyk61t1j         , gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(64         ) l7jhaqngq3ln4es0         (cl1hpce , i984chc2gxtcivks        , t8b69o0ss     , gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(64      ) tlxfjudygg3x             (vumxz5fuj , cyudxl51e             , qb3k8_95n0k5gblo   , gf33atgy, ru_wi);

  ux607_gnrl_dfflr #(32   ) qgn4562n             (vumxz5fuj , nv33gk9s6_             , cxea1bdq1t2   , gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1                  ) vcj5axt7oqxq          (vumxz5fuj , tv7ak8mtfqswt          , e6scnj06m       , gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1                  ) dvhkwlqft931uz          (vumxz5fuj , axbsuznhe7w6rrd          , f5yetvw_f7       , gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1                  ) iqn10kmwrodxpt          (vumxz5fuj , j49by1lxo4ie9_ho          , h2j202k2_h2       , gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1                  ) k48tf7sgaewm_vbv         (vumxz5fuj , rtjejhmafpq7db         , i5w9n6x9c      , gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1                  ) w27xswaf5jg7e         (vumxz5fuj , vnc88f08k1s0obtnvb         , ycw1qucy1      , gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1                  ) cjusycc5w8ra3gqcg         (vumxz5fuj , u5pfnkzvz6fsvmgw4         , a7kf63mkflg      , gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1                  ) p91lt0r6bwukklzb         (vumxz5fuj , zlk2yur1jgjwg         , vmze27ob2cy      , gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1                  ) w1hv72r_t68z254c_vv   (vumxz5fuj , ow91ik9ily4bugcc43pp   , m18d45glia74ly, gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1                  ) pmcebpdipymvef        (vumxz5fuj , bf8iyrsqp4a2s         , b129regxq_4_      , gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(105 ) datvhtahg69o_s5da6 (amk_mv9we , j7l4qmkctu4k_1q6c       , u3ha2g0qwmeq4s    , gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(50) wkl9pc33k6jbo_a87x7 (amk_mv9we , x6t2ufv1z2uufogo       , kzjz3lqozt3dmzo    , gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1                  ) mo8i_nh0qy07rxg2rvt5_x(vumxz5fuj,  pu764metopn524rq4hg2c24  , m4ym0905s8pyqg9bhvs , gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1                   )   l2yt7wnn9j7a         (vumxz5fuj, q5_q35rctah_,       zdykvgl_mc          , gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1                   )   xl1scr9gp400fwr      (vumxz5fuj, hm3iwty3s1d4si2p4,    k0ab90pinn8       , gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1                   )   xazuisqsaokwhpgnv5x(vumxz5fuj, bod813pzaejozw9p1, xg4pg_p97h     , gf33atgy, ru_wi);

  ux607_gnrl_dfflr #(48 )   yw7enchstkr77hefl    (rrurxkl633, eph11j28sez0oftr7b,  tcd_45_gx4ssqq     , gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(64          )   nl0_78lzx_q3129_     (cl1hpce, lq6932o27hlk9v4f1m,   lk_h0xurtx      , gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1                   )   q37vzbyuij09c_wt0w  (vumxz5fuj, sll07sleuwo2fkitj,ax4ahtf316zoev   , gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1                   )   ls7yyg_p3eyukrqpfh2  (vumxz5fuj, v2e4q5r07qxd6fxruqia3f,h7jd3bxg3vb5ki   , gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1                   )   tm3lzvahk0x9snr_r7w  (vumxz5fuj, e5nqx8gg2u3gxy0y4c,mwxgcnv_5_jd   , gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1                   )   tylvk2slxa9jvza2926   (vumxz5fuj, ajka24wmafrwpta96cf2, jqfj544dp2cb    , gf33atgy, ru_wi);

  ux607_gnrl_dfflr #(1                  ) rxwv9hlswbjuzzzu851h     (vumxz5fuj , vh0cb71_xnjsewqur3     , hw87q7y3ka1ce3cf  , gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1                  ) fkglhiensw5ly2o8mfj4     (vumxz5fuj , gbgabhg8e_ul0e24r6jq     , t34t4sxf0vge  , gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(4      ) in087sdgbxzqur           (vumxz5fuj , z8xxe17sssy8tr8q219       , c1suh2jqglqdt6    , gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(48) hnt4v972qb0vh4hxj_9       (vumxz5fuj , juyjh9cdf4vvzhq       , i5uwzakbdn    , gf33atgy, ru_wi);

  ux607_gnrl_dfflr #(8                  ) oy8nx5nhq6saipgz61       (vumxz5fuj , mn3tic51ckga0gc       , jw77minock       , gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(3                  ) u83u3wmwys08libr972lb2tr  (vumxz5fuj , k0be3wres3xocvs9tpkn4fu  , a2mv_cpge41qs2p9lx  , gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(64      ) bhjy7_8py17fkkhrb1    (vumxz5fuj , rx4zxlit4v_5k4fclu    , sl4ljoqdgrgf5xq    , gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1                  ) hbzientvoid8tk1jmc47fn61ku(vumxz5fuj , vq3a19my9wldb5hug_nnbu0, rj8vqubs4fbhoqdmdbutku, gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(64      ) f1568wqw41pfla4y4br8     (vumxz5fuj , k_7iagb48feg9b3wj    , ltkf0drscru5nbk40    , gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(2    ) fwb2jo95cn8_umydy    (vumxz5fuj , ephp7dpea6ymyg0eucjv0    , xx4eq74chgxf9    , gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1                  ) xb6zw3xr98nh         (vumxz5fuj , kr13pzf9ml9ic_vbl         , suca9h8s7z2         , gf33atgy, ru_wi);

  wire g2uelalc59 = s0aynip0upf & vumxz5fuj;
  ux607_gnrl_dfflr #(1)                   fzxikiprqbzf7j9             (vumxz5fuj , pwppbjb8emt8vd9_w      , p428idthlk91      , gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(19) rq96f3keqpb4fujnnh5     (g2uelalc59 , z69pfny03ofcxvjyygmo6    , uiug3i4kuqimc    , gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(64) msy9xika388u4246ydfn (g2uelalc59, t9kvx890cyg  , ylghhwm40190t, gf33atgy, ru_wi);

  wire io8nnxty6dsz4n7fp_fyb19 = rtxazwz & s0aynip0upf;
  wire ilruiseabv5xbxz2uk8x1i = n2e11ebegn & s0aynip0upf;
  ux607_gnrl_dfflr #(64) n338figwjevypxyje8ji (io8nnxty6dsz4n7fp_fyb19, d0vtqvwh6t2[64-1:0], bplid7_q2mwu6f9, gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(64) w80ml0of2j5onev5g (ilruiseabv5xbxz2uk8x1i, swbwo112tnd[64-1:0], xfmtyw53vycvz7ow, gf33atgy, ru_wi);


  wire uwuie868 = cdlm5zrwv & vumxz5fuj;
  ux607_gnrl_dfflr #(1)                   kpcmk1lpy2nle1_r6c       (vumxz5fuj , z1et08p41uxcl76      , cs5oy2n8k08rtw      , gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(48) xor52un3mjou400adq     (uwuie868 , jymdjzitd0hv0e9uhul    , ebpafsre29c1c    , gf33atgy, ru_wi);

  
  wire dcosew6bka_yzfrg4k = rtxazwz & cdlm5zrwv;
  wire no_rbrxekhdasy0vblmu = n2e11ebegn & cdlm5zrwv;
  wire qspml1_58he2g9txiz = y4rl0n0q & cdlm5zrwv;
  ux607_gnrl_dfflr #(64) paja6r1ziaz066ab2 (dcosew6bka_yzfrg4k, d0vtqvwh6t2[64-1:0], u_x7t53qamy1ma_, gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(64) p05r65fj06tgbiyelie (no_rbrxekhdasy0vblmu, swbwo112tnd[64-1:0], lezhwkr_wxtgf, gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(64) he4pyt6lozp53xdi6l (qspml1_58he2g9txiz, k9n6vqknux9[64-1:0], k8nsdxg9w21, gf33atgy, ru_wi);

      ux607_gnrl_dfflr #(1                  ) qopwqdv3urxenoo_o      (vumxz5fuj, mylxtynzir7dvcouvb5thi   , gcuafcqpbtm4jn4wl   , gf33atgy, ru_wi);
      ux607_gnrl_dfflr #(1                  ) y3qsyfyuzx24euefb1bbj    (vumxz5fuj, o5yttui8un64i2r3s3yxxxjc25iwv , dsvgzb_ckrnd_7h3gwn52m , gf33atgy, ru_wi);



  generate
    if (t5462hhws9i6ynbxi == 0) begin: yk74rpnqrlfspp
      ux607_gnrl_dfflr #(5) h23ulh0a0vxbd (vumxz5fuj, uzn8ik3rkkwib6p , xkx07g_p, gf33atgy, ru_wi);
      ux607_gnrl_dfflr #(1                  ) u5jtabipbq5kqx         (vumxz5fuj , u4k7uyzg9lp3zlf         , b3qg60ck8hbf         , gf33atgy, ru_wi);
      ux607_gnrl_dfflr #(1                  ) pc1u7oqusmw8q           (vumxz5fuj , k_igx5_oeq1ag3m          , yegbnqo2n4          , gf33atgy, ru_wi);
      ux607_gnrl_dfflr #(1                  ) zwa3jmhhbwlpyma7       (vumxz5fuj , th3snuy_v19o06eanj      , va2_bl8hseu5      , gf33atgy, ru_wi);
      ux607_gnrl_dfflr #(1                  ) v62ojgl6ekmov7        (vumxz5fuj , w37tf6nz0oty_z89xv1        , kr65vpwn31r279        , gf33atgy, ru_wi);
      ux607_gnrl_dfflr #(1                  ) mtme1q15snt21rm        (vumxz5fuj , pfeci7n4c83yiwln58        , fm4d1r6ip9d3        , gf33atgy, ru_wi);
      ux607_gnrl_dfflr #(1                  ) sst1bnuk9h3ib         (vumxz5fuj , mzu7xfmjf4mwa0b         , ujgkuoavh         , gf33atgy, ru_wi);
      ux607_gnrl_dfflr #(1                  ) vnshm144gsrksbsxzcexv     (vumxz5fuj , g3t8ql0mi58ddizau_8t3     , t7y6dm970g6nyutdm     , gf33atgy, ru_wi);
      ux607_gnrl_dfflr #(1                  ) bg8ricpidysphdu_i         (vumxz5fuj , gg468ty1pm6_zgec         , og5hyvaovkaj         , gf33atgy, ru_wi);
      ux607_gnrl_dfflr #(1                  ) kr_6_w85z8b8x6j         (vumxz5fuj , jtvucg9wp5nxn         , xvh8ja0ivjz         , gf33atgy, ru_wi);
      ux607_gnrl_dfflr #(1                  ) at36i0y9oyxa77jcr6       (vumxz5fuj , ofe8xctslv6q5w48ky       , ch9pg0w3st        , gf33atgy, ru_wi);
      ux607_gnrl_dfflr #(4*8    ) xhpfbliib1udhhs__9ljyfj   (vumxz5fuj , lot9xvzuqrd5jm0scdx5t   , hxp04fxso6sgjraa5   , gf33atgy, ru_wi);
      ux607_gnrl_dfflr #(1                  ) qyp_xxwhuchqe        (vumxz5fuj , akk0_n8kvb1w0wxrz    , bidv0g7keket    , gf33atgy, ru_wi);
      ux607_gnrl_dfflr #(9 ) txqbnvr22_brxoi        (vumxz5fuj , w42z5c2wv916u4df79p        , yy98t18hg5sfal        , gf33atgy, ru_wi);

        assign w722m1qcnuznp = {64{1'b0}};
        assign cistktgs2yjqga_2e = 1'b0;

      assign bihnkz = {64{1'b0}};

      assign n5c5v69zesumwty   = 1'b0;
      assign dnyg2nba4qnttvpy_ = 1'b0;
      assign m1m8zl_robbyztr01mtvt73 = 1'b0  ; 
      assign qi_vhihdg1g7krvsdp      = 1'b0  ; 
      assign dr7shdz251oj346h   = 1'b0  ; 
      assign d3um711skad08s3cghqj  = 1'b0  ; 
      assign eqxz7pvl8qvj63dwx_nh  = 1'b0  ; 
      assign jf16idqnvj2k5c3jix = 64'b0  ; 
      assign xq7_8a4tmvq72qzi  = 1'b0;
      assign jvbb9wysosshvb9 = 1'b0;
      assign qj3kcyyo_mj4n4g = 1'b0;
      assign ng6l_wwjcq763yj = 1'b0;
      assign o93a_6syaiqzt83d7 = 1'b0;
      assign wwq0ynqkhyyd88ysee = 1'b0;
      assign nhml4wi8atuicrq9 = 1'b0;
      assign ewn2ga5jg8g602f3 = 64'b0;
      assign w0e45bp2c_69hv = 1'b0;
      assign n50a0572igbciguq5  = 1'b0  ; 
      assign dd3aq4w2_otde7    = 1'b0  ; 

      assign dt6w0zkcz72w6ctu_l = 1'b0; 
      assign foftuihyj2l66w_oto2_n = 1'b0; 
      assign yjmz9fbw8j9ck09ty4j9k48f0j = 1'b0;
      assign er2z0hm5khvf9haqza4z6wxj  = 1'b0  ; 
      assign bi0ec7mchd7wzkb3_9begl  = 1'b0  ; 
      assign eljv84ctnizg2rl5rqnm23qboa_ = 64'b0  ; 

    end else if (t5462hhws9i6ynbxi == 1) begin: yk74rpnqrlfspp
      ux607_gnrl_dfflr #(64         ) ef8o5dsk4d      (vumxz5fuj & (~vh0cb71_xnjsewqur3)  , plk8ixck4wj7c , bihnkz , gf33atgy, ru_wi);
      ux607_gnrl_dfflr #(1                  ) xqoarg69pxdxas8hku75cv4   (vumxz5fuj , wkixlev_tj12x_lfp6p04t   , xq7_8a4tmvq72qzi , gf33atgy, ru_wi);
      ux607_gnrl_dfflr #(1                  ) utgiud4l_p_e9djgm7474s11  (vumxz5fuj , jzx45r8bb79aj5ddz7h_565f  , jvbb9wysosshvb9, gf33atgy, ru_wi);
      ux607_gnrl_dfflr #(1                  ) ul3jyp7xvnfu7p3onugyib       (vumxz5fuj , s6in6vliinq9udhsofa      , qj3kcyyo_mj4n4g  , gf33atgy, ru_wi);
      ux607_gnrl_dfflr #(1                  ) w8dpkekzz03wa9uur1y_     (vumxz5fuj , cuxay1hemfm214cwu1513x     , ng6l_wwjcq763yj  , gf33atgy, ru_wi);
      ux607_gnrl_dfflr #(1                  ) yg9td2jxwoy5kgqh6ba9f4     (vumxz5fuj , cnp1c4afdljmpemgot3sa     , o93a_6syaiqzt83d7  , gf33atgy, ru_wi);
      ux607_gnrl_dfflr #(1                  ) zz30jhkl2512pp28nv_0a     (vumxz5fuj , wsh7h1p7b0zifvs0kwabih   , wwq0ynqkhyyd88ysee, gf33atgy, ru_wi);
      ux607_gnrl_dfflr #(1                  ) c80nbs3zehgh53_idkrsn      (vumxz5fuj , qhk0gez3kmex8twzly7mxn    , nhml4wi8atuicrq9, gf33atgy, ru_wi);
      ux607_gnrl_dfflr #(64      ) pn1iweyft797qz_cg     (vumxz5fuj , rafwujb8lw59lcbn9vsz8o   , ewn2ga5jg8g602f3, gf33atgy, ru_wi);
      ux607_gnrl_dfflr #(1)                   wj6hmbbxqfvuw8oxl       (vumxz5fuj , dqpwtmmizdh6bvzsx6     , w0e45bp2c_69hv, gf33atgy, ru_wi);
      assign b3qg60ck8hbf      = 1'b0;
      ux607_gnrl_dfflr #(1                  ) pc1u7oqusmw8q           (vumxz5fuj , k_igx5_oeq1ag3m          , yegbnqo2n4          , gf33atgy, ru_wi);
      ux607_gnrl_dfflr #(1                  ) zwa3jmhhbwlpyma7       (vumxz5fuj , th3snuy_v19o06eanj      , va2_bl8hseu5      , gf33atgy, ru_wi);
      ux607_gnrl_dfflr #(1                  ) v62ojgl6ekmov7        (vumxz5fuj , w37tf6nz0oty_z89xv1        , kr65vpwn31r279        , gf33atgy, ru_wi);
      ux607_gnrl_dfflr #(1                  ) mtme1q15snt21rm        (vumxz5fuj , pfeci7n4c83yiwln58        , fm4d1r6ip9d3        , gf33atgy, ru_wi);
      ux607_gnrl_dfflr #(1                  ) sst1bnuk9h3ib         (vumxz5fuj , mzu7xfmjf4mwa0b         , ujgkuoavh         , gf33atgy, ru_wi);
      ux607_gnrl_dfflr #(1                  ) vnshm144gsrksbsxzcexv     (vumxz5fuj , g3t8ql0mi58ddizau_8t3     , t7y6dm970g6nyutdm     , gf33atgy, ru_wi);
      ux607_gnrl_dfflr #(1                  ) bg8ricpidysphdu_i         (vumxz5fuj , gg468ty1pm6_zgec         , og5hyvaovkaj         , gf33atgy, ru_wi);
      ux607_gnrl_dfflr #(1                  ) kr_6_w85z8b8x6j         (vumxz5fuj , jtvucg9wp5nxn         , xvh8ja0ivjz         , gf33atgy, ru_wi);
      ux607_gnrl_dfflr #(1                  ) at36i0y9oyxa77jcr6       (vumxz5fuj , ofe8xctslv6q5w48ky       , ch9pg0w3st       , gf33atgy, ru_wi);
      ux607_gnrl_dfflr #(4*8    ) xhpfbliib1udhhs__9ljyfj   (vumxz5fuj , lot9xvzuqrd5jm0scdx5t   , hxp04fxso6sgjraa5   , gf33atgy, ru_wi);
      ux607_gnrl_dfflr #(1                  ) qyp_xxwhuchqe        (vumxz5fuj , akk0_n8kvb1w0wxrz    , bidv0g7keket    , gf33atgy, ru_wi);
      ux607_gnrl_dfflr #(9 ) txqbnvr22_brxoi        (vumxz5fuj , w42z5c2wv916u4df79p        , yy98t18hg5sfal        , gf33atgy, ru_wi);

        assign w722m1qcnuznp = {64{1'b0}};
        assign cistktgs2yjqga_2e = 1'b0;
        assign xkx07g_p = {5{1'b0}};

      assign n5c5v69zesumwty   = 1'b0;
      assign dnyg2nba4qnttvpy_ = 1'b0;
      assign m1m8zl_robbyztr01mtvt73 = 1'b0  ; 
      assign qi_vhihdg1g7krvsdp      = 1'b0  ; 
      assign dr7shdz251oj346h   = 1'b0  ; 
      assign d3um711skad08s3cghqj  = 1'b0  ; 
      assign eqxz7pvl8qvj63dwx_nh  = 1'b0  ; 
      assign jf16idqnvj2k5c3jix = 64'b0  ; 
      assign n50a0572igbciguq5  = 1'b0  ; 
      assign dd3aq4w2_otde7    = 1'b0  ; 

      assign dt6w0zkcz72w6ctu_l = 1'b0; 
      assign foftuihyj2l66w_oto2_n = 1'b0; 
      assign yjmz9fbw8j9ck09ty4j9k48f0j = 1'b0;
      assign er2z0hm5khvf9haqza4z6wxj  = 1'b0  ; 
      assign bi0ec7mchd7wzkb3_9begl  = 1'b0  ; 
      assign eljv84ctnizg2rl5rqnm23qboa_ = 64'b0  ; 

    end else if (gdctpuyrfi_b) begin: qhx9o35h2bu3u_l3n
      wire ezfdn1gnnda66 =vumxz5fuj & (~vh0cb71_xnjsewqur3); 
      ux607_gnrl_dfflr #(64         ) ef8o5dsk4d               (ezfdn1gnnda66 , plk8ixck4wj7c               , bihnkz , gf33atgy, ru_wi);
      ux607_gnrl_dfflr #(1                  ) ifrj9_35w2as8fq9nz    (vumxz5fuj, rgip60bn9st8htirgmhnohyj      , n5c5v69zesumwty   , gf33atgy, ru_wi);
      ux607_gnrl_dfflr #(1                  ) vqra4dcfxkcgxxf6415dub9  (vumxz5fuj, duo6acmepph_0ahl_0ebyyjh    , dnyg2nba4qnttvpy_ , gf33atgy, ru_wi);
      ux607_gnrl_dfflr #(1                  ) og8rk82ofwzd09irtdalogh3ls(vumxz5fuj, fxsynukaasxx8lt57bwdodyn3cem  , m1m8zl_robbyztr01mtvt73  , gf33atgy, ru_wi);
      ux607_gnrl_dfflr #(1                  ) y6bp99r33l3q857tw     (vumxz5fuj, oel93f4rkl6esczbag9yld       , qi_vhihdg1g7krvsdp       , gf33atgy, ru_wi);
      ux607_gnrl_dfflr #(1                  ) s1xggvoe1jbvmfa730huzv  (vumxz5fuj, vmp6zvyj46lrfmg3bl_kecu59    , dr7shdz251oj346h    , gf33atgy, ru_wi);
      ux607_gnrl_dfflr #(1                  ) vozyj3csob4_x6msp28tc3ah4 (vumxz5fuj, gj_lc7e2uh1cdx5b2bmynhvw   , d3um711skad08s3cghqj   , gf33atgy, ru_wi);
      ux607_gnrl_dfflr #(1                  ) a65q1_8_m46m6duwza0i9l (vumxz5fuj, b7ker79ak62g5qei_oa7kxdm0   , eqxz7pvl8qvj63dwx_nh   , gf33atgy, ru_wi);
      ux607_gnrl_dfflr #(64    ) v4z3871yyhpwy2eeq6szaxzsq_(vumxz5fuj, i3rcr_tmnynzs9lr254bac9x2b  , jf16idqnvj2k5c3jix  , gf33atgy, ru_wi);
      ux607_gnrl_dfflr #(1                  ) b31l0kch_1ooa_ww81ibql_   (vumxz5fuj, ti5a3yv8_m3rzzigzeuzrt1     , n50a0572igbciguq5    , gf33atgy, ru_wi);
      ux607_gnrl_dfflr #(1                  ) z4b18y1nq0nfi7wcl     (vumxz5fuj, cb86_62ddnv8i2whbc       , dd3aq4w2_otde7    , gf33atgy, ru_wi);
      ux607_gnrl_dfflr #(1                  ) owlk5rj5148st6hf979kd(vumxz5fuj, i_2lk2qupeba0sjgw6sdnbedc  , dt6w0zkcz72w6ctu_l  , gf33atgy, ru_wi);
      ux607_gnrl_dfflr #(1                  ) cti6libnf1qs1s41_0qtbdj1hexi(vumxz5fuj, a46z1a4rlrucmwj5ju3o83orp8jx2e  , foftuihyj2l66w_oto2_n  , gf33atgy, ru_wi);
      ux607_gnrl_dfflr #(1                  ) el46sqt53j261k44tyvr6_klirob(vumxz5fuj, p8zi9oi86dxmkaq4uqhu8j1hl0e  , er2z0hm5khvf9haqza4z6wxj  , gf33atgy, ru_wi);
      ux607_gnrl_dfflr #(1                  ) f4plrsbzxdxljreix5s4n1zm5uijj(vumxz5fuj, plmzz80_s0_tb0kwjjgu5p7uktpi2  , bi0ec7mchd7wzkb3_9begl  , gf33atgy, ru_wi);
      ux607_gnrl_dfflr #(1                  ) stroegmwky0r7tpa29p1ur0oak(vumxz5fuj, ti9h9knu4vrm6k3vqry9vfxbc4b  , yjmz9fbw8j9ck09ty4j9k48f0j  , gf33atgy, ru_wi);
      ux607_gnrl_dfflr #(64    ) pnipvjar7bmjfd_2iubynsx9wgw(vumxz5fuj, z_r1pp7wjooqw6n7rnoyv7nka81o, eljv84ctnizg2rl5rqnm23qboa_  , gf33atgy, ru_wi);
      ux607_gnrl_dfflr #(1                  ) xqoarg69pxdxas8hku75cv4    (vumxz5fuj, wkixlev_tj12x_lfp6p04t   , xq7_8a4tmvq72qzi , gf33atgy, ru_wi);
      ux607_gnrl_dfflr #(1                  ) utgiud4l_p_e9djgm7474s11   (vumxz5fuj, jzx45r8bb79aj5ddz7h_565f  , jvbb9wysosshvb9, gf33atgy, ru_wi);
      ux607_gnrl_dfflr #(1                  ) ul3jyp7xvnfu7p3onugyib       (vumxz5fuj , s6in6vliinq9udhsofa      , qj3kcyyo_mj4n4g  , gf33atgy, ru_wi);
      ux607_gnrl_dfflr #(1                  ) w8dpkekzz03wa9uur1y_      (vumxz5fuj, cuxay1hemfm214cwu1513x     , ng6l_wwjcq763yj  , gf33atgy, ru_wi);
      ux607_gnrl_dfflr #(1                  ) yg9td2jxwoy5kgqh6ba9f4  (vumxz5fuj , cnp1c4afdljmpemgot3sa     , o93a_6syaiqzt83d7  , gf33atgy, ru_wi);
      ux607_gnrl_dfflr #(1                  ) zz30jhkl2512pp28nv_0a     (vumxz5fuj , wsh7h1p7b0zifvs0kwabih   , wwq0ynqkhyyd88ysee, gf33atgy, ru_wi);
      ux607_gnrl_dfflr #(1                  ) c80nbs3zehgh53_idkrsn      (vumxz5fuj , qhk0gez3kmex8twzly7mxn    , nhml4wi8atuicrq9, gf33atgy, ru_wi);
      ux607_gnrl_dfflr #(64      ) pn1iweyft797qz_cg     (vumxz5fuj , rafwujb8lw59lcbn9vsz8o   , ewn2ga5jg8g602f3, gf33atgy, ru_wi);
      ux607_gnrl_dfflr #(1)                   wj6hmbbxqfvuw8oxl       (vumxz5fuj , dqpwtmmizdh6bvzsx6     , w0e45bp2c_69hv, gf33atgy, ru_wi);


      ux607_gnrl_dfflr #(1                  ) pc1u7oqusmw8q           (vumxz5fuj , k_igx5_oeq1ag3m          , yegbnqo2n4          , gf33atgy, ru_wi);
      ux607_gnrl_dfflr #(1                  ) zwa3jmhhbwlpyma7       (vumxz5fuj , th3snuy_v19o06eanj      , va2_bl8hseu5      , gf33atgy, ru_wi);
      ux607_gnrl_dfflr #(1                  ) v62ojgl6ekmov7        (vumxz5fuj , w37tf6nz0oty_z89xv1        , kr65vpwn31r279        , gf33atgy, ru_wi);
      ux607_gnrl_dfflr #(1                  ) mtme1q15snt21rm        (vumxz5fuj , pfeci7n4c83yiwln58        , fm4d1r6ip9d3        , gf33atgy, ru_wi);
      ux607_gnrl_dfflr #(1                  ) sst1bnuk9h3ib         (vumxz5fuj , mzu7xfmjf4mwa0b         , ujgkuoavh         , gf33atgy, ru_wi);
      ux607_gnrl_dfflr #(1                  ) vnshm144gsrksbsxzcexv     (vumxz5fuj , g3t8ql0mi58ddizau_8t3     , t7y6dm970g6nyutdm     , gf33atgy, ru_wi);
      ux607_gnrl_dfflr #(1                  ) bg8ricpidysphdu_i         (vumxz5fuj , gg468ty1pm6_zgec         , og5hyvaovkaj         , gf33atgy, ru_wi);
      ux607_gnrl_dfflr #(1                  ) kr_6_w85z8b8x6j         (vumxz5fuj , jtvucg9wp5nxn         , xvh8ja0ivjz         , gf33atgy, ru_wi);
      ux607_gnrl_dfflr #(1                  ) at36i0y9oyxa77jcr6       (vumxz5fuj , ofe8xctslv6q5w48ky       , ch9pg0w3st       , gf33atgy, ru_wi);
      ux607_gnrl_dfflr #(4*8    ) xhpfbliib1udhhs__9ljyfj   (vumxz5fuj , lot9xvzuqrd5jm0scdx5t   , hxp04fxso6sgjraa5   , gf33atgy, ru_wi);
      ux607_gnrl_dfflr #(1                  ) qyp_xxwhuchqe        (vumxz5fuj , akk0_n8kvb1w0wxrz    , bidv0g7keket    , gf33atgy, ru_wi);
      ux607_gnrl_dfflr #(9 ) txqbnvr22_brxoi        (vumxz5fuj , w42z5c2wv916u4df79p        , yy98t18hg5sfal        , gf33atgy, ru_wi);

      assign b3qg60ck8hbf      = 1'b0;

        ux607_gnrl_dfflr #(64  ) qx27hh20qdgdx3wr    (uwuie868 , lq6932o27hlk9v4f1m , w722m1qcnuznp  , gf33atgy, ru_wi);
        ux607_gnrl_dfflr #(1           ) qfruijqggdsa0mj18nlx7yp     (vumxz5fuj, txcys7e9ezk6xikpy2hu987,   cistktgs2yjqga_2e       , gf33atgy, ru_wi);

        assign xkx07g_p = {5{1'b0}};



    end else begin: uu6n368x9tf27mn
      ux607_gnrl_dfflr #(64         ) ef8o5dsk4d      (vumxz5fuj & (~vh0cb71_xnjsewqur3)  , plk8ixck4wj7c , bihnkz , gf33atgy, ru_wi);
      assign b3qg60ck8hbf      = 1'b0;
      ux607_gnrl_dfflr #(1                  ) pc1u7oqusmw8q           (vumxz5fuj , k_igx5_oeq1ag3m          , yegbnqo2n4          , gf33atgy, ru_wi);
      ux607_gnrl_dfflr #(1                  ) zwa3jmhhbwlpyma7       (vumxz5fuj , th3snuy_v19o06eanj      , va2_bl8hseu5      , gf33atgy, ru_wi);
      ux607_gnrl_dfflr #(1                  ) v62ojgl6ekmov7        (vumxz5fuj , w37tf6nz0oty_z89xv1        , kr65vpwn31r279        , gf33atgy, ru_wi);
      ux607_gnrl_dfflr #(1                  ) mtme1q15snt21rm        (vumxz5fuj , pfeci7n4c83yiwln58        , fm4d1r6ip9d3        , gf33atgy, ru_wi);
      ux607_gnrl_dfflr #(1                  ) sst1bnuk9h3ib         (vumxz5fuj , mzu7xfmjf4mwa0b         , ujgkuoavh         , gf33atgy, ru_wi);
      ux607_gnrl_dfflr #(1                  ) vnshm144gsrksbsxzcexv     (vumxz5fuj , g3t8ql0mi58ddizau_8t3     , t7y6dm970g6nyutdm     , gf33atgy, ru_wi);
      ux607_gnrl_dfflr #(1                  ) bg8ricpidysphdu_i         (vumxz5fuj , gg468ty1pm6_zgec         , og5hyvaovkaj         , gf33atgy, ru_wi);
      ux607_gnrl_dfflr #(1                  ) kr_6_w85z8b8x6j         (vumxz5fuj , jtvucg9wp5nxn         , xvh8ja0ivjz         , gf33atgy, ru_wi);
      ux607_gnrl_dfflr #(1                  ) at36i0y9oyxa77jcr6       (vumxz5fuj , ofe8xctslv6q5w48ky       , ch9pg0w3st       , gf33atgy, ru_wi);
      assign hxp04fxso6sgjraa5 = 8'b0;
      assign yy98t18hg5sfal = 9'b0;
        assign w722m1qcnuznp = {64{1'b0}};
        assign cistktgs2yjqga_2e = 1'b0;
        assign xkx07g_p = {5{1'b0}};
    end


  endgenerate

  assign jdngc81st67hk8p = mxpzil60c4_2b;
  assign u4t194j1c9najq = am9icjqa;
  assign gkzjw6iff1idxo = enabtauddm3i;
  assign jcj76rmi3pqujm3v = xkx07g_p;
  
  
  assign p8to9sivjjwpc0pn2bvf21se3 = m4ym0905s8pyqg9bhvs;   

  assign v8zi5h4rj36jt = nsph0 ;
  assign livvja2ywo91o8v = yk8g9nis ;
  assign t5p9q190fm = ny6lnci ;



  assign dckyl_qt92wqvghtw3 = frgsqzgn0 ;
  assign vyug4w9rb9kj6bmwwu = ay1h7j45ex4sqr ;
  assign h40f1u8xaz57o3c = ivik66aksp ;
  assign bv8rdomgcr9w6r2z = yfbph0f2bzthnh ;
  assign ujgn98iv8k5xidjk = oyd81my_twgbtz ;

  assign fw_dplmj46w6 = bihnkz;

  assign ptu54kun7juh0           = ijomb1x0;   
  assign tsns5phts_z2fnf           = rdlfxqf8;   
  assign rsdyvyptjiksvewu           = ciaqg62qrzne;   
  assign zf1w750jg2mtdij           = r4r2y8p;   
  assign pw6i533r0oou6ub            = yegbnqo2n4;   
  assign getq71b86zu18ri7x        = va2_bl8hseu5;   
  assign iouqv7uynzgvde_v             = mbdfs7v8w;    

  assign h_4gbwx46f8brur_wc      = sl4ljoqdgrgf5xq    ;    
  assign ruzuip2lmd_5bjdch       = ltkf0drscru5nbk40    ;    
  assign nabilb10azux1hnithsys     = hxp04fxso6sgjraa5    ;    
  assign pcmvrs0wuwr_x06ql         = jw77minock    ;    
  assign du9lzthd93rvmfcw7rz0wap    = a2mv_cpge41qs2p9lx;   
  assign vir1r5sxmryfghdpp_u82bq6   = o93a_6syaiqzt83d7;
  assign t7xboey2yuqaq15sxya1b5      = wwq0ynqkhyyd88ysee;
  assign v4icsnfwb3y76_4utq       = nhml4wi8atuicrq9;
  assign u4560ic2z4t9ft8jb0rvw      = ewn2ga5jg8g602f3;
  assign de7s4aih29brxnb18p        = w0e45bp2c_69hv;
  assign v175vi3kjhjhl37_p       = ng6l_wwjcq763yj;
  assign soumhrmo71_bkr9v6s5       = qj3kcyyo_mj4n4g;
  assign fqx1jny69kgy_gimut      = xx4eq74chgxf9;
  assign sd2su0k2v13e1jhtkwj          = yy98t18hg5sfal;
  assign r26sxdceh7f2t6xroiyejiud7e  = rj8vqubs4fbhoqdmdbutku;   
  assign q2vmic6hc_08xqnvwhw          = bidv0g7keket;

  assign hb36pq8e0n24raht15       = wza0m_ubqdukti34;  
  assign xphk4z06widyipxfcjr       = s1u27hydhjys;  
  assign xcu8n5tos13pfc6jhw22       = u13lvaym24h7;  

  assign lbx9pnfl2z4is68kam      = bgn0kteb_8_x8gy6;
  assign hl9x8gmcd9k2ttm0hui2j      = mprd8f9bcmzkm_m;
  assign ioka849821_gx48yl9gk      = ergtosintr_qu;

  assign j9fcegru44_r74xlm2sbp     = jprib8qcyar3osk6;  
  assign uw1jajj_fvu9278tlptmv_     = p2usgr1j2bdu2daclo8;  
  assign tdwhghf609ku2jek72pn3     = idmjx9akqjlxnru2v;  
  assign cc7_9__0hrnupts              = zdyk61t1j;     
  assign pba2_zyealgm_jf64t          = t8b69o0ss; 
  assign zpdph1sve               = qb3k8_95n0k5gblo;      
  assign o9d_zhwhmsph               = cxea1bdq1t2;      
  assign dte0cay394mhjhkr         = c1suh2jqglqdt6;
  assign tp46wehs200pll2qi           = b3qg60ck8hbf;
  assign vyis_kjmkr7org4mer          = kr65vpwn31r279; 
  assign n20czkexgpbptzj5w          = fm4d1r6ip9d3; 
  assign uvysjueb4qilrx7           = ujgkuoavh ; 
  assign qd0yrkr028oru_36lsp9       = t7y6dm970g6nyutdm ; 
  assign zkhg8302rekq3           = og5hyvaovkaj ; 
  assign yjox8n6veh2dfp4           = xvh8ja0ivjz ; 
  assign xa_tll8bjyk6hu8         = ch9pg0w3st; 
  assign cmbn4qx1zcverw            = e6scnj06m; 
  assign r9098zakm9jc            = f5yetvw_f7; 
  assign ye_x11o9y0je9god            = h2j202k2_h2; 
  assign fwpoqfymdxr45bq2         = i5uwzakbdn;
  assign rnub9co3myzraj2l           = i5w9n6x9c;
  assign azbeqtr4zo_xorty8           = ycw1qucy1;
  assign fv_51fuukywshp7hm           = a7kf63mkflg;
  assign w20nxrvpdf716_           = vmze27ob2cy;
  assign x2ypwv3n6g8jsweuweebmhq     = m18d45glia74ly;
  assign dwvp6uc1acommla           = b129regxq_4_;
  assign x9t5ge71i97il9r8         = u3ha2g0qwmeq4s;
  assign n7fla3l_dqx9jnxul4         = kzjz3lqozt3dmzo;
  assign vg7c1san7ef_              = zdykvgl_mc;
  assign umwzm3ilav51kmk7r           = k0ab90pinn8;
  assign c8l2f5n1fhxm76kt3vlu6jp  = cistktgs2yjqga_2e;
  assign hibevegtudxlh_nk6e8e         = tcd_45_gx4ssqq;  
  assign y6lolb8cmealsn6ev          = lk_h0xurtx;
  assign x2bck2rbbpoyqbz62ld0tg       = ax4ahtf316zoev;
  assign abkeecplc6ueo97vo24tg       = h7jd3bxg3vb5ki;
  assign b_fk_j1filrux_uod       = mwxgcnv_5_jd;
  assign oaedrllyjbu5y92f        = jqfj544dp2cb;
  assign plgwduxqtms73miw0         = xg4pg_p97h ;
  assign mf_okovo5c__xpv1x          = h9_wdq7h6 ;
  assign i1_2srs1sequ9t          = k28peem24d9ts ;
  assign a4aa8t_dofc7_82w          = y7eur82cjk9r ;

  assign q6sud8b_vapga5ru5c           = cs5oy2n8k08rtw;
  assign latkf6ie2l8fv5dg98qec         = ebpafsre29c1c;  
  assign azmawprujj_u7q6ofj          = u_x7t53qamy1ma_ ;
  assign wigxwsu_39gcyutr_re          = lezhwkr_wxtgf ;
  assign l0_j3191k35720flisiv          = k8nsdxg9w21 ;
  assign cf059q4pm79who8jb          = w722m1qcnuznp ;


  assign pket_pq2m99ayix3fk5yps       = hw87q7y3ka1ce3cf;
  assign ty49bqt9pydf4fr50f89       = t34t4sxf0vge;
  assign itofghyluwwiwmqnj_4imeao     = n5c5v69zesumwty;
  assign j47kiegbvv22z361yv9n5   = dnyg2nba4qnttvpy_;
  assign r75dlj23fr96kve4fzd8xpw2zn  = gcuafcqpbtm4jn4wl  ;
  assign mx7juirxj661i6i9lns4hnnyw0ep= dsvgzb_ckrnd_7h3gwn52m;

  assign frehkmd0xqj4qeyqqodmp0onx7 = m1m8zl_robbyztr01mtvt73 & ycw1qucy1; 
  assign ms95k2pmbvtrb33p5oa2q      = qi_vhihdg1g7krvsdp      ; 
  assign r928tvy6d88uh6s9qun65udol2   = dr7shdz251oj346h   ; 
  assign jtgchf8072p4v1h9xclp0t  = d3um711skad08s3cghqj & ycw1qucy1; 
  assign jekm9yqqqogc7_czwax0r6an_f  = eqxz7pvl8qvj63dwx_nh & ycw1qucy1; 
  assign vs9f2qtmvyxt6ycc5e_z47fnjr = jf16idqnvj2k5c3jix ; 
  assign wvywyxp28r9wdwncg13zbc_6= n50a0572igbciguq5 ; 
  assign suaktr_howpmkqxx3p5j4  = dd3aq4w2_otde7   ; 

  assign mnym6ha4fxtg2oqq9hlac5s1  = dt6w0zkcz72w6ctu_l; 
  assign p6wfurur4eut85r8tktdi03zxb = foftuihyj2l66w_oto2_n; 
  assign xxr9qx83ggzl9q98ig_ys5w60a = er2z0hm5khvf9haqza4z6wxj; 
  assign lozr9fiy6p7y8rinc582m2bt2ha_xmf = bi0ec7mchd7wzkb3_9begl; 
  assign u78ade2idh660umk_1m66fdlksb9b = yjmz9fbw8j9ck09ty4j9k48f0j; 
  assign z3j5lbdgqwmp5zmv4g_zn29fgvintdc = eljv84ctnizg2rl5rqnm23qboa_; 



  assign pdns51exd9ffhf5pykv42sq     = xq7_8a4tmvq72qzi;    
  assign k09nslb_nkoy4r0t34xu6    = jvbb9wysosshvb9;    

  assign ussyj508sxu9v0           = suca9h8s7z2 ; 

  assign jm4ru1fdiqtw706w8        = p428idthlk91;
  assign j021ufdslrlb4m5c5h2      = uiug3i4kuqimc;
  assign crr9jljkvi3gsixv1_v8       = bplid7_q2mwu6f9;
  assign sca7p0942a6kocjqqvat       = xfmtyw53vycvz7ow;
  assign go_m73qp_w0p7abohs24       = ylghhwm40190t;





  assign p1kjflyurzeuxj          = s1u27hydhjys;
  assign yvjlu1e9eng5_5tme         = mprd8f9bcmzkm_m;
  assign hh8nc68zrpki2m9r        = p2usgr1j2bdu2daclo8;  
  assign v8wv99vga5gkl8xhk7x9in      = uamf3ccv7ouhi18;
  assign ahfx5rs9jkdyw3b8ztscfx     = s73raoa0ilom1wyi;
  assign ts3_k4ergzh8upz7         = uc9k3lw_iehx;
  assign ktqya1x1mfi5j3q7          = dtypmpwq1q2j;
  assign z6njhanl_m_hv48x5i9y      = 1'b1;
  assign dvm_h24fnflt11prmyvme     = jxogr1vy8jotyh8ivd2u;
  assign uvyubcp0tbk9yirhz         = x4owqbu74zh_xxr;
  assign ivoui15mvw3de5ds44          = avpvrch0prpui67;




wire wxhj90zyzedojn50gn, ylk4alw9to8n2a0x;
generate
if(t5462hhws9i6ynbxi == 0) begin: evkm_k2x24
  ac6zxmzb4w0hgrfychpxv_xj # (
   .tcebpmbl7g(0),
   .mhdlk(1),
   .onr7l(1)
  ) w92h1x_zwb9kh (
    .veibgbyke(e7nqb0p7cffw4lrkd), 
    .bw6ftrau0(cvqaktep17ac), 
    .eef2g8(h91pmjbyad1itr37), 
    .qbjvs30wtb(1'b0),
    .wqljp(wxhj90zyzedojn50gn),
    .h9378(ylk4alw9to8n2a0x),
    .dqgck5s(),

    .gf33atgy  (gf33atgy  ),
    .ru_wi(ru_wi)  
   );



    wire ofuz9yi1xj0ychlty = ((wza0m_ubqdukti34 ) & ( ycw1qucy1))
                          ;
    assign akdv8vv97zk549v     = ((~ofuz9yi1xj0ychlty) & wxhj90zyzedojn50gn);
    assign ylk4alw9to8n2a0x = ((~ofuz9yi1xj0ychlty) & k_wnu24cz94zwh8);
    assign pysgbgu5mzucuewf1    = wxhj90zyzedojn50gn;    


end
else if(gdctpuyrfi_b == 1) begin: gkgb_21bseosn
  ac6zxmzb4w0hgrfychpxv_xj # (
   .tcebpmbl7g(0),
   .mhdlk(1),
   .onr7l(1)
  ) w92h1x_zwb9kh (
    .veibgbyke(e7nqb0p7cffw4lrkd), 
    .bw6ftrau0(cvqaktep17ac), 
    .eef2g8(h91pmjbyad1itr37), 
    .qbjvs30wtb(1'b0),
    .wqljp(wxhj90zyzedojn50gn),
    .h9378(ylk4alw9to8n2a0x),
    .dqgck5s(),

    .gf33atgy  (gf33atgy  ),
    .ru_wi(ru_wi)  
   );



    wire thbe_978hpwxcic = (wza0m_ubqdukti34 
                         |  s1u27hydhjys
                         |  (u13lvaym24h7 & (~m4ym0905s8pyqg9bhvs))
                         )
                          ;
    assign akdv8vv97zk549v     = ((~thbe_978hpwxcic) & wxhj90zyzedojn50gn);
    assign ylk4alw9to8n2a0x = ((~thbe_978hpwxcic) & k_wnu24cz94zwh8);
    assign pysgbgu5mzucuewf1    = wxhj90zyzedojn50gn;    
   end
 else if (t5462hhws9i6ynbxi == 1) begin: njkssg06u37tleou4w
  ac6zxmzb4w0hgrfychpxv_xj # (
   .tcebpmbl7g(0),
   .mhdlk(1),
   .onr7l(1)
  ) w92h1x_zwb9kh (
    .veibgbyke(e7nqb0p7cffw4lrkd), 
    .bw6ftrau0(cvqaktep17ac), 
    .eef2g8(h91pmjbyad1itr37), 
    .qbjvs30wtb(1'b0),
    .wqljp(wxhj90zyzedojn50gn),
    .h9378(ylk4alw9to8n2a0x),
    .dqgck5s(),

    .gf33atgy  (gf33atgy  ),
    .ru_wi(ru_wi)  
   );





    wire thbe_978hpwxcic = (ej5tfrzf8ad7noezo8gdkb1xg4 | (ekmvur7r4qz7ea7htd&ndvqmbwgzq08mbdaxnn4))
                         ;
    assign akdv8vv97zk549v     = ((~thbe_978hpwxcic) & wxhj90zyzedojn50gn);
    assign ylk4alw9to8n2a0x = ((~thbe_978hpwxcic) & k_wnu24cz94zwh8);
    assign pysgbgu5mzucuewf1    = wxhj90zyzedojn50gn;  

 end else begin:q05tvvewoxcik9
   ux607_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(1)
  ) w92h1x_zwb9kh (
    .i_vld(cvqaktep17ac), 
    .i_rdy(h91pmjbyad1itr37), 
    .i_dat(1'b0),
    .o_vld(akdv8vv97zk549v),
    .o_rdy(k_wnu24cz94zwh8),
    .o_dat(),

    .clk  (gf33atgy  ),
    .rst_n(ru_wi)  
   );
    assign pysgbgu5mzucuewf1    = 1'b0;    
    assign wxhj90zyzedojn50gn = 1'b0;    
    assign ylk4alw9to8n2a0x = 1'b0;    
 end
 endgenerate

  assign g65q46nnz7gip0zyo = wxhj90zyzedojn50gn;

endmodule                                      























module ac6zxmzb4w0hgrfychpxv_xj # (


  parameter tcebpmbl7g = 0,
  parameter mhdlk = 1,
  parameter onr7l = 32
) (
  input           veibgbyke,
  input           bw6ftrau0, 
  output          eef2g8, 
  input  [onr7l-1:0] qbjvs30wtb,
  output          wqljp, 
  input           h9378, 
  output [onr7l-1:0] dqgck5s,

  input           gf33atgy,
  input           ru_wi
);

  genvar i;
  generate 

  if(mhdlk == 0) begin: kum1oxhw1b434q

      assign wqljp = bw6ftrau0;
      assign eef2g8 = h9378;
      assign dqgck5s = qbjvs30wtb;

  end
  else begin: r1f9lplxw0lya5z

      wire d35brwhbkm;
      wire xlzi7_mjg;
      wire xayqet0sd;
      wire ycgzbt;
      wire d0x7t39v;


      assign d35brwhbkm = bw6ftrau0 & eef2g8 ;

      assign xlzi7_mjg = wqljp & h9378;

      assign xayqet0sd = (d35brwhbkm | xlzi7_mjg   ) |  veibgbyke;
      assign d0x7t39v = (d35brwhbkm | (~xlzi7_mjg)) & (~veibgbyke);

      ux607_gnrl_dfflr #(1) hdti_6iaq (xayqet0sd, d0x7t39v, ycgzbt, gf33atgy, ru_wi);

      assign wqljp = ycgzbt;

      ux607_gnrl_dffl #(onr7l) tn7qvilprku (d35brwhbkm, qbjvs30wtb, dqgck5s, gf33atgy, ru_wi);


      if(tcebpmbl7g == 1) begin:lvfon_zgkwp229

          assign eef2g8 = (~ycgzbt);
      end
      else begin:ulbqsqnmhe2qhizmyx

          assign eef2g8 = (~ycgzbt) | xlzi7_mjg;
      end
  end
  endgenerate


endmodule 



















module pkdsokaky2kt15iive(
  input  [5-1:0] w42_wd9um28vh,
  input  [5-1:0] ssjx8h5cj3q4ffem,
  input  [5-1:0] rwby8vkzgm4y4r,
  output [64-1:0] vuv0917fanv19,
  output [64-1:0] j2xzlc7dmxgmtn6kmk,
  output [64-1:0] tkxnzh2vh65vfutt3,
  input  j8mbnycgbc8k4exus50,
  input  [5-1:0] uup8_48koujjsde7s4,
  input  [64-1:0] unb_5mvf3gc1403brsa,
  input  nlxthgp55i6f26ozu4n,
  input  [5-1:0] bhxoyk3s_9ylb3,
  input  [64-1:0] y9hqso2yg_rpfqu,
  input  ub63nbp2x73net910cs,
  input  [5-1:0] pi6em2fjks8g1zb87,
  input  [64-1:0] u04hsk__lriad8ii,

  output [64-1:0] rfe2lglwm,
  output [64-1:0] oxa8a6mj5,


  input  gc4b3kdcan6do88ta_,
  input  gf33atgy,
  input  ru_wi
  );

  wire [64-1:0] fbu76k [0:32-1];
  wire [32-1:0] leab8mqf;
  wire [64-1:0] fd91wbm1bxxy [0:32-1];

  wire [32-1:0] dio6f7bff1;
  wire [32-1:0] gk661s__xwp;
  wire [32-1:0] ju71blrrvb;



  genvar i;
  generate 

      for (i=0; i<32; i=i+1) begin:ubs_7gmy192w

        if(i==0) begin: g7cih43

            assign fbu76k[i] = 64'b0;
            assign fd91wbm1bxxy[i] = 64'b0;
            assign dio6f7bff1[i] = 1'b0;
            assign gk661s__xwp[i] = 1'b0;
            assign ju71blrrvb[i] = 1'b0;
            assign leab8mqf [i] = 1'b0;
        end
        else begin: oky_oycgk0rvj

            assign dio6f7bff1[i] = j8mbnycgbc8k4exus50 & (uup8_48koujjsde7s4 == i[5-1:0]) ;
            assign gk661s__xwp[i] = nlxthgp55i6f26ozu4n & (bhxoyk3s_9ylb3 == i[5-1:0]) ;
            assign ju71blrrvb[i] = ub63nbp2x73net910cs & (pi6em2fjks8g1zb87 == i[5-1:0]) ;

            assign leab8mqf[i] = dio6f7bff1[i] 
                             | gk661s__xwp[i]
                             | ju71blrrvb[i]
                             ;
            assign fd91wbm1bxxy[i] =   ({64{dio6f7bff1[i]}} & unb_5mvf3gc1403brsa) 
                                | ({64{gk661s__xwp[i]}} & y9hqso2yg_rpfqu)
                                | ({64{ju71blrrvb[i]}} & u04hsk__lriad8ii)
                                ;

            ux607_gnrl_dfflr #(64) ddzbam3h39f (leab8mqf[i], fd91wbm1bxxy[i], fbu76k[i], gf33atgy, ru_wi);
        end

      end
  endgenerate

  assign vuv0917fanv19 = fbu76k[w42_wd9um28vh];
  assign j2xzlc7dmxgmtn6kmk = fbu76k[ssjx8h5cj3q4ffem];
  assign tkxnzh2vh65vfutt3 = fbu76k[rwby8vkzgm4y4r];


  assign oxa8a6mj5 = fbu76k[1];
  assign rfe2lglwm = fbu76k[3];


  wire [64-1:0] adtau = fbu76k[0];
  wire [64-1:0] f49g58 = fbu76k[1];
  wire [64-1:0] rhgpt = fbu76k[2];
  wire [64-1:0] ollg7 = fbu76k[3];
  wire [64-1:0] xw = fbu76k[4];
  wire [64-1:0] qfmfb5 = fbu76k[5];
  wire [64-1:0] q1z9nzm = fbu76k[6];
  wire [64-1:0] cf6_ = fbu76k[7];
  wire [64-1:0] zq5iq = fbu76k[8];
  wire [64-1:0] ksc = fbu76k[9];
  wire [64-1:0] llw = fbu76k[10];
  wire [64-1:0] hcm2g84 = fbu76k[11];
  wire [64-1:0] rsq0n = fbu76k[12];
  wire [64-1:0] gdrdah = fbu76k[13];
  wire [64-1:0] ys7m = fbu76k[14];
  wire [64-1:0] aa8b73lt = fbu76k[15];
  wire [64-1:0] kzib = fbu76k[16];
  wire [64-1:0] mbigdy = fbu76k[17];
  wire [64-1:0] lf_yup = fbu76k[18];
  wire [64-1:0] j2tdf6cz = fbu76k[19];
  wire [64-1:0] si7g9wy1 = fbu76k[20];
  wire [64-1:0] afy6p = fbu76k[21];
  wire [64-1:0] p6aa8 = fbu76k[22];
  wire [64-1:0] cj9rozp4 = fbu76k[23];
  wire [64-1:0] a4c = fbu76k[24];
  wire [64-1:0] uno = fbu76k[25];
  wire [64-1:0] g904q85c = fbu76k[26];
  wire [64-1:0] egvo = fbu76k[27];
  wire [64-1:0] rk8z = fbu76k[28];
  wire [64-1:0] y3voy9l = fbu76k[29];
  wire [64-1:0] c_sbw3x9 = fbu76k[30];
  wire [64-1:0] kut = fbu76k[31];
  
  wire [64-1:0] nsv6t1_qdn_9 = fbu76k[0];
  wire [64-1:0] po3j538u = fbu76k[1];
  wire [64-1:0] p8o0_330gs = fbu76k[2];
  wire [64-1:0] v172ktljmnc = fbu76k[3];
  wire [64-1:0] p__wpn = fbu76k[4];
  wire [64-1:0] onpzsh_1vla = fbu76k[5];
  wire [64-1:0] m7o6c1 = fbu76k[6];
  wire [64-1:0] vrwxs314m4 = fbu76k[7];
  wire [64-1:0] nx8kfo39x7 = fbu76k[8];
  wire [64-1:0] y7x_60uvr38 = fbu76k[9];
  wire [64-1:0] btwin5wu = fbu76k[10];
  wire [64-1:0] e4yvsmyqy = fbu76k[11];
  wire [64-1:0] ac8s0g = fbu76k[12];
  wire [64-1:0] dmzvl9bxxfa = fbu76k[13];
  wire [64-1:0] fu7j595o = fbu76k[14];
  wire [64-1:0] nqfhlj1v = fbu76k[15];
  wire [64-1:0] jr0bnqhb = fbu76k[16];
  wire [64-1:0] bb855azalfz = fbu76k[17];
  wire [64-1:0] ubpvkwalpw = fbu76k[18];
  wire [64-1:0] loadfy = fbu76k[19];
  wire [64-1:0] ccwqq95kvj = fbu76k[20];
  wire [64-1:0] x7ycj11ozi = fbu76k[21];
  wire [64-1:0] nckhyppprc = fbu76k[22];
  wire [64-1:0] vh60h5r = fbu76k[23];
  wire [64-1:0] rp116vqit = fbu76k[24];
  wire [64-1:0] hm0vdu = fbu76k[25];
  wire [64-1:0] imqz29r = fbu76k[26];
  wire [64-1:0] eujduw3l6 = fbu76k[27];
  wire [64-1:0] gfe04i3 = fbu76k[28];
  wire [64-1:0] p349rzblig = fbu76k[29];
  wire [64-1:0] o1xbxqh = fbu76k[30];
  wire [64-1:0] zrj6l2yp = fbu76k[31];

endmodule




















module pxp_0xj1 (



  input  jjzotrbn, 
  output hw1_k1jmu,
  input  [32-1:0] j3oz8j2,
  input  [64-1:0] bwjyqadn,   
  input  u2k4dyp52s_m ,
  input  djvj1e_ ,
  input  bktu0z1mk56 ,
  input  ipht6ss_sh6h,
  input  piwiqvrjoq,              
  input  al4xeg8mukgfg,               
  input  ryc6z1c7rmzrnlno,               
  input  rhufxsnopy0n,               
  input  wbhvg_1r9435,               
  input  s1woka0byzgo,             
  input  qhyq467foflgyn5y,               
  input  [64-1:0] binjv97px9r7dt04h0,
  input  ajl4tppx98ihuirj_mxih,
  input  sa2f4h4xeakpfnunl,               
  input  nrebzehsuam,
  input  [5-1:0] cpt0qfwiz,   
  input  [5-1:0] vf7a_1kae4zv5,   
  input  [5-1:0] djv9nstr,   
  input                          gy5zhpbrnl ,   
  input                          qv70a7n8p ,   
  input                          anlbkc8jny ,   


  input                          k405wpjt ,   
  input                          epi4op2w5ban9o ,   
  input                          heqeu11d07lcg2ss ,   
  input                          exzr5we0sujvtby ,   
  input                          anvecdxcx1ouoa0,   
  input                          x240tjzbog6i9q,   
  input                          uimia9sdhaq9x,   
  input  [5-1:0] bq9_5ksloh67_2ti,
  input  [5-1:0] qosgyc25p4fzq8b4,
  input  [5-1:0] cqk3fh13g1cxf9j,






  input  a02zzbowpjn06h,
  output st4f16aums5,
  output p05ld2ghmwh,



  output qbsr1jytrqtsbk4ttb8nz,

  output av1w8ld09cfofn,
  output im2b5l0h98avl6t4sj,
  output bw65wl7fvekfymd8vqx,
  output [64-1:0] pecbpcoa04vq,
  output [64-1:0] tb_snaxyfs,
  output [64-1:0] zc4mldgm25r,
  output [32-1:0] d23wb5yh1iyvf,
  output [1:0] srim3bfnzhve,
  output fvqwdz2hdbb,
  output cy3nuhzm_v2p73mt,

  output [64-1:0] ollg7,
  output d3n7pwgwcgze9cr4,
  output [64-1:0] amc4c8vcbecv1i,  
  output pby60vfdze02,
  output [64-1:0] vm3pyzc9nt95,
  output rbz4pv_atxqopdwt,
  output [64-1:0] qs1xgat7r8xow,

  input  [64-1:0] wd9dvepxj,

  output rm1dxjejhq7dh3q5m,
  output rvr30vvllni,
  output aw82i964do,

  input  dyl5g2vgrvy4mb3,
  input  r5hpbriny8m67sv9e_ylgo1,
  input umnrzb6pv8dzc,


  output                                   x8rpm78rvvycis, 
  input                                    h7lpiwlxyb79qyr06, 
  output [74-1:0] canacnkc7zibtkn418i, 
  input                                    bkkiffh6ob85nh79doya_, 
  input  [5:0]                             qhqqh0lyehgtfop1tc, 
  

  output                                   sxhicsqvufwfbnk0, 
  input                                    c5wzn6bil69i9toc, 
  output [74-1:0] x03ux1utw4qem5kk3c, 
  input                                    pjic5x84bqxpvdduy4r2s, 
  input                                    w5az87bw32r0tjbo0tdrv2ouvx, 








  output  hwpkcsh2atrq , 
  output  v3e6l1k7eo9k3 , 
  output  hxrmt706n071lic0f7, 
  input  [4*8-1:0] jt4l0g4njcsrt720n,
  output [4*8-1:0] w7uciar2_6p9xc5mc,
  input  [7:0] m9cdnl05ykr_3p,
  output [7:0] ex6ixmgf331,
  input  [2:0] akh3h7anvh7892ugn,
  output [2:0] vfu1cc_k9n55lt38g_vii,
  input   o_d157fc5_l,
  output  texy7g6tpvcgwtyd,
  input  [9-1:0] s68_9qhgnb_o,
  output  [9-1:0] q52oeddgdt76b,
  input  [2-1:0] oypxxr_e_rms7ai,
  output [2-1:0] gkps1gyqdwgzcvr0c,
  output  gfod0nmy6eta29jeeg6mr2,
  output  n4soswat5yihd74b,
  output [64-1:0] if0fog4bug_zkykpi,
  output q97rqfy8n7ixfm2a5wev4nd5sylpcq3j,
  output lln3b7iev7jpvogh964ro_9bc_3y,
  output hujgg6hjnhtbspbkekuz5_u,
  output v3pnt81kfrgbaanm1mhh51w,
  output [64-1:0] i08eq60d_snxeq8si_ezod,
  output dgnjyd9xs8efyxm0tdlsvfq4eop,
  output y8wz7aud_fd6dfiakjtx2i0g,
  output a3xib90kwk4_hm1,
  output nfzexr8q9g893gi,
  output [64-1:0] opkkwp3eg8g3448t,
  input   zsgl59ydqwjln,
  output  b9yq2alidby7zgom1,

  output  tvqijouldcgiz2dxdco7,  
  output  zkxlkidschdubxpkpm,  
  output  xmcrni1qngfvh9pil9j,  
  output  btkcf2uqr61gkiqhde0lai,  
  output  [64-1:0] h01d94xsxbxe_req,  
  output  w1casjl7bz73brz,  
  output  hjri7cufo9ckntq,  
  output  yghffofulqa77bd7aw07badta1a,
  output  rrl7evvmayt1_vvp74iq9h6_cjf,
  output  [27-1:0] zddoxp22m1o11x30gbe,
  output  [16-1:0] hwfethpzkuauejcgtbl6o,  

  input   n3ak8l6cvn0s4,
  output  hsxh9536ho4bw8o,
  output  r_edve7v9jcr26q6zk,  
  output  vrqfzuog2k4pos133,  
  output  bmw2yi333716crywk,  
  output  k2sr7sw1plcmnki5ajtscw,  
  output  [64-1:0] jkzw_f9anx55,  
  output  t8muv9e6d7yk_whqa0,  
  output  hzdfp71n6g3f5fsg5,  
  output  lwdhmuzyvcvv14mjbl0h2a41z,
  output  xy48dugh009wtmazqug3kpy2a5h_,
  output  [27-1:0] l4ztejmt2__wxqm2rw,
  output  [16-1:0] s3ujdp2a8n69bm6engxok,  


  output emc_bywzarijbo,
  output qo5p9t6s74zxpo,

  output tw5xnp59d8x,


  output [8*32-1:0] pcr4upio7_tx37   , 
  output [8*1-1:0]          uzklqlncpqqm1rav,
  output [8*1-1:0]          ortueunvnkx_l5m_j,
  output [8*1-1:0]          hwuhtb7ucto_utk56,
  output [8*2-1:0]          i1env2kmns7qvvuuc,
  output [8*1-1:0]          g3s3vpafvy3i,

  output                                 bz8qao4o4xqslni1d3,
  output [27-1:0]          vpecdc5kos, 
  output [1:0]                           pccd7o463jfc_dpc5va, 
  output                                 k5ovx8tintgvetip, 
  input                                  f97le_hyejv7saw9vslna, 
  input                                  yruel3nusosm39gnmb9ev_, 
  input                                  oeux55k_cre0he7w7jip5b1, 
  input  [55-1:0]     r8z2r_ud53zj8mrpk, 
  input                                  bu1949pq_9946o1_e2q_uvr8p4, 
  input                                  b4isf5u8b8pj34e09f72vxe38zg, 

  input                                  kvpemhoim1tq5y8mzwvix5, 
  
  output                                 z1l_kkshyf_56cwmaq2dm,
  output [16-1:0]          w7u50np_chxy7wq5n9et_q,
  output [20-1:0]            l2dse4sd3runnrb1rcbydauc, 
  output                                 kr1rhzlb5gr_wty1pe392s5oqet, 
  output [1:0]                           ox2ptuhum_e2aodz8wine6h, 
  output                                 g_qmxgznvfin609fmm97kuc2dm02, 
  output                                 i9oln6xm1pi9dzsd61s1kg4dmo7j, 
  output [1:0]                           hei_cs0rbwsv, 
  output                                 yf_5vs18cke5xg660my, 
  output                                 deo3wn_907tw886r,  

  output w92a5o09fp9dg6   ,
  output eglor15f7p2ivpny5dc   ,
  output ous_emkpecrqhg5e7,
  output doh50j3p7c7yl7uk9,
  output s7eq8f6z1uyi2in,

  output  um8zsjyxn_4p,  

  input  [64-1:0] v09gw6e6rfjf05qg,
  input  fcjh1nct4r,
  output x_cq40qmp6a,
  output z1l80uwh6vyyg34,
  input  rn1o3sl83,
  input  zz5wo47gw146x4,
  input  fgr486jx5kevbua,
  input  pvfk1_6o89lmby,
  input  xx87vzbpchg,

  
  
  input  c5ewdqztjw9za,
  input  rn2mt6nngsc9w5cz,

  output  [64-1:0] qeb3z0x5,
  output  ibhfuwrztbm8p4gg,
  output  [3-1:0] i8_5wt0vppx,
  output  osv2437qj_3nuf,


  output  b7g_vsn0zoewh6g1,
  output  [2-1:0] onnv64ydiajl,
  input   [2-1:0] r21i4by0bu3ks,
  input  [64-1:0] hn85hkp2yav,

  input  [64*4-1:0] azll7rq5fab5ou,
  input  [64*4-1:0] n6a0r_0zddzrme8,
  output ns0i7siujgkrghjpqv6,


  input  t5trf35s8vy,
  input  zbac123pv78sbz3,
  input  z4e_m564fxae0kpbjr,
  input  zmwq3e9oijvo7d7,
  input  hixy2y36a1pn0,
  input  ozwene1gdpatk6g,
  input  sxvvsxtbhyvt,

  output j0qaxhuqtdi,
  output pbzpk52jinfscit4mm,
  output gwj6ow6qvbhs0tc31,
  output iwdkm52x_w4hpak_a2_w,
  output [12-1:0] mm0ssgy582fv_j,
  output [64-1:0] ir2913p9xpmq_1bvfd1,
  input  [64-1:0] bsjo0v5e0t556pph,
  input  mwegg_7inaca6povsw,
  input  wnkp7091zrsevkbl,


  input  pydatzxqqi,
  input  c4ughu0qm5sfai,


 input [64-1:0] er2ibckhm98h98,
 input [64-1:0] tmi776v7orl,


 input [64-1:0] ndn228hd1n2x,
 input [64-1:0] kwk_z0jwwa2r,
 input [64-1:0] fnbi_cp8jq6t9ropn,


 output [5-1:0] cjo14q6bim0c,   
 output [5-1:0] yqawr6m8r98vjx73,   
 output [5-1:0] wuzzw7m7hpf4p6q31,   
 output [48-1:0] zscjnjl4ffiey84zel2,  
 output [64-1:0] qy0ycb_z4ngy2ll8pqo,
 output nb2chelz4_ijwumv9murokla,
 output bcrcin74qehflgu36ch9ghyv,
 output fbzipldpa3ewvv31mgr,
 output nlptjpg_zybrljgsnky1iwvhf,
 output zgv8w7jqb5wr6l2elow5znmm,
 output rpceina94e3bcz2ov7g1t_iom,


 output                           c4i0yanuek7va0ztp ,
 output [48-1:0] n5x33q1l9ewebt6692qaofd8,  
 output [64-1:0]          eqhoch739wo4sqhno2u,
 output [64-1:0]          qj1fn7kk041c_7kez4t2fkt,
 output [64-1:0]          q2qa0la3s98x10a2aqsb73g,
 output [64-1:0]          ajk1fk4kecwsdaeiybv,





  input                          vz63qkw5s3m8urb9, 
  input  [64-1:0]        iojqlhtwx45_siz,
  input  [4 -1:0] ydtm1yuxqj7fmxvqc,

  input                         o4qff84vfbn, 
  output                        x74_jhmpouk, 
  input  [64-1:0]       z5tnbveujliw633sxlb8,
  input  [4 -1:0]l8ng5e_pa1fg07__37,
  input                         erdoc9bbdnq8065yw , 
  input                         zqx1cj9lvt0e,
  input                         zsxgccndqw2suf6,
  input  [64-1:0] y9389ymcyh2ia2082yx1_,
  input  [64 -1:0]   uiu4_g7j41kz,
  input                         ro93aearv5754gz9w , 
  input                         rqy9v1_k_o74etonfc , 
  input  [4:0]                  ytp8_jsqr2sjmu08gdn,
  input                         b0ylmw5xa8oytsw3j6n,












  input                         flcopog5zzpohfautwy, 
  output                        gtb8f_h0g28itdr8k, 
  input                         wf15djwi2hw25nz_  , 
  input                         t1q5qmk9jzpf6glng4y,
  input [64-1:0]        xsmx4zoewhbt07jxq,
  output                        xmbe_e4vm6ofjbn7lq,

  output y_0q8d40rrzolo1y6,
  input  ao17frh5wnr0wddz3,
  output  mmludd_fnt2yevok8a1a0,
  input   buwj9_8l8bwj80kkinq9p,


  output um28jgd2x4mbs,
  output [64-1:0] l_imk5zs8ejjka,
  output [64-1:0] lz3vnoxnz_z,
  output yhbtmo4kyz_ewog3,
  output cd4d2_i3rcc1_p,
  output [5-1:0] wyu42gj62n994v0wo_,
  output x9cmkt53yq483z1,
  output cxmwxfttqy2t7ura   ,
  output b5wruck8tj9sa   ,
  output bxentpryfwb3d  ,
  output o2a43mjdbgea1  ,




  output                         o21b8ypt1xiu5ml63d,


  output                         badsf4ksbp3k6p_p5hnj2i, 
  input                          ed4kcy8s9nrisftgx_q, 
  output [32-1:0]   bdqo1tgw2_bpi2e8alini, 
  output                         jp5nha2l14e7kx2jzpke,   
  output                         c1gmncmorg16sachdas,  
  output                         za9xg3zsqni_aeqmke,  
  output [64-1:0]        a4a48egkdkec8d9b_9, 
  output [8-1:0]     xwfmltfzahuj4qfn4qf2, 
  output                         p648zxn2luyxy8mt992a,
  output                         uxlldm0w_h7kicit8gvhqv2,
  output                         yvu98r_7ji4o250r_u,
  output                         zdpamqgv7ddf1n3x5t2q,
  output                         wpsukhyqhl92dzoam7cm,
  output                         v3oo69y614hgiemyyld,
  output [1:0]                   ggxoqcj7ytp1a4pjf7ee,
  output                         l3c127qdc9a2mfc13,
  output [4 -1:0] oq9b5zfhza9yvdoj,
  output [4:0]                   szrgf24or2mbt7w_yleh_vt,

  output                         sg33s7pt45jp_ ,

  output                           p1kjflyurzeuxj,
  output                           yvjlu1e9eng5_5tme,
  output [4-1:0]       hh8nc68zrpki2m9r,

  output                           v8wv99vga5gkl8xhk7x9in,
  output                           ahfx5rs9jkdyw3b8ztscfx,
  output [4-1:0]       ts3_k4ergzh8upz7,
  output [64-1:0]          ktqya1x1mfi5j3q7,

  output                           z6njhanl_m_hv48x5i9y,
  output                           dvm_h24fnflt11prmyvme,
  output [4-1:0]       uvyubcp0tbk9yirhz,
  output [64-1:0]          ivoui15mvw3de5ds44,

  output                           n3zlo14nquu5l7zf3,

  output                           a_1o1o8345o28hui,
  output                           t8p1kh0tvb2ej56s  ,
  input                          p7ah58va5_2njbtv,
  input [64-1:0]         u981qrwkgi5h0e72b__gg19w,
  input                          p0i2i3v3j1tclelx51,
  
  
  
  
  
  
  
  

  
  
  


  input                            f0jwv0n5olimpf4vnvqpb4hs,



  output  yixt0a_xmh        ,
  output  ej7frm_ut9j6y    ,
  output  izjeme5aukvcc    ,
  output  uzevp4zrbs9gi,

  input   uc5qxb4d2b28ye5,
  output  o2qkf90r783,


  output habgbg2jn3qi,
  output dg4hzu_,
  output h7fseh5_df0hbx,




  input enwn0u48p2_ls5az80,
  output [7:0] f_i1959b4xizzq9jea,
  input [9:0] b4lwcgm6l21pi,
  input [7:0] hjrk_rwjkqj3zk_b,
  input zwcbp7zqfei5xz,
  input znzjygllppv1s0a8cqub3c, 
  output gfy3zost37aq8qmr,
  output dz0zrf512290tvcy4q,
  output dxi_ue3gf5zqqqxwgq2a,
  output ix299qulxi5    , 
  output jjj61w03m77lv    ,
  output dn8riluj40uunvq5,
  input miax48k27o484e8a,
  output fzdb65fcrotwcaccus_cwo,
  output [7:0] tcy_87vt9vet39knuw,
  input  fc_4ns_w1nh4h02z_dgg,
  input  jqsukc5b5drcc1e78,
  input  gnn46rd7vvofruqij,
  

  output y8_gkxsfle,

  output dkmuhc79d2wm0wubp,
  output u2demhkod_er3kf6b,
  input  uz7pt71lvqit85od,
  output [4-1:0] v3uvhtx7e5vbtvie,
  output [64-1:0] tmqkgmlzi018,
  output [64-1:0] lx_olubu7t8h,
  output [64-1:0] dd1p3tnenmm9r,
  output [3-1:0] l60zv02z95hlayri,
  input  l1xzyldaa9dr2q7mla,
  input  a5z_23_ryr_m29hhia_p ,

  output vejdvgqormu727s,
  output [64-1:0] ar9ro1ql86jzmq_p,
  output [5-1:0] qz1gqv6vh5qturw6v1mz,
  output ptyuk4efbbdu9asp0b8cmreeh,  
  

  input                          y7rd1k0an54clel_5q6, 
  output                         com03bquiktu249yb0, 
  input  [64-1:0]        tzg0yjgx9bn98i,
  input  [4 -1:0] c2mipfm_6z5ef4p3aoz,
  input                          y3z8rf7c6hvsiux , 
  input  [5-1:0]                 x8_a2j7z3gz3l0tfjqp,

  input  xq0mj5mg2_512eu4, 
  output e11m1298jo38qcwq9er2, 
  input  [64-1:0] ec94_mk193di7tj,
  input  [4 -1:0] m2sw40fca0wvnmy,
  input  ywhfwlbfro2dmuvf , 
  input  [5-1:0] nodrapn01yl1vxle30p,

  input  ex_g_cnadtiu1r9u,
  output orzasugx5h5pio22_,
  input  [64-1:0] dxwtzud_wfj8jqk0,
  input  [4 -1:0] gi8o690aydhqi8,
  input  zl1r9cfvuhltjq ,
  input  [5-1:0] dn074lh73rzchvrqzm8,


  output f71k3zhdtjavw19c52g45, 




  input  [31:0]           ij_sgq3rtvw2,
  input  [31:0]           k9jntnqwqp,



















  input  gc4b3kdcan6do88ta_,
  input  dk2xhkj77a,
  input  stlp3kak,
  input  gf33atgy,
  input  ru_wi
  );








  wire                         se2buoxmq91dbic3y2m5hu;  
  wire                         e9u0rtvt8jrygyc8s;  
  wire                         eyvp_wq1ero7byc8pxubqtg;
  wire                         g0gwombfdn5ycvw4m1vh7f95; 
  wire                         umtp4mg0svcx_tzytl9f2gx_9qa; 
  wire [32-1:0]   ave0oxjdt4lz6czd61woyw2yb; 
  wire                         hc665sbb0domfwj0scqo_bhyan0;   
  wire [64-1:0]        ehzuy3rj6cnownydmlhhqorz; 
  wire [8-1:0]     a8hb7l400suw5vjdy40x_cjbtdzv; 
  wire                         srz_pttv795yabd3rlohv25jpcoj;
  
  wire                         w9feuue3j76drwahit30vtv396w;
  wire                         caj02kz7j7ejw81vsf0fla;
  wire                         evt2fcz8mh_y8u4scgguyq287kcm;
  wire                         wrqq_2zdqd0x7l_8uyy75putmx;
  wire                         f9gyp2oa2mz_rqxqxrizc1l;
  wire [1:0]                   rn2r2g1hhe3zfa2usi0x_mw;
  wire                         gy3d5ed4dpwebmbht825jpu;
  wire [4 -1:0] fcfcmwdw40u0wskca41p_6qb7m3;
  
  
  

  wire  l_giy79jkzkxy7j  ;
  wire  cw9xa748nw    ;
  wire  x1huhi29x9mco   ;
  wire  fpo04urqz74     ;
  wire  a2i6e7_7    ;
  wire  cque110xwd150_ ;
  wire  m705cbtazx7y  ;
  wire  etp831o_vh94  ;
  wire  w3p1po3pu   ;
  wire  nxy2oljfg0lssc  ;
  wire  n2s7mr_zvl9k  ;
  wire  mzwwsw0h6m1  ;
  wire  lydg_n0cr655 ;
  wire  tb62wswspbytv ;
  wire  [64-1:0]      jttn_e63nm4n4lm9; 

  wire                         oa95jvzldxkjxnka5;
  wire [32-1:0]        hjbzyjew4g2fmth4l66ng8;
  wire                         dl59edtk0_9k5jd65gxp;
  wire                         unzbnfwje52jxr_9yt38_bmn;
  wire                         qtcuhd18j5hjtx41o9tjmv0cm434;
  wire                         srphqbnx3w67orxkuwvoz;
  wire                         jbju6a9hecf_f8kg2bsz4;
  wire                         w66c528fqa9qnfz1btjnm;



  
  wire                         qhvzepznvxpv9_wyiu767h7;
  wire                         lwjhzma3f8s38cp0iw7a471x;
  wire [64-1:0]        kcliouozy4gzxf4ji1d_1ug;
  wire [4 -1:0] t208_ksfx0p48awxbbi41vdc6k;
  wire                         p6887dnv76xwdpql2ru4c ;
  wire                         lkdi90h27rm6bstdc_lv43xs9hw;
  wire                         p1todm057e8_laqnquniw6y0rw6;
  wire                         uvbcza18x9h661vyy9t1uik595c;
  wire [64 -1:0]  ff37q45o11p27pc_tlfpgr8yspb0w;
  wire [64 -1:0]  bv8onmahmkg35l9opjmw5v1axpaj;
  wire                         d_arhdx13m6c57bz_fusjchynkad;
  wire                         vx75xcy7pymxftm_8zyk4pytv9kuyd;
  
  wire j2_lz0mpsxf4xotgqf1ngx;
  wire hcugdkhp9szims1nk8rhakn;
  wire dw2ygdedledlm7ps830qgbwonu; 
  wire ygvgcd3cyi2ipiz53hbsp;

  
  
  wire                                   vs6ryzcr0bwqs5so                ; 
  wire [32-1:0]                  j25ub196dc_agl8oovaex4               ; 
  wire                                   pi2nokcm8qf7och7l4g               ; 
  wire                                   c0i0hs5tz64_ce5f0z              ; 
  wire                                   dmzdczrqcueolg3dzufj_by5rmf         ; 
  wire                                   a1sqko6fok9qzpbtyuw0              ; 
  wire                                   bquohubxiv2rsayn62v              ; 
  wire                                   kqyojh1maxy0x834htg             ; 

  wire                                   refz65mt7g99f_cb9h                ;
  wire                                   e2rgt3d7pxx8bv6_w1v7                 ;
  wire                                   d6ltnbdw_4ll2                     ;
  wire                                   lmrvfbh6ipddvrrollz4_              ;
  wire                                   zh907qs92c1ixb_97gmdepk            ; 
  wire [27-1:0]      phofig8d5zd_8v9g8                   ; 
  wire [1:0]                             hey6uxy22wzzlom6mekyg2y            ; 
  wire                                   qerr94cedlotaj08239y                ; 
  wire [26-1:0]    js0ml55dtie8qenb4eoj2             ; 
  wire [64-1:0]                  ticm3jrqt6tjtf6                  ; 
  wire [64-1:0]                  hpaul9bznamp4qkl                  ; 
  wire                                   vq7jwn83uus_ac4s4ghf            ; 
  wire                                   gzh3us4_ux10aey                    ; 
  wire                                   np3fnkgbpsuf8nkgnf                ; 
  wire                                   hpk3eafyque5ubt_c62flnny           ; 
  wire [27-1:0]      sfezv1xz2ghvo8pkt                  ; 
  wire [1:0]                             vagaza053272juvmo59v8w20s           ; 
  wire                                   rzf45534z36ejq96260               ; 
  wire [26-1:0]    frzfsbt7hp3n4aj3zvvumnh0s            ; 
  wire [64-1:0]                  zkuxqezrmlhyyjjgx                 ; 
  wire [64-1:0]                  u3h5tvu1g2q93141j9o                 ; 
  wire                                   pjh0wad7t_5du3cync_0c           ; 
  wire                                   wmkgrgf631pbq                   ; 
  wire                                   oyq1p3qa2iffjuqns0jkgg               ; 
  wire                                   evji0n54bi8hm_n24uk853qw9c      ; 
  wire [27-1:0]      s9psy03yyyxh7qrmosmb1             ; 
  wire [1:0]                             sqkbogq1h4psprgoosl2lmrpj9_      ; 
  wire                                   n5gj_lxl9078ky9b2zawd0          ; 
  wire [26-1:0]    b0fkq6hghv6az5l_j1j2c12imdd6       ; 
  wire [64-1:0]                  argq10f3h723e0jtlrdbu53            ; 
  wire [64-1:0]                  e7iar94ylidlt25a9g9n            ; 
  wire                                   qj6kqe1holct34gfb0q9p9a04_alrzg      ; 
  wire                                   bmkssziw1_8am7ea6dv              ; 
  wire                                   xefc2nul9m648jueckdrui_l          ; 
  wire                                   c9k79dqw2z4f63_8lcp4w            ; 
  wire [26-1:0]    ly39gmn8_bufgxi162s47mj5md         ; 
  wire [20-1:0]         u6f8hwzstewuo7nl0iywamw              ; 
  wire                                   owio9cfz6lmpk7katn_gtlo9             ;
  wire                                   dna64e9sa3ona8c40stq             ;
  wire                                   yqonk7rjhe328d_deg1             ;
  wire                                   fvuwaqmgv_r72l8z4ys0lq59             ;
  wire                                   x5_495u23v2cqjqs7nx9m3s             ;
  wire                                   j9pnp242pb8iiimxe87y                ;
  wire                                   qvfjqeg7co1udtegoqx2t09jmc       ;
  wire                                   m6_yvtzjevmj_c4bel_9vu0kkk_t     ;
  wire                                   woq47beoqkpu1um82nv58l1u_hyj4      ;
  wire [26-1:0]    a1r66jlym5w100htq8lfn_o0rapdf5s   ;
  wire [20-1:0]         trt0bnwhmoe0r7apy2x_p9hltd;
  wire                                   wqjorkypks0nndgahingvyvil3dvqo;
  wire                                   obokll126527kg6wlw1t6vfh8;
  wire                                   msh4030y2dhqf78kyckys0c2ue0ic;
  wire                                   oebo4piph5o2byr1030bgmb0ye31c6;
  wire                                   tlmtrlht_1gsijvzms1twiewyym;
  wire                                   ez_fxjs3_wlsve__62ua9tqsfa6k89twfir;
  wire                                   p3nsxkqv6seglstz4ge77tdjcngbig0w30rq;
  wire                                   qjw2q0j88rjr42lautsqnca            ; 
  wire [26-1:0]    imkm56ujne9v4m6n08w1yf5622         ; 
  wire [20-1:0]         txk1r9aiq_7l2nkw101w_              ; 
  wire                                   ih4hmwugasiodbx5da9_40kx             ;
  wire                                   x5vjq7mshfwr0h3q514t7mhdt             ;
  wire                                   qrxtk7e03100_uwkx73sg7             ;
  wire                                   i7qiq2q9c6hbeful9qu9lb             ;
  wire                                   yr0s3skqk7cdqflsrbsxg9znu             ;
  wire                                   adqieke11qo0elfz93hlouwjc0       ;
  wire                                   w93gdpnnxuydy53eu0s9nxw7xdct7     ;

  wire                                   s47txxhzt1zertcfln5                 ;
  wire                                   w0s0l3_vvnnjgr_7cg2               ;

  wire                                   b0ry73kp6sc2;
  wire                                   hr64e6c3gy ;
  wire                                   cz1hh6af7xp2;
  wire [1:0]                             st2zalpx0uf; 
  wire                                   ni01kj42oob2x;
  wire                                   ah8kjlmvnaxzbi;
  wire                                   fkuqlh34r;
  wire [16 -1:0]           hnc10arn_rd;
  wire [20 -1:0]             b2ulqcjb;
  wire [1:0]                             w30ye15yns15;

  wire                                   vdtkg4_jnsbu0p8wqnasmncdouhwmk;
  wire                                   dll7vburbug9zho0oh3rpr0pnjnnh;
  wire [64-1:0]                  wqbvx_uqjrfzj8cjke712tpq;
  













  wire [64-1:0] dy_nwgv6;
  wire [64-1:0] f_ljupvj_wh;
  wire [64-1:0] v1tu43o;







  wire [5-1:0] f2x5pi_qvq5;
  wire [5-1:0] rw6_l_0bzu7h_k;
  wire [5-1:0] k0a54ytxmfbhg;
  wire [5-1:0] rig48lgqgq8oxt = f2x5pi_qvq5;   
  wire [5-1:0] zaub9z0lm4s93y = rw6_l_0bzu7h_k;   
  wire [5-1:0] j_69hsshtbv = k0a54ytxmfbhg;   
  wire [5-1:0] kd6v2vk601xpnm ;   



  wire sb8ax73d3ud = gy5zhpbrnl;
  wire f9_w27gbcq__ = qv70a7n8p;
  wire iq9sj_i8z1k712 = anlbkc8jny;






  wire dqyc8po_8fx = jjzotrbn & hw1_k1jmu;
  wire jdilf8e00vb3v8b5wy =  sb8ax73d3ud ; 
  wire knvph84tf1ry6cw3yr =  f9_w27gbcq__ ; 
  wire crn_7p36v3mpr  =  iq9sj_i8z1k712 ; 
  wire c8xzhxo1hdq9yc5_ = jdilf8e00vb3v8b5wy & dqyc8po_8fx; 
  wire u2l_1mg4um_jvsz_ = knvph84tf1ry6cw3yr & dqyc8po_8fx;
  wire bn4gs0qptrej1g = crn_7p36v3mpr & dqyc8po_8fx;
  wire [5-1:0] wf1tajpedkiof25 = cpt0qfwiz;
  wire [5-1:0] x16252ur82ajlgnoa = vf7a_1kae4zv5;
  wire [5-1:0] h9me0s065bzyb669 = djv9nstr;
  wire [5-1:0] o5r84zerdxtf;
  wire [5-1:0] muhxao8ez6o_4;
  wire [5-1:0] nosygh5mqqgj7g7;
  ux607_gnrl_dfflr #(5) t1ajzj4xsxst1u2njum4(c8xzhxo1hdq9yc5_, wf1tajpedkiof25, o5r84zerdxtf, gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(5) xxc6jnsjttv72ij5(u2l_1mg4um_jvsz_, x16252ur82ajlgnoa, muhxao8ez6o_4, gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(5) lyzatn8zi425mebdszp_7(bn4gs0qptrej1g, h9me0s065bzyb669, nosygh5mqqgj7g7, gf33atgy, ru_wi);

  assign f2x5pi_qvq5 = jdilf8e00vb3v8b5wy ? cpt0qfwiz : o5r84zerdxtf;
  assign rw6_l_0bzu7h_k = knvph84tf1ry6cw3yr ? vf7a_1kae4zv5 : muhxao8ez6o_4;
  assign k0a54ytxmfbhg = crn_7p36v3mpr  ? djv9nstr : nosygh5mqqgj7g7;

  wire rnx27onf2lbe;
  wire g_o2wra9n9s = k405wpjt;


  wire i7pubsxfsb4uys;
  wire [5-1:0] jc4yg1pkylr2gonwcd = bq9_5ksloh67_2ti;
  wire [5-1:0] nd3cgvec1pogf2 = qosgyc25p4fzq8b4;
  wire [5-1:0] f7crsrzernrwgmepy = cqk3fh13g1cxf9j;
  wire [5-1:0] pw085ct76po3c;
  wire kfz3mojvfh2fsfd;
  wire [48-1:0] g5usf8ixwjaxjs1m;  
  wire [64-1:0] pxhhgm9746n;
  wire nykwng_3anppxi  = epi4op2w5ban9o;
  wire shpynlimbt55rj4  = heqeu11d07lcg2ss;
  wire jycwup76klyed6d2  = exzr5we0sujvtby;
  wire fgm5kq4y725x6yylw = anvecdxcx1ouoa0;
  wire awld9ngcypgfxa = x240tjzbog6i9q;
  wire v5m66onlnmxeejfhn = uimia9sdhaq9x;

  wire d40y0va2l7xzj   ;
  wire [48-1:0] hhj5975j18r0n  ;


 wire wzcablvbov0zio = g_o2wra9n9s & (~rnx27onf2lbe);
 wire j5jswvt7ahm_iw0l4noh7hi = wzcablvbov0zio & nykwng_3anppxi & fgm5kq4y725x6yylw;
 wire kklg95ydii_hyz_wjg = wzcablvbov0zio & shpynlimbt55rj4 & awld9ngcypgfxa;
 wire gf1pz3n62zkjsykks7h92m = wzcablvbov0zio & jycwup76klyed6d2 & v5m66onlnmxeejfhn;
 wire zvnl8r316zxiqhn4avn3x = j5jswvt7ahm_iw0l4noh7hi & dqyc8po_8fx;
 wire hmakr66bx296ugqqe72 = kklg95ydii_hyz_wjg & dqyc8po_8fx;
 wire md4d9y8uf1q_udklshht = gf1pz3n62zkjsykks7h92m & dqyc8po_8fx;
 wire [5-1:0] xhv2ftbxji78ahyjyhulux = bq9_5ksloh67_2ti;
 wire [5-1:0] hnt2ut9n45ct3cbdgq4w = qosgyc25p4fzq8b4;
 wire [5-1:0] k_7iup5p8ivubmxl_yt = cqk3fh13g1cxf9j;
 wire [5-1:0] sd1q3796ad87z_81;
 wire [5-1:0] t1u2equ5qaj721ozxroou;
 wire [5-1:0] fzzthsme4xnzp1g7;
 ux607_gnrl_dfflr #(5) xtelriwli2rymfw_kmw_(zvnl8r316zxiqhn4avn3x, xhv2ftbxji78ahyjyhulux, sd1q3796ad87z_81, gf33atgy, ru_wi);
 ux607_gnrl_dfflr #(5) doojy862_8u69mdi_rg_nm0v(hmakr66bx296ugqqe72, hnt2ut9n45ct3cbdgq4w, t1u2equ5qaj721ozxroou, gf33atgy, ru_wi);
 ux607_gnrl_dfflr #(5) aw42v24_x83g0tc0m8fv(md4d9y8uf1q_udklshht, k_7iup5p8ivubmxl_yt, fzzthsme4xnzp1g7, gf33atgy, ru_wi);
 assign cjo14q6bim0c = j5jswvt7ahm_iw0l4noh7hi ? bq9_5ksloh67_2ti : sd1q3796ad87z_81;
 assign yqawr6m8r98vjx73 = kklg95ydii_hyz_wjg ? qosgyc25p4fzq8b4 : t1u2equ5qaj721ozxroou;
 assign wuzzw7m7hpf4p6q31 = gf1pz3n62zkjsykks7h92m ? cqk3fh13g1cxf9j : fzzthsme4xnzp1g7;




  wire                         u2a25670eeoaaxpdc;
  wire [64-1:0]        dl2wnjpp4e2270jy;
  wire [5-1:0] fy1at1kp6l7l_r5w__q;
  wire                         nruhqt4v8aa4ul498;
  wire [64-1:0]        sf3mcfi86e2vz;
  wire [5-1:0] j5zkfgic67jhz8;
  wire                         aw3rv1bswmks;
  wire [64-1:0]        etusjysf1bvjmp5;
  wire [5-1:0] u3fyvcviv3tk65gmcth;

  pkdsokaky2kt15iive heje9e9heregeo1z_uj(
    .rfe2lglwm   (ollg7),
    .w42_wd9um28vh (f2x5pi_qvq5),
    .ssjx8h5cj3q4ffem (rw6_l_0bzu7h_k),
    .rwby8vkzgm4y4r (k0a54ytxmfbhg),
    .vuv0917fanv19 (dy_nwgv6),
    .j2xzlc7dmxgmtn6kmk (f_ljupvj_wh),
    .tkxnzh2vh65vfutt3 (v1tu43o),

    .oxa8a6mj5          (l_imk5zs8ejjka),

    .j8mbnycgbc8k4exus50 (u2a25670eeoaaxpdc  ),
    .uup8_48koujjsde7s4 (fy1at1kp6l7l_r5w__q),
    .unb_5mvf3gc1403brsa (dl2wnjpp4e2270jy ),

    .nlxthgp55i6f26ozu4n (1'b0          ),
    .y9hqso2yg_rpfqu (64'h0 ),
    .bhxoyk3s_9ylb3 (5'h0 ),

    .ub63nbp2x73net910cs (aw3rv1bswmks  ),
    .u04hsk__lriad8ii (etusjysf1bvjmp5 ),
    .pi6em2fjks8g1zb87 (u3fyvcviv3tk65gmcth),

    .gc4b3kdcan6do88ta_     (gc4b3kdcan6do88ta_),
    .gf33atgy           (stlp3kak          ),
    .ru_wi         (ru_wi        ) 
  );




  wire fpwql5ik7_sp0;
  wire dwci8hbxok739;



  wire [19-1:0] eaxqugrf_ryu5rxxw41;
  wire tkm5u9dl8zav4;
  wire [64-1:0] t05leas4w4r;
  wire [32-1:0] zk9uk90j08ogqpn;
  wire mg0onistbzu9ys;
  wire g3btysb7vvv;
  wire yjgkn7vcv;
  wire b6cv9yeaga7hf;




  wire fqizcmmfg ;
  wire tbuacpjktio ;
  wire ciftsjs2bvaxns ;
  wire k_y4yq3crp_zqtg;


  wire vfye1vj155_k;
  wire vujduks2o30;
  wire y4zqru1tedm;
  wire q1coyps2cz7xe;
  wire sibtd2rf5j;
  wire hgvdw0qnels8;
  wire aiok9wht8yx8u6dz1e;
  wire [50-1:0] mg4yq4mui7ruja;
  wire [105-1:0] z8t7w6zr5woh649;
  wire oli3_udj80h6urj;
  wire m05tjqf24b1fabuu0e;
  wire rphjsg75001l2;

  wire ch8qv98q9xu469etyz8oj;
  wire [48-1:0]  zj0wqwminaxn;

  wire nnng_p6632p;
  wire jw1vgacy_r0vr;
  wire [64-1:0] bdhv0j4zhtx9nxmz;

  wire [15:0] ru3mfqrzh6 = nrebzehsuam ? j3oz8j2[31:16] : 16'h0;
  wire [15:0] q9933q2hmd = j3oz8j2[15:0];
  wire [32-1:0] k_pblo0 = {ru3mfqrzh6, q9933q2hmd};

  wire nt2l7qcrv0wofhii = y4zqru1tedm & zj0wqwminaxn[6:6];
  wire [64-1:0] n0b78w3x6yz3b = 
                                    (nt2l7qcrv0wofhii & ciftsjs2bvaxns & mg0onistbzu9ys) ? 32'h00000000 :
                                     dy_nwgv6;

  wire [64-1:0] zrhbyythja =  f_ljupvj_wh;



  wire                    werzz_4cg4m65i ;
  wire                    i5ogs4ipdqkwou0;
  wire                    qzdlalytscynhz1 ;



  jgz9v2pi3n5adi7j41 b2163wfvtrtbqnnjbc0fx (

    .qbsr1jytrqtsbk4ttb8nz(qbsr1jytrqtsbk4ttb8nz),

    .b0ry73kp6sc2  (b0ry73kp6sc2 ),
    .hr64e6c3gy   (hr64e6c3gy  ),
    .cz1hh6af7xp2  (cz1hh6af7xp2 ),

    .k0xug5g      (k_pblo0),
    .qhyq467foflgyn5y (qhyq467foflgyn5y), 
    .sa2f4h4xeakpfnunl (sa2f4h4xeakpfnunl), 
    .u2k4dyp52s_m      (u2k4dyp52s_m ),
    .djvj1e_      (djvj1e_ ),
    .bktu0z1mk56      (bktu0z1mk56 ),

    .s1woka0byzgo   (s1woka0byzgo),
    .al4xeg8mukgfg     (al4xeg8mukgfg  ),
    .piwiqvrjoq    (piwiqvrjoq ),
    .wi_dfzp70x09hm1m  (werzz_4cg4m65i   ),
    .jdyqycv3wdp2sgy(i5ogs4ipdqkwou0 ),

    .ld01d40_n3   (),
    .o8rwk067   (),
    .r1on2k03r  (),
    .gw7452ctd577  (),
    .b1roq8tr9r   (),
    .j_ku88w81rg   (),
    .ng_pudjzgnamv0es(),

    .jw1vgacy_r0vr   (jw1vgacy_r0vr),

    .t9xs6bqphiru  (x9cmkt53yq483z1),
    .ls1dudpc     (),
    .tzjssx03b     (cxmwxfttqy2t7ura   ),
    .cni2453cuofb     (b5wruck8tj9sa   ),
    .kt04okvuth    (bxentpryfwb3d  ),
    .kq9gup8pu2    (o2a43mjdbgea1  ),


    .rnx27onf2lbe     (rnx27onf2lbe),  
    .g_o2wra9n9s        (       ),
    .nykwng_3anppxi  (              ),
    .shpynlimbt55rj4  (              ),
    .jycwup76klyed6d2  (              ),
    .i7pubsxfsb4uys  (i7pubsxfsb4uys),
    .jc4yg1pkylr2gonwcd (              ),
    .nd3cgvec1pogf2 (              ),
    .f7crsrzernrwgmepy (              ),
    .pw085ct76po3c  (pw085ct76po3c),
    .g5usf8ixwjaxjs1m   (g5usf8ixwjaxjs1m),
    .pxhhgm9746n    (pxhhgm9746n ),
    .fgm5kq4y725x6yylw (              ),
    .awld9ngcypgfxa (              ),
    .v5m66onlnmxeejfhn (              ),
    .kfz3mojvfh2fsfd  (kfz3mojvfh2fsfd),
    .m05tjqf24b1fabuu0e (m05tjqf24b1fabuu0e),

    .d40y0va2l7xzj    (d40y0va2l7xzj    ),
    .hhj5975j18r0n  (hhj5975j18r0n  ),





    .mg0onistbzu9ys (mg0onistbzu9ys),
    .g3btysb7vvv (g3btysb7vvv),
    .yjgkn7vcv (yjgkn7vcv),
    .sb8ax73d3ud (         ),
    .f9_w27gbcq__ (         ),
    .b6cv9yeaga7hf (b6cv9yeaga7hf),
    .iq9sj_i8z1k712  (),
    .hgvdw0qnels8  (hgvdw0qnels8),

    .rig48lgqgq8oxt(          ),
    .zaub9z0lm4s93y(          ),

    .j_69hsshtbv(          ),
    .kd6v2vk601xpnm (kd6v2vk601xpnm),
    .t05leas4w4r   (t05leas4w4r),
    .fpwql5ik7_sp0  (fpwql5ik7_sp0),
    .dwci8hbxok739  (dwci8hbxok739),
    .zk9uk90j08ogqpn(zk9uk90j08ogqpn),
    .fqizcmmfg (fqizcmmfg ),
    .tbuacpjktio (tbuacpjktio ),
    .ciftsjs2bvaxns (ciftsjs2bvaxns ),

    .eaxqugrf_ryu5rxxw41(eaxqugrf_ryu5rxxw41),
    .tkm5u9dl8zav4  (tkm5u9dl8zav4  ),

    .z8t7w6zr5woh649   (z8t7w6zr5woh649),
    .mg4yq4mui7ruja   (mg4yq4mui7ruja),
    .sibtd2rf5j     (sibtd2rf5j  ),
    .vfye1vj155_k  (vfye1vj155_k),
    .vujduks2o30  (vujduks2o30),
    .y4zqru1tedm  (y4zqru1tedm),
    .q1coyps2cz7xe  (q1coyps2cz7xe),

    .qzdlalytscynhz1 (qzdlalytscynhz1),

    .oli3_udj80h6urj  (oli3_udj80h6urj),
    .rphjsg75001l2  (rphjsg75001l2),
    .ch8qv98q9xu469etyz8oj (ch8qv98q9xu469etyz8oj),
    .zj0wqwminaxn(zj0wqwminaxn),

    .nnng_p6632p    (nnng_p6632p   ),
    .bdhv0j4zhtx9nxmz (bdhv0j4zhtx9nxmz),
    .k_y4yq3crp_zqtg(k_y4yq3crp_zqtg) 
  );



  wire vvsvl34lm1_1h; 
  wire r_p2yyjhd3; 

  wire [4-1:0] hn_32518x9i;
  wire [64-1:0]    qpscc8xem;
  wire [64-1:0]    u3wdadynlf;
  wire [64-1:0]    igvq6tvqkm;
  wire [64-1:0]    xz5xffoimfam1;
  wire [64-1:0]    iaekulscp0d5;
  wire                     gkx4s0wv_05dt7e;
  wire [5-1:0] lnwarwpyiph_rhx;


  wire [64-1:0] u5115crirpno;



  wire                    qdh2itqlmn859kps6;
  wire                    g2515ltnbxvz;
  wire                    u8cs2vcqau77o ;
  wire                    k0tpiu_dns7fesh ;
  wire                    h9v5a720moqn805 ;
  wire                    q3l2pm3uzu4 ;
  wire                    dsff_1r8ibc2u1kl52;
  wire                    altukww2cr3  ;
  wire                    gosrdaw5huebw9  ;
  wire                    uf9szdd1w73  ;
  wire                    qh5uw_vgky8ctx9s ;
  wire                    ncr4iqrzig1xhs584u;
  wire                    g59aakolhtnl6vjex;












  wire [64-1:0]      y2ee2w8tps_6;



  wire                          o7wl_069n_sy5rue7;
  wire                          nt344pvhrf4_gj1h1pp;
  wire  [5-1:0] j2vhfgh92_ia2leet_11;
  wire  [5-1:0] o5j_0q84lvbq1m6zqcrttm;
  wire  [5-1:0] oxmshd1ilks70i3zxfapd;
  wire  [5-1:0] nu1oenmx9659cv65 ;
  wire                          gv5x7tbabwro1zc6cvwa ;
  wire                          t2qvskf77dx_qfcl1 ;
  wire                          j3iskguxr07s_auk4h ;
  wire                          bqrsuxkxg7wfhxfo3_k ;

  wire                          f136__ouz2d6kha2 ;
  wire                          ldzmdnb_744cs12l0t ;
  wire                          so92sz9arx155dg58 ;
  wire                          dqhqa5vyv4o5r73gsbmlg ;
  wire                          isjfto67rigtgkzl5 ;
  wire                          w9cz5plbg7bt3u34h6d_ ;
  wire                          c1a4qnyxrjj1h_g8  ;



  wire                          q_wc5085zblpey;
  wire                          srowfx3o2v3rl;
  wire                          od2labe2838d;
  wire                          nb3g7kcdyt7bwtvq;
  wire                          u4vwxxdwlql;
  wire [4-1:0]   ofxcqyaipegys;
  wire [4-1:0]   jyp69_3c6ce00h7e;


  wire                          ipoo1harz8;
  wire [4-1:0]   e8fbphi7t5pf39a9p;
    wire                          t1kvrmw3rk07cq   = ipoo1harz8;
    wire [4-1:0]   roif50sqz2l = e8fbphi7t5pf39a9p;

  wire [4-1:0]      otg3fn806ut;
  wire                          vi03qlql8tkd5    ;

  wire [64-1:0] zz7qeo73h2suy9k30jfzo;
  wire [4*8-1:0] m8yvt2y7rtjci4j6g1k0by;
  wire [7:0] kdi4n7teicbpfh90v5_hm;
  wire [2:0] ybptxmszcng89e3sisfytlxnl_j;
  wire ebpt710a8zup4xs8xzo;
  wire [2-1:0] mbghtxhocdjiarvwm96k8n5;
  wire [9-1:0]  md5rsuwww5y3iwkgy03x6;
  wire b9dlu6jwb4xgx25wfn5okd_7xyqlk;

  wire feq1g7m2cy1erl;
  wire qwcb6hcmvfqmf032z;
  wire [4-1:0] ppx8euepv0evvizd;
  wire f1yknbdsst7yvsgvm210;



  zu3cpta_6amki_tj3nyfxw7 ijvjeq924fk_weqrgde6awlw(
    .j2f1_e0en     (bktu0z1mk56),
    .aw82i964do     (u2k4dyp52s_m),
    .y8_gkxsfle     (djvj1e_),

    .x6eruzvd5     (bwjyqadn    ),
    .kw2010ymt1iz5   (1'b0  ),
    .yeo38qe8mley55  (1'b0 ),
    .rvfxw53dft5    (1'b0   ),
    .r6dop3ru22     (1'b1   ),
    .n6a0r_0zddzrme8 (n6a0r_0zddzrme8),
    .azll7rq5fab5ou (azll7rq5fab5ou),

    .coeuovgdaw1  (werzz_4cg4m65i  ),
    .o_gen1so7__xgr3pw2(i5ogs4ipdqkwou0),
    .gf33atgy(gf33atgy),
    .ru_wi(ru_wi)     
  );





  wire  qfspmfi47b5jx99i0, ngy4ipxc1vxym69lu  ;
  wire blu0a55bvxo3cmeyj = qfspmfi47b5jx99i0 | ngy4ipxc1vxym69lu;
  wire w1et7pt4n96m3703shs = blu0a55bvxo3cmeyj ;
  wire d9_s5e6qdqa7haet4s = ngy4ipxc1vxym69lu;
  wire bq9gnoi981qw397qkojrj = ngy4ipxc1vxym69lu;

  assign um28jgd2x4mbs = 1'b0;
  
  wire v_zbcmfxuliycnh;
  v3jar7rg0a6jqc jmu9tbv104qn9vd3(

  .r5hpbriny8m67sv9e_ylgo1 (r5hpbriny8m67sv9e_ylgo1),
  .dyl5g2vgrvy4mb3       (dyl5g2vgrvy4mb3),





  .vi03qlql8tkd5      (vi03qlql8tkd5),


  .p1oz3zlyx9z099ko                  (jjzotrbn), 
  .i7xpott8rcin                  (hw1_k1jmu), 
  .i4ph1cg8ey91ao                 (ipht6ss_sh6h),
  .v367rhzcrd1qq5y                 (vfye1vj155_k),
  .m6ow3ped_b3ynpgtz                 (vujduks2o30),
  .po8t3bdmxflhl2                 (y4zqru1tedm),
  .acploblvq3_mum6ni                 (q1coyps2cz7xe),
  .d5hyfhqo_lj0prgy                 (oli3_udj80h6urj),
  .pf_xchk7690b64ux                (rphjsg75001l2),
  .dg8l11o4gz7pp4nz6q                (ndn228hd1n2x),
  .l_w_v2dy7wxfnyy_ka5                (kwk_z0jwwa2r),
  .zrckh33wcln3qe0gwm                (fnbi_cp8jq6t9ropn),
  .nog5k2tkaj_                   (zj0wqwminaxn),


  .so8hgqibdpmm                  (mg0onistbzu9ys),
  .jyc3e55o28bdrj7ce                  (g3btysb7vvv),
  .y4er8_lympr8x7vr4                  (sb8ax73d3ud),
  .fxa5t2739h1y                  (f9_w27gbcq__),
  .pdyldj59mo6vg0bdw                 (rig48lgqgq8oxt),
  .dxnb4vitu85cv                 (zaub9z0lm4s93y),
  .xfxtnu32e4                    (n0b78w3x6yz3b),
  .bzyabkjyg5aufwj                    (zrhbyythja),
  .l2t6z9zsi2w0_zq                  (b6cv9yeaga7hf),

  .kshl17el0r504ln0s0                (hgvdw0qnels8),

  .jjab0msl5gufous                  (yjgkn7vcv),
  .ng2go_dzj8ezoh                  (iq9sj_i8z1k712),
  .y0sg1fz2ziwsp                 (j_69hsshtbv),
  .be99yq3n56                     (v1tu43o),


  .k1hmos4y13oq40h(3'b0),
  .ir18j9t6197l06(kd6v2vk601xpnm),
  .a1nhqrkfzavps(t05leas4w4r),
  .d0fq7icjv8j5ogee(32'b0),
  .ee8ig_qwdt           (bwjyqadn),
  .kn1fenl59sz01m7vnq2em_s  (binjv97px9r7dt04h0),
  .u_rd99v1d167myvqms9  (jt4l0g4njcsrt720n),
  .yauc7c8wjjqclo3tp       (o_d157fc5_l),
  .m_h2ikgwk1idzghe517   (oypxxr_e_rms7ai),
  .sjpycsle28a3pm_p       (s68_9qhgnb_o),
  .u9fj6h2fgqotisf      (m9cdnl05ykr_3p),
  .z2kxp5om4aw87pz8o18n1z6h (akh3h7anvh7892ugn),
  .vuxawlqfs_00v7_hzu3nxvoz  (ajl4tppx98ihuirj_mxih),
  .hyt20f5h_uwl66fhu4_      (qzdlalytscynhz1),
  .qmscup3rxdd9panua6h      (piwiqvrjoq),
  .odgwr675x09tn       (al4xeg8mukgfg ),
  .lzddtts2zym6c0cpur   (ryc6z1c7rmzrnlno),
  .i11dangz7fq7x35giy       (rhufxsnopy0n ),
  .zyh78crm605f5vguk       (wbhvg_1r9435 ),
  .p_cayjjoaokcjaec     (s1woka0byzgo),
  .ciy8of6we8nbld        (u2k4dyp52s_m  ),
  .dcpzocokm__mx7iua        (djvj1e_  ),
  .isem4fqob1u88i        (bktu0z1mk56  ),
  .rqmodrsg4hiv3yd (k_y4yq3crp_zqtg),
  .e6dhhsva7_jc3yex    (dwci8hbxok739),
  .m01780lmcvgmej7gv   (werzz_4cg4m65i   ),
  .vmc4uk3dtr_i3b6a1ojb (i5ogs4ipdqkwou0 ),

  .ssbpxp6oebc9u      (g_o2wra9n9s),
  .mp__ij57saap5pzjguck(nykwng_3anppxi),
  .bzxq5cchssdayz9w(shpynlimbt55rj4),
  .j35b4l1vciavqz_c8d(jycwup76klyed6d2),
  .q3fqrzgv4ce7343pb4(i7pubsxfsb4uys),
  .lou99zfk5t2fgui5tdozk(jc4yg1pkylr2gonwcd),
  .vx_07j3zzi0_m3lyq2tj(nd3cgvec1pogf2),
  .zo2kgt18lgbbaee80oq(f7crsrzernrwgmepy),
  .cez5fjfkhrstof7vn (pw085ct76po3c),
  .woaibn5hs0f9zh9obi(fgm5kq4y725x6yylw),
  .rczetx728pgbbuyhj(awld9ngcypgfxa),
  .l4y91rsecb8o3de_m(v5m66onlnmxeejfhn),
  .i90ggmn3seqiequ3ikr (kfz3mojvfh2fsfd ),

  .glf9eqlzf6ocu2fgv_jen              (tkm5u9dl8zav4   ),
  .fn921s9pkxbuyodk3cs              (v_zbcmfxuliycnh  ),



  .d3le01r9nrj56s4d(vvsvl34lm1_1h), 
  .awd7cj8qhsnpdq2i(r_p2yyjhd3),

  .mhnv1zj1t2xbsvq6pgtez4d(1'b0),
  .h76iv7j9x_gukyjc7q75qp_kags(1'b0),

  .fssz5redtt2z0j3bm                (qpscc8xem),
  .vahtdoye9yd23j                (u3wdadynlf),
  .tc85_x5h95y20zrlyv5                (igvq6tvqkm),


  .cqiq85nw82tognls5    (),
  .e8htsab8ol_n9_vmg55h(),
  .v8h7kn3z48bhc41oj0m              (gkx4s0wv_05dt7e),
  .s_ngsncbxs5sazdn09m2              (lnwarwpyiph_rhx),
  .tml6nm8cttakxkfl21                (u5115crirpno),
  .qjdagljhhzu7oqkdf8dt( ),
  .pj2f1w77r_add                 (y2ee2w8tps_6              ),
  .euzjqpru0y77ampkkzy_xt        (zz7qeo73h2suy9k30jfzo    ),
  .mizeob9j8ozttr2_5f1bf4zfgw0j       (m8yvt2y7rtjci4j6g1k0by),
  .kbdkmakcambtuegb3yt           (kdi4n7teicbpfh90v5_hm),
  .i6zm27hf33zy3u5g9qudq24sqm285    (ybptxmszcng89e3sisfytlxnl_j),  
  .hl3g_tq2rbkqa9ohkpb            (ebpt710a8zup4xs8xzo),
  .zrnrmtty0nzt9spsnhdcm1fcb        (mbghtxhocdjiarvwm96k8n5),
  .m9w2x58qenx6t_2bi2            (md5rsuwww5y3iwkgy03x6),
  .sw9yrs02t82mjdszv19xlcnijsm    (b9dlu6jwb4xgx25wfn5okd_7xyqlk),
  .ta29h0x4_ymr6ur6mk04               (hn_32518x9i            ),
  .lgm4pk95gcg3msfburvh            (qdh2itqlmn859kps6         ),
  .r9xo5zxa6yk5sahklgriapc            (g2515ltnbxvz         ),
  .qhr7po23q4sobg2liu8pg             (u8cs2vcqau77o          ),
  .fat5whs4wafix5rmfhm4837957         (k0tpiu_dns7fesh      ),
  .wtormxdkxhzy97pmh             (h9v5a720moqn805          ),
  .dskiex0swz5vysk4mc5             (q3l2pm3uzu4          ),
  .w313qpi6k9c_3uaxaj_ew           (dsff_1r8ibc2u1kl52        ),
  .hzx0lxqvh33f51vttk0y              (altukww2cr3           ),
  .vzwsikmnhz1uumkd9              (gosrdaw5huebw9           ),
  .vfq4rm5ouxjqvse7              (uf9szdd1w73           ),
  .p0q6b5s2pyhh9h5qc724n             (qh5uw_vgky8ctx9s          ),
  .m755tv316f55fgbeul39qh        (ncr4iqrzig1xhs584u   ),
  .bvwm3a9jzm7y_sjdaeqvzzvxeg      (g59aakolhtnl6vjex ),



  .hwu6b9ql3l7sw43wkk0lg          (1'b0),
  .a4rzfgrj8wj0hf3kl4wtn          (1'b0),
  .dp3lxnqfh_zuqs0qfwzb8(1'b0),
  .g5uxvsehmtgyorg3wb                 (otg3fn806ut),
  .jya9awf7h3oxy2ame3                 (o7wl_069n_sy5rue7),
  .gjbc27bxx6tkh_1w1               (nt344pvhrf4_gj1h1pp),
  .i9h3d3za76przvk_l70p              (dqhqa5vyv4o5r73gsbmlg),
  .euc_83pmnhwvr32xx              (isjfto67rigtgkzl5),
  .o2psmcgly2h0shgva5              (w9cz5plbg7bt3u34h6d_),
  .f9fubli1q2_q74eh               (c1a4qnyxrjj1h_g8 ), 
  .rev7x95ee0q6067               (gv5x7tbabwro1zc6cvwa), 
  .bpr67a65mrtg6l5byk3               (t2qvskf77dx_qfcl1), 
  .qe_d8g8bvqcuzvaepz               (j3iskguxr07s_auk4h), 
  .l56hg65h6fdq8htrj6gb               (bqrsuxkxg7wfhxfo3_k), 

  .hrlh00uvgxvc0v3fhap               (f136__ouz2d6kha2), 
  .xnnfhu8lpo04_jagyvmf               (ldzmdnb_744cs12l0t), 
  .keve1s8kiyssv8a               (so92sz9arx155dg58), 


  .fnkzuyagjhoinc95_              (j2vhfgh92_ia2leet_11),
  .x70ugsspg9qc0ccmj              (o5j_0q84lvbq1m6zqcrttm),
  .bhpc3d1wahnkux0bil5x              (oxmshd1ilks70i3zxfapd),
  .wtrlpn7minfboagr               (nu1oenmx9659cv65 ),
  .feq1g7m2cy1erl(feq1g7m2cy1erl),

  .gf33atgy             (gf33atgy  ),
  .ru_wi           (ru_wi) 
  );

  wire alu_cmt_wfi;
  wire j39tby_g7kqga33w_m;

  wire                         s_7qgktcx5l9b;
  wire                         swk0us69_ctq2k;
  wire                         zcqvodebks4c; 
  wire                         eru3qosawo7xqc6t999;
  wire                         j29miwazgbxlk8;
  wire                         wsvr7r5n5ep12y; 
  wire                         i6zt9kqe09i5ky; 
  wire [5-1:0] ybf0zo9v_845pqb_jh; 
  wire [5-1:0] cw3uprz8e2rwau3z7; 
  wire [5-1:0] bsnlk54ub6j_e7; 

  wire                         q58rcdx67tyrer; 
  wire                         c4juuyd55lxion9c; 
  wire [5-1:0] tk22_ghwl49rxxdnop; 
  wire                         keta7gjvl7x; 
  wire                         no1k1_uyge8hlp; 
  wire                         xg63_va9bynd285dre; 
  wire [5-1:0] mwzhu7wrbq1rkp; 
  wire                         s1j5549fqdsj5ad; 
  wire                         msqwr_9vjwohg; 
  wire                         onnke16xcq5904dt; 
  wire [5-1:0] fy0rb852ky8dy1; 
  wire                         qgpl_3pohcjc3g; 
  wire                         kf18wkamz8k9bxuv2j; 
  wire                         w5151c0ak9j8c; 
  wire [5-1:0] u0oho0bfx9igpi; 

  wire m631c388smkc86tlvjo8cy0euyc,gose7syxzsxbsjpxu9gf46ryn,xltf9w3ak66b70kftwbyhk8hfkvrk, qd5sbh8mupp_n4y95vo;
  wire [4-1:0] hl8tx_5fn5baqsm5i614qe_, ydctapy4pueuwk6n3mwwodl2o, v5654pk52c83hd4wif_iicjko, fs6jojwsl0l32t7brm38vh;
  wire [64-1:0] s7vgjm2azmcc3uzzdc_7;

  wire [64-1:0] jwwku_el5h5h2lx6e0kyi;




  wire                          ua_r8723rm_0699y9ue0qself  ;
  wire  [4 -1:0] rlwzlq3wmb1t76we1pgot2d6_   ;
  
  wire                          boie2le90zg6moigey_xh5kjc6  ;
  wire  [4 -1:0] jpa3mq_tg3w9jebkjw0qy4zhw   ;
  
  wire                          vn7agcnzu58a7jbm9n9em4kadk_  ;
  wire  [4 -1:0] ec2k88gmpr185bkl8ndglqu_p6l3   ;
  
  wire                          yqlpqui4nfbe0t93srqmvngkzf4y1  ;
  wire  [4 -1:0] n2nv4gollbb6vbo938tfa19gk   ;

  wire                         iy6jwb45n967lh; 
  wire                         nv4qt_e1adenv0c; 
  wire [5-1:0] z8h5zyhj54howg; 
  wire                         f28m69gb9k8l_ic;

  wire                     e45zjh64jxwnli64ak;
  wire [4-1:0] dg8pvkc6n2uz2w2f;
  wire                     p1jdw9loxkz60taq_vkp_3;
  wire [4-1:0] eo5skx1ygvzuasbjgnyl ;


  wire woon4h3ivznl_qiu7i_9;
  wire                     a42c0ps3vi3,h5i09w3ul0070, srr68v2d6ti;
  wire [4-1:0] p7165rjkv,il76519zb__bx,a2q31s2sx9u1;




  wire kf2bfg0y804sefov7qwk95xq;
  wire [4-1:0] u9jwgutri3owj857elesn;



 moqpszi6cm8qllh02c2ny2 zuwetofs7yg8b5h12w5w2ml(
  .jfb7utzuy3zdlp(blu0a55bvxo3cmeyj),


  .z4423w2ovxgs284(o7wl_069n_sy5rue7), 
  .s9k46re7yyb4d9(nt344pvhrf4_gj1h1pp), 

  .l_clnlob7ji8v9527(a42c0ps3vi3),              
  .pnc251fe9pp3tm(kf2bfg0y804sefov7qwk95xq), 
  .h4sfadnxw7z3wz14(srr68v2d6ti),              
  .cpi07x9cy64pn2(p7165rjkv),              
  .eyd9fc4vjxutcl(u9jwgutri3owj857elesn),   
  .pyhxgdg6s29imj(a2q31s2sx9u1),              





  .a_rhsk184ulq9ofyz   (m631c388smkc86tlvjo8cy0euyc),
  .radwr7skyhm3jqso5    (hl8tx_5fn5baqsm5i614qe_),
  .ovpwjtytlapia4s3cl   (gose7syxzsxbsjpxu9gf46ryn),
  .zdid44qi3bv7q4phl    (ydctapy4pueuwk6n3mwwodl2o),
  .uo331eh1sm8wclmxid   (xltf9w3ak66b70kftwbyhk8hfkvrk),
  .lgrrvklyk4mm3aai    (v5654pk52c83hd4wif_iicjko),
  .aseeilkazdwwcb4raoo2   (1'b0),
  .ijxk119_taxeoqx0n    (4'h0),
  .d67xmgrcefvmtl4jvxtz   (ua_r8723rm_0699y9ue0qself),
  .brw5ihk9eaoddaefi7    (rlwzlq3wmb1t76we1pgot2d6_),  
  .kgrl1ycpn2xb_uhommxp   (boie2le90zg6moigey_xh5kjc6),
  .spknpgo66_t6t3dm__y    (jpa3mq_tg3w9jebkjw0qy4zhw),  
  .dj75s2vvoi93lk6c1i   (vn7agcnzu58a7jbm9n9em4kadk_),
  .ql612i235fqhavkhdu    (ec2k88gmpr185bkl8ndglqu_p6l3),
  .gawf4cwltls4ro8y_u   (yqlpqui4nfbe0t93srqmvngkzf4y1),
  .przse28gs3o6cuvfp21u    (n2nv4gollbb6vbo938tfa19gk),

  .rz544x9yj6wtz        (qd5sbh8mupp_n4y95vo), 
  .nkffqtpacz_8         (fs6jojwsl0l32t7brm38vh ),

  .lr9ry0wds3k88rvde7n  (f1yknbdsst7yvsgvm210),
  .smjqotzwkn9j4hf2ev_     (ppx8euepv0evvizd),


  .ipht6ss_sh6h           (ipht6ss_sh6h    ),
  .sbtst18g6wurw5m36lm8 (woon4h3ivznl_qiu7i_9),


  .qomzw_wq7v_mblz0qrfi  (swk0us69_ctq2k),
  .f015ahr7wg2fbe5_c5ja8(j29miwazgbxlk8),
  .g_sda8atgrsb3n64a1e(cw3uprz8e2rwau3z7),
  .r3d0cws3w3xmt0koa6l6g5  (s_7qgktcx5l9b),
  .yzu_ab6e_rylfgno7k0o2(eru3qosawo7xqc6t999),
  .ih20zj50pzg1yxubdakxiz(ybf0zo9v_845pqb_jh),
  .k9fd4y9sg2l8f8pi29mz  (zcqvodebks4c),
  .jcs6ikpya0beppu6gdyf(wsvr7r5n5ep12y),
  .do0utstzhn7g1d7unzt(i6zt9kqe09i5ky),
  .jenm8icl2nmc7a1huf5(bsnlk54ub6j_e7),
  .llha0lc4h8ie3t0l8  (             ),
  .g97p2rs03luvt0no8_ksk(               ),
  .mosdlr9l78vgfsp3tj1(               ),
  .t9le19upn_tsza2pzh3zii  (keta7gjvl7x),
  .ip8580r8cp1_26jkauyh1wb(no1k1_uyge8hlp),
  .x1k7b9da53adlb0frcz(mwzhu7wrbq1rkp),
  .zjz6klk8496qrc03ps2snhs(xg63_va9bynd285dre),
  .hv33acidoo0f1j4kpbs  (s1j5549fqdsj5ad),
  .j1otk5cqg9j9l3e8ynv(msqwr_9vjwohg),
  .ky4jzzww3o0e66ldnngw1p(fy0rb852ky8dy1),
  .xkeclsgck5wllhwobaopvb0(onnke16xcq5904dt),
  .vpst0pbni2odvl7nr  (qgpl_3pohcjc3g),
  .dd92276i_tlq259bo27zu(kf18wkamz8k9bxuv2j),
  .zv9jo3fw_4ik299ra2irk87(u0oho0bfx9igpi),
  .alnssn8w7d9iksq1ou7y2u(w5151c0ak9j8c),
  .e5fsovqfl70bx4m4ahb3o  (q58rcdx67tyrer  ),
  .nlb0f26rp9onx17ui5yzy(c4juuyd55lxion9c),
  .irsej5jxvp566dv071e6(tk22_ghwl49rxxdnop),

  .hh0mpxxw3c00cet       (iy6jwb45n967lh  ),
  .k1rpfwk8imnpek5     (nv4qt_e1adenv0c),
  .kayddlyy2ps8dzeq46a     (z8h5zyhj54howg),
  .t7m_v9aew2ud1e0u     (f28m69gb9k8l_ic),



  .gy5zhpbrnl      (gv5x7tbabwro1zc6cvwa ),
  .qv70a7n8p      (t2qvskf77dx_qfcl1 ),
  .ojbpo5z6urt      (bqrsuxkxg7wfhxfo3_k ),
  .cpt0qfwiz     (j2vhfgh92_ia2leet_11),
  .vf7a_1kae4zv5     (o5j_0q84lvbq1m6zqcrttm),
  .fhhe7189lmum      (nu1oenmx9659cv65 ),



  .cp7yy8bv2o8n     (dqhqa5vyv4o5r73gsbmlg),
  .ypmn53drey     (isjfto67rigtgkzl5),
  .msz_o10r_pkr     (w9cz5plbg7bt3u34h6d_),
  .q7qac2db3cbk      (c1a4qnyxrjj1h_g8 ),
  .yrmykp4o9t      (j3iskguxr07s_auk4h ),
  .rqj15_sdahil     (oxmshd1ilks70i3zxfapd),


  .zzxn5x18ahgk4     (otg3fn806ut), 



  .i0fdxue89ury      (q_wc5085zblpey  ),
  .z4ufug6cvdodh      (srowfx3o2v3rl  ),
  .kbmj0dq2hvlwx78s    (ofxcqyaipegys),
  .rod5c8pxpam5dt9n9y    (jyp69_3c6ce00h7e),

  .zuht4f9qjrazipld4u     (od2labe2838d ),
  .g4qik0dwtex1gpiep     (nb3g7kcdyt7bwtvq ),
  .f__fcmmb1thlj     (u4vwxxdwlql ),
  .vt96ugjl7qf4rqnj3      (ipoo1harz8  ),
  .xu91lmfwk_nbjrz_    (e8fbphi7t5pf39a9p),




  .skcjh3xhs73ucsbh77 (vi03qlql8tkd5 ),
  .s9kw_2m8ozw73_mbk1o0o  (),

  .gf33atgy          (gf33atgy  ),
  .ru_wi        (ru_wi)
  );





  















  wire [3-1:0] phk590vi2;





  wire ngiuqj2j6rsgfaeu27;
  wire ka4_ngr35vo6rrkp72;
  wire [5-1:0] jhes_c10xw065fcx;
  wire zc9t_vib9_fw44d;
  wire cwmxezrc3jv6hzxcfc;
  wire uig3ujuyq0_61kqb;
  wire xc2becmsn4fcniw6ks;


  wire ap889z2q8jbzn4dhurkzl;
  wire [64-1:0] y_jjs1fut37ilha91qtxkacsoxy;  
  wire rnodgdrxyr_tulm0nnnign;
  wire t0o4cn_ndv2lmnp;
  wire aa5a1tnclwe351p5ujs;
  wire [64-1:0] my5_v4hhb7oc51;
  wire [32-1:0] lmv45fhtl015bg;
  wire [64-1:0]    yd4wqg2e0i386ccq6y9;
  wire tv3_4qrynvnaoy4riz;
  wire uv_3uzx5ti04u5nd;      
  wire [31:0] ne5matgyfjvw3elazxt7p;
  wire y_gvnr7uidhcof1;
  wire zh_0_4wrffapmbs;
  wire nrze6rcjz4m65z;
  wire cjxy_cr6jzz17mr8 ;
  wire g0ovdu1w9dcoqg ;
  wire uxdt29u4dd96ukc ;
  wire r_cdggxn_7syt0g;
  wire uvw8h6lqr2ou0;
  wire cmv9vkluc86swnlc;
  wire rwip45nhuhbz2jkd4;
  wire x3r6u6q7ck5ud8wbii;
  wire p0ga7mahvd8zjma;
  wire hlxcm16byj04fp0;
  wire o4lqcf45nah3boccbw;
  wire alu_cmt_ifu_misalgn;
  wire qjg3a6detqucp4byrgs;
  wire qn6g68ul7q8pz3pvopdmh0m;
  wire [64-1:0] co8g52huetu0l9justjw5wcy19yi;
  wire ihmezohdr7mg9_blli7;

  wire oozkxp7aywu4l0hz73uedbtyiad;
  wire kxmzp6o3alj05dfq9d_e8ci;
  wire d2gcdo57ra3yxudimcwal0;
  wire ob__kc7kdtjxp74ajo7ql548o;
  wire v85ovm_7gp20oi4vj;
  wire j5wtbhk36xx9j2h1kgsniu9p0d9xzj ;
  wire qh0m9d6yrl5kb_1vvecw1kb1wrbm ;
  wire kihyrfzcb87yz3qnxq7c0o11at5u ;
  wire ho49hpl6ijpiop4thzf8rh6apio4u ;
  wire wk2sssl74c1xyhbm7pf29qtbpws1 ;
  wire vxcgun4z0ztx7nmvm;
  wire fq2y4oplmud5drf9s;










  wire rb050tnl;
  wire a94vd35etec4;
  wire el7_p8jit09;
  wire [12-1:0] e1go3iu;

  wire [64-1:0] l9erxxpnphqd26vg9;
  wire [64-1:0] hig2gwwbeuhnt65xrp;
  wire [64-1:0] z0yhjfv_e0yaa2r;
  wire [64-1:0] guuvp01vkcryglsu1p3;
  wire [64-1:0] vf5xcr67bqhzlo43_;

  wire [64-1:0] bj7h5jqg66r51jxki6emra;
  wire [64-1:0] zmfo8cca_77pc;

  wire [64-1:0] vmx1fh4kmh4c;

  wire v35y3qnk7mx3l1695;

  wire af5qc04tmn51e4u2h1z;

  wire ya8t4ev_aidf0t0x4or;






  wire r0s7d8cr68i2qs1z;
  wire kakelc68be0x7tdm9b9o;
  wire j3j1czgoam48vhs8auo;
  wire gm1r5itc44uxw_y0_msk;


  wire [64-1:0] p6rw9no76a3m;
  wire [64-1:0] vyxop00ua6vr;

  wire tywculgjyor8ndw   ;

  wire [64-1:0]  pldoasxyzlvx2;
  wire [64-1:0] tvh1llq2i3_y;
  wire [64-1:0]  bde41te346q515l;
  wire z1cj655u31   ;
  wire lhu2z948o3n   ;

  wire exltui35irvvmodu205vw;
  
  
  wire [64-1:0] nb3w1rq_ny95rvrt;
  wire [4-1:0] p_yx415so7q1vohijb;
  

  wire [64-1:0]    mne0dg23_1aal06pio ,em0guzjh3x0tokxd ;
  wire [4-1:0] pc67uztpd_zg6bsal,hno6u0yd_gjy_1t;

  wire [64-1:0] onacehe6tcgr,pv44129rj0uy831j6;
  wire [64-1:0] tyvyxz0mf,iaejzw1j2jb5i,aucihtckush;

  wire [64-1:0] oajzut537ryb591kzk,qos_22gbinvor4;

  wire [64-1:0] jwbql4ta0c;
  wire [32-1:0] kmfvezt2;
  wire qw6ymq0u4qknlwh,td_th3xz1iyqn_w,e25k01aox4_;
  wire [5-1:0] pdwodu8jbockhftk7;
  wire bwd5a_yj_liikyo,piiqrjby8_d9dndhct,b7fov0er1gnx,xyq4s_ubn1sx2s;
  wire o8rffdg1904azl0q,f0ziihie9il3138m;
  wire gldc_bv5wpppiij9;
  wire ljghmx9gec8jr0of;
  wire i6yx610m2nd7razu,luf9wadz1xvpbt,r8b6cghj00gkt7, rdce2xlm_syu,zcl5hta0nld, x882ucszl6qqk9m7,zlp9p2qtwrt0ra6c7,yd1xmujxb33j01a4c;
  wire ohftngf40mc7275vq;
  wire y3lf5lq_1tfm1iea;
  wire hv3n9x664ena;
  wire fa9nldm69zre__ccuu82h,jfnkyxema4_sqj5v2v;
  wire [4-1:0] omler2igyskatx;
  wire k_u427htf3nny,snxyhe6q4j0ik6is,di_rao90w5qbjlfn9,r43_rk2c1l4t;

  wire s2mopc8npltdcmohj94  ;
  wire ab20niin2uxlfv9w5s5n7y;

  wire                           lvamcxldxlbi7k3r;
  wire                           c_vdpq9m03rq493zpv2165d3;
  wire [50-1:0] rcp57t3vlm6czu6;
  wire [105-1:0] ja6yz91tkse7r9tt;
  wire ho405be3bp1ma;
  wire t4zsjo_uj3n_m5;
  
  wire p_gj56fnt4qky4n6sxai;
  wire pjz1nevm60h9ihnmunx4;
  wire [48-1:0] ytygj4ti9khaqpbhp;  
  wire [64-1:0] d9hqn06qm44jqmxo;
  wire hpf6iii62xdb170ho7ax;
  wire ckkfhtew3eup3984z;
  wire dved_rrjqsz_ib5rx8;

  wire                           ob602_qjqak28zc1l;
  wire [48-1:0] hu2q59l06nvqg7i7f;  

  wire o99cbvjf8lyjdj,y6tqh4z7ck7gj;
  wire kzdc2z8f1n1qrac7;
  wire [48-1:0]  vqp0990pwh3u9u4f;
  wire                                  fq4r9kho3s5rkyx;
  wire [19-1:0] b1_o25pwqim0zl2p159psk;
  wire  w0p_8cae4cqs_1hdeoydtp,g7rjoc9tw3_k7r1i21ghnsfcv;
  wire  hncm6yp50zjrhz9dcp1t1q,g_wqbz93wfi5bmx7bczdub7;
  wire                           yh8eetxf0xs392  ;
  wire                           gjfmlxjpnnka6o8odi  ;
  wire                           mbwb4j_f4iygi4phniwt  ;
  wire                           t8qh_jt867ifbzdy0  ;
  wire [4-1:0]    a6eyass0uv3sh81xwu;
  wire [4-1:0]    zhaca_k1wq3sy5wznci2pu; 
  wire [4-1:0]    l276zv1sj136kk9s9_unb3; 
  wire                           g_cuqgaizsk_nq6fwir1_ ;
  wire                           rrubg3ioxxvdto3bjmpfsy ;
  wire                           if5n6cmdrvnn2c0vt09 ;


  assign  aiok9wht8yx8u6dz1e = 
                              (sibtd2rf5j & mg4yq4mui7ruja[26])
                             & (lvamcxldxlbi7k3r & rcp57t3vlm6czu6[26])
                             & (kzdc2z8f1n1qrac7 & iq9sj_i8z1k712)
                             & (pdwodu8jbockhftk7 == kd6v2vk601xpnm)
                             ;


  wire [64-1:0]    jz2qz87howt08ld8lq    ;
  wire  [64-1:0] ksgamvgvgr9n02_txmv    ;
  wire                      lgs2ndps7oi98rleg8tshcz;
  wire                      y9bk3uc02upz;

  wire jol0q6b5zk9uuu_  = gldc_bv5wpppiij9 & (gjfmlxjpnnka6o8odi 
                                    | mbwb4j_f4iygi4phniwt
                                    | t8qh_jt867ifbzdy0
                                     );







  wire gkfhdl1lvs93nq2q = 
                       ((k_u427htf3nny | di_rao90w5qbjlfn9 ) & jol0q6b5zk9uuu_) 
                     | (y9bk3uc02upz)
                     | (r43_rk2c1l4t)
                     | (fq4r9kho3s5rkyx)
                     | (lvamcxldxlbi7k3r)
                     ; 
  wire jvi2i2xkdm88aoes = 
                      (k_u427htf3nny & (~y9bk3uc02upz) & (~jol0q6b5zk9uuu_))
                    | (di_rao90w5qbjlfn9 & (~y9bk3uc02upz) & (~jol0q6b5zk9uuu_))
                    | (snxyhe6q4j0ik6is & (~gjfmlxjpnnka6o8odi))
                     ;






  wire hnsixpix0gzu  = di_rao90w5qbjlfn9 & jvi2i2xkdm88aoes;
  wire a6qybr3pioqo0 = di_rao90w5qbjlfn9 & gkfhdl1lvs93nq2q;

  wire bjqlln4lucs2dyr;
  wire icczfaorqi6bmvsm5c4h,o_adoo65svxjvftm_rm3,evh7l6yf2zeh1opg8dw;
  wire                                lbuuy3oqfy7m98dnu6x6;
  wire                                k48o66po4ld1pl217myx5me3;
  wire [50-1:0] rj9754hija256ughfk96zd;
  wire [105-1:0]   ai272s0_wt92lhlok1_j2;
  wire r7y76nl0xxu4lp4 = (jvi2i2xkdm88aoes & k_u427htf3nny); 





  wire n7xyejmco0cd85m_d = ((~w0p_8cae4cqs_1hdeoydtp) & icczfaorqi6bmvsm5c4h);
  wire flxli77po8atcjwdr = 1'b1;


  wire                     lkvz9_caztnpkd5y1a,dvloyy6lickuq8759jcfc6 ;  
  wire [64-1:0] du9nxa6qo7knx2et1gw6, a9rvmf7a9nbie6nd923;
  wire [4*8-1:0] qrodgqtao6oexta13898,q7iyngsmbckvi2tht2wb5nh,elfo368_wilpagxfb_udyc10aej;
  wire [7:0]                 s4ec4uwf6ke9r_tpu    ,mq09q0m1l74z182ajkt2udd    ,h33etngddojmz59z88a1yv3    ;
  wire [2:0]                 o8s3z5xdvprqa0193p0    ,xsziw9gaor0xrlm1hvlpjr    ,qbwq6loiooi7x8oz3mm    ;
  wire kxcwjr8ri3x86f, reu5ooijp0czeggc974, qcs_9_0j844qh49kucr_8;
  wire b6p6azv95fkv2o7od5rkww9t, blw41o7zqxmgmztc9cwl593q4;
  wire b81kg80kxviv6w2l2dt8qq, jxknblho9wokk6irza7q48k6h;
  wire [2-1:0] crpiujipdzd_h3djv_bjup, m5mjr032v1z_erq3mxi07t3v, vmcutkgts6eafpyi257frl0pq;
  wire [9-1:0] sh7px5ghy0tmin8 , kccav9va65o92d7d9d    , nmn1jadde_4_xom6aqb    ;
  wire h_iyw8puc0v6p12hca799v99;

  wire                     r9hdxtws4mibgldl,jf9ko0etxomcrj25,i7qg9zxylz7rpfw286 ;
  wire                     tcveomov4rt0zai5ns;
  wire [4-1:0] nlbav8h239dt2a   ;
  wire [64-1:0]    rwtwoy92pmk4i    ;












  wire                           tb198r6lzk1sr77g4         ;
  wire                           abn9qjx8er38bt0stedss         ;
  wire                           nz4yhqimnsh10c6gso429         ;
  wire                           e0eyarvfj_jnbe           ;
  wire dd8pb3i1ec_uv5  ;
  wire s62ahm8e0we20r;
  qy_752rpwt4qqgs1gejira_te o61okcsx2t8btek447pam71bv (
    .j2f1_e0en      (zcl5hta0nld),
    .aw82i964do      (rdce2xlm_syu), 
    .y8_gkxsfle      (y3lf5lq_1tfm1iea), 
    .azll7rq5fab5ou  (azll7rq5fab5ou   ),
    .dd8pb3i1ec_uv5  (dd8pb3i1ec_uv5  ),
    .s62ahm8e0we20r(s62ahm8e0we20r) 
  );

  assign nz4yhqimnsh10c6gso429 = (dd8pb3i1ec_uv5 | s62ahm8e0we20r) & (tb198r6lzk1sr77g4 | abn9qjx8er38bt0stedss); 

  assign e0eyarvfj_jnbe = ~zcl5hta0nld & t5trf35s8vy & (tb198r6lzk1sr77g4 | abn9qjx8er38bt0stedss);    


  wire uys2_c7rmnm5gjf6t;



  wire h41082ijgnoh480fx5t;
  wire e0xd37xbhk4bxmxa9_93qr;
  wire gsbir68u7ok8gu2xesw0zek;

  wire vcn_k11zjsoeq1mbk6c7hfmmtm = (e0xd37xbhk4bxmxa9_93qr & tb198r6lzk1sr77g4) | (gsbir68u7ok8gu2xesw0zek & abn9qjx8er38bt0stedss) | uys2_c7rmnm5gjf6t;






  assign o8rffdg1904azl0q     = gldc_bv5wpppiij9 & (~e9u0rtvt8jrygyc8s) & (~nz4yhqimnsh10c6gso429) & (~e0eyarvfj_jnbe) & (~e2rgt3d7pxx8bv6_w1v7) & (~vcn_k11zjsoeq1mbk6c7hfmmtm);
  assign ljghmx9gec8jr0of = f0ziihie9il3138m     & (~e9u0rtvt8jrygyc8s) & (~nz4yhqimnsh10c6gso429) & (~e0eyarvfj_jnbe) & (~e2rgt3d7pxx8bv6_w1v7) & (~vcn_k11zjsoeq1mbk6c7hfmmtm);


b0gv4gv3sqckul0vbemwxr #(
  .gdctpuyrfi_b (0),
  .l_7qc0w_2x6i(1),
  .t5462hhws9i6ynbxi(0)
  )x28em0c_brupbhar4un_vhc(
  .cu1owrury8wsed               (nlbav8h239dt2a           ),
  .mt1z8r_sz               (pc67uztpd_zg6bsal       ),
  .uc9k3lw_iehx               (fs6jojwsl0l32t7brm38vh   ),
  .radwr7skyhm3jqso5         (ydtm1yuxqj7fmxvqc    ),
  .zdid44qi3bv7q4phl         ({4{1'b0}}  ),
  .x4owqbu74zh_xxr         (eo5skx1ygvzuasbjgnyl    ),

  .b43m7n67rav8he           (r9hdxtws4mibgldl      ),
  .qcutfgh43gov5u4urt           (jf9ko0etxomcrj25  ),
  .s73raoa0ilom1wyi           (qd5sbh8mupp_n4y95vo  ),
  .dnwb40nhmse7rcj0epzjo     (vz63qkw5s3m8urb9       ),
  .omeribg0gbgvpn78urilv_a     (1'b0),
  .jxogr1vy8jotyh8ivd2u     (p1jdw9loxkz60taq_vkp_3    ),

  .kl8zh4diafqs                (rwtwoy92pmk4i            ), 
  .jiartjoiycj2                (mne0dg23_1aal06pio        ), 
  .dtypmpwq1q2j                (s7vgjm2azmcc3uzzdc_7   ), 
  .uwl7jm0d1lv0xpo            (r7y76nl0xxu4lp4 ), 
  .u2l80pdclhyu1bl            (n7xyejmco0cd85m_d ), 
  .uamf3ccv7ouhi18            (1'b1        ), 

  .pkw60eo867gghh          (iojqlhtwx45_siz     ), 
  .strg8286lgex8p4_0m          ({64{1'b0}} ), 
  .avpvrch0prpui67          (jwwku_el5h5h2lx6e0kyi  ), 


  .lot9xvzuqrd5jm0scdx5t       (m8yvt2y7rtjci4j6g1k0by   ),
  .mn3tic51ckga0gc           (kdi4n7teicbpfh90v5_hm       ),
  .k0be3wres3xocvs9tpkn4fu      (ybptxmszcng89e3sisfytlxnl_j),
  .akk0_n8kvb1w0wxrz            (ebpt710a8zup4xs8xzo        ),
  .cuxay1hemfm214cwu1513x         (1'b0        ),
  .s6in6vliinq9udhsofa         (1'b0        ),
  .ephp7dpea6ymyg0eucjv0        (mbghtxhocdjiarvwm96k8n5    ),
  .w42z5c2wv916u4df79p            (md5rsuwww5y3iwkgy03x6        ),
  .k_7iagb48feg9b3wj         (64'h0),
  .cnp1c4afdljmpemgot3sa     (1'b0),
  .wsh7h1p7b0zifvs0kwabih        (1'b0     ),
  .qhk0gez3kmex8twzly7mxn         (1'b0     ),
  .rafwujb8lw59lcbn9vsz8o        (64'b0),
  .dqpwtmmizdh6bvzsx6          (1'b0),          

  .plk8ixck4wj7c              (64'h0           ), 
  .e7nqb0p7cffw4lrkd            (w1et7pt4n96m3703shs          ), 
  .ej5tfrzf8ad7noezo8gdkb1xg4 (qwcb6hcmvfqmf032z        ), 
  .ekmvur7r4qz7ea7htd           (alu_cmt_wfi             ),
  .ndvqmbwgzq08mbdaxnn4        (j39tby_g7kqga33w_m           ),
  .dorqi70cvs05s           (gv5x7tbabwro1zc6cvwa        ),
  .pgfbjdj832ly_           (t2qvskf77dx_qfcl1        ),
  .z0yti764_a15nwanb           (j3iskguxr07s_auk4h        ),

  .k5yu5na0oo41y           (f136__ouz2d6kha2        ), 
  .n8g2a10i7cbowtvjhc           (ldzmdnb_744cs12l0t        ),
  .pzlsmt96uolwfb47           (so92sz9arx155dg58        ),
  .uzn8ik3rkkwib6p           (oxmshd1ilks70i3zxfapd       ),
  .kh00jq7wde_slaj           (qpscc8xem                ), 
  .rezwnhzl7vmkg           (u3wdadynlf                ), 
  .nq_d1dxi6n86s           (igvq6tvqkm                ), 

  .z8xxe17sssy8tr8q219         (otg3fn806ut                ),
  .rx4zxlit4v_5k4fclu      (zz7qeo73h2suy9k30jfzo    ),
  .vq3a19my9wldb5hug_nnbu0  (b9dlu6jwb4xgx25wfn5okd_7xyqlk),
  .mn8sk0gr9oh54zn_o       (q_wc5085zblpey              ),
  .oetzq1g528ymdza0maph       (srowfx3o2v3rl              ),
  .x11xtpe4e78unv1ahgzinz4n     (ofxcqyaipegys            ),
  .ialrcyi5grz5o0hc0jyjuwv     (jyp69_3c6ce00h7e            ),
  .bwsazwvhtn9in7lpyjssdk       (ipoo1harz8              ),
  .wfpum3du8gc8hr_xuerx     (e8fbphi7t5pf39a9p            ),
  .aly0oms0x8r1kmmdgyob      (od2labe2838d ),
  .vckb4tc8r10z7n621obxkju      (nb3g7kcdyt7bwtvq ),
  .f3lw5s13_0u5q6o4ep      (u4vwxxdwlql ),

  .u4k7uyzg9lp3zlf           (qh5uw_vgky8ctx9s             ),
  .rtjejhmafpq7db           (vfye1vj155_k              ),
  .vnc88f08k1s0obtnvb           (vujduks2o30              ),
  .u5pfnkzvz6fsvmgw4           (y4zqru1tedm              ),
  .zlk2yur1jgjwg           (q1coyps2cz7xe              ),
  .ow91ik9ily4bugcc43pp     (ch8qv98q9xu469etyz8oj        ),
  .bf8iyrsqp4a2s           (sibtd2rf5j              ),
  .pu764metopn524rq4hg2c24   (aiok9wht8yx8u6dz1e      ),
  .j7l4qmkctu4k_1q6c         (z8t7w6zr5woh649            ),
  .x6t2ufv1z2uufogo         (mg4yq4mui7ruja            ),
  .q5_q35rctah_              (g_o2wra9n9s                 ),                    
  .hm3iwty3s1d4si2p4           (oli3_udj80h6urj              ),                    
  .txcys7e9ezk6xikpy2hu987  (1'b0              ),                    
  .eph11j28sez0oftr7b         (g5usf8ixwjaxjs1m            ), 
  .lq6932o27hlk9v4f1m          (pxhhgm9746n             ), 
  .sll07sleuwo2fkitj       (fgm5kq4y725x6yylw          ), 
  .v2e4q5r07qxd6fxruqia3f       (awld9ngcypgfxa          ), 
  .e5nqx8gg2u3gxy0y4c       (v5m66onlnmxeejfhn          ), 
  .ajka24wmafrwpta96cf2        (kfz3mojvfh2fsfd           ), 
  .bod813pzaejozw9p1         (m05tjqf24b1fabuu0e        ),
  .z1et08p41uxcl76          (d40y0va2l7xzj  ),
  .jymdjzitd0hv0e9uhul        (hhj5975j18r0n),

  .juyjh9cdf4vvzhq         (zj0wqwminaxn            ),
  .pwppbjb8emt8vd9_w        (tkm5u9dl8zav4           ),
  .z69pfny03ofcxvjyygmo6      (eaxqugrf_ryu5rxxw41         ),
  .cvqaktep17ac            (vvsvl34lm1_1h              ),
  .h91pmjbyad1itr37            (r_p2yyjhd3              ),
  .mtsy6_whdwum2fu            (b6cv9yeaga7hf               ),
  .k_igx5_oeq1ag3m            (fpwql5ik7_sp0               ),
  .th3snuy_v19o06eanj        (dwci8hbxok739           ),
  .xxggjmznfu9b_             (nnng_p6632p                ),
  .imj0glh0tzynz           (ipht6ss_sh6h                ),
  .t9kvx890cyg              (t05leas4w4r                 ),
  .i984chc2gxtcivks          (bdhv0j4zhtx9nxmz             ),
  .cyudxl51e               (bwjyqadn                    ),
  .nv33gk9s6_               (k_pblo0),
  .w37tf6nz0oty_z89xv1          (qdh2itqlmn859kps6            ),
  .pfeci7n4c83yiwln58          (g2515ltnbxvz            ),
  .mzu7xfmjf4mwa0b           (u8cs2vcqau77o             ),
  .g3t8ql0mi58ddizau_8t3       (k0tpiu_dns7fesh         ),
  .gg468ty1pm6_zgec           (h9v5a720moqn805             ),
  .jtvucg9wp5nxn           (q3l2pm3uzu4             ),
  .ofe8xctslv6q5w48ky         (dsff_1r8ibc2u1kl52           ),
  .axbsuznhe7w6rrd            (fqizcmmfg               ),
  .j49by1lxo4ie9_ho            (tbuacpjktio               ),
  .tv7ak8mtfqswt            (ciftsjs2bvaxns               ),
  .vh0cb71_xnjsewqur3       (1'b0                    ),  
  .gbgabhg8e_ul0e24r6jq       (1'b0                    ),  

  .rgip60bn9st8htirgmhnohyj     (1'b0                    ),
  .duo6acmepph_0ahl_0ebyyjh   (1'b0                    ),
  .mylxtynzir7dvcouvb5thi  (ncr4iqrzig1xhs584u         ),
  .o5yttui8un64i2r3s3yxxxjc25iwv(g59aakolhtnl6vjex       ),

  .fxsynukaasxx8lt57bwdodyn3cem (1'b0                    ),
  .oel93f4rkl6esczbag9yld      (1'b0                    ),
  .vmp6zvyj46lrfmg3bl_kecu59   (1'b0                    ),
  .gj_lc7e2uh1cdx5b2bmynhvw  (1'b0                    ),
  .b7ker79ak62g5qei_oa7kxdm0  (1'b0                    ),
  .i3rcr_tmnynzs9lr254bac9x2b (64'h0      ),
  .ti5a3yv8_m3rzzigzeuzrt1 (1'b0      ),
  .cb86_62ddnv8i2whbc   (1'b0      ),

  .i_2lk2qupeba0sjgw6sdnbedc (1'b0                    ),
  .a46z1a4rlrucmwj5ju3o83orp8jx2e (1'b0                    ),
  .ti9h9knu4vrm6k3vqry9vfxbc4b (1'b0                    ),
  .p8zi9oi86dxmkaq4uqhu8j1hl0e (1'b0                    ),
  .plmzz80_s0_tb0kwjjgu5p7uktpi2 (1'b0                    ),
  .z_r1pp7wjooqw6n7rnoyv7nka81o (64'h0  ),

  .kr13pzf9ml9ic_vbl            (jw1vgacy_r0vr      ),
  .wkixlev_tj12x_lfp6p04t      (1'b0     ),
  .jzx45r8bb79aj5ddz7h_565f     (1'b0     ),



  .akdv8vv97zk549v            (gldc_bv5wpppiij9         ),   
  .k_wnu24cz94zwh8            (ljghmx9gec8jr0of         ),   
  .g65q46nnz7gip0zyo          (                        ),   
  .v8zi5h4rj36jt              (tyvyxz0mf               ),
  .livvja2ywo91o8v              (iaejzw1j2jb5i               ),
  .t5p9q190fm              (aucihtckush               ),

  .jdngc81st67hk8p            (qw6ymq0u4qknlwh             ),
  .u4t194j1c9najq            (td_th3xz1iyqn_w             ),
  .gkzjw6iff1idxo            (e25k01aox4_             ),
  .jcj76rmi3pqujm3v           (pdwodu8jbockhftk7       ),
  .ptu54kun7juh0           (o99cbvjf8lyjdj            ),
  .tsns5phts_z2fnf           (y6tqh4z7ck7gj            ),
  .rsdyvyptjiksvewu           (kzdc2z8f1n1qrac7            ),

  .fw_dplmj46w6              (                        ),
  .zf1w750jg2mtdij            (xyq4s_ubn1sx2s            ),   

  .dckyl_qt92wqvghtw3          (oajzut537ryb591kzk),
  .vyug4w9rb9kj6bmwwu          (qos_22gbinvor4),

  .h40f1u8xaz57o3c          (),
  .bv8rdomgcr9w6r2z          (),
  .ujgn98iv8k5xidjk          (),
  .pysgbgu5mzucuewf1           (yh8eetxf0xs392            ),   
  .pw6i533r0oou6ub            (bwd5a_yj_liikyo             ),   
  .getq71b86zu18ri7x        (piiqrjby8_d9dndhct         ),   
  .iouqv7uynzgvde_v             (b7fov0er1gnx              ),    

  .h_4gbwx46f8brur_wc      (ksgamvgvgr9n02_txmv       ),
  .nabilb10azux1hnithsys     (qrodgqtao6oexta13898      ),
  .pcmvrs0wuwr_x06ql         (s4ec4uwf6ke9r_tpu          ),
  .du9lzthd93rvmfcw7rz0wap    (o8s3z5xdvprqa0193p0),  
  .q2vmic6hc_08xqnvwhw          (kxcwjr8ri3x86f           ),
  .v175vi3kjhjhl37_p       (                      ),
  .vir1r5sxmryfghdpp_u82bq6   (                          ),
  .soumhrmo71_bkr9v6s5       (                        ),
  .fqx1jny69kgy_gimut      (crpiujipdzd_h3djv_bjup       ),
  .sd2su0k2v13e1jhtkwj          (sh7px5ghy0tmin8           ),
  .r26sxdceh7f2t6xroiyejiud7e  (lgs2ndps7oi98rleg8tshcz   ),
  .ruzuip2lmd_5bjdch       (),
  .t7xboey2yuqaq15sxya1b5      (),
  .v4icsnfwb3y76_4utq       (),
  .u4560ic2z4t9ft8jb0rvw      (),
  .de7s4aih29brxnb18p        (),  

  .hb36pq8e0n24raht15       (gjfmlxjpnnka6o8odi        ),  
  .xphk4z06widyipxfcjr       (mbwb4j_f4iygi4phniwt        ),  
  .j9fcegru44_r74xlm2sbp     (a6eyass0uv3sh81xwu      ),  
  .uw1jajj_fvu9278tlptmv_     (zhaca_k1wq3sy5wznci2pu      ),  
  .xcu8n5tos13pfc6jhw22       (t8qh_jt867ifbzdy0        ),  
  .tdwhghf609ku2jek72pn3     (l276zv1sj136kk9s9_unb3      ),  
  .lbx9pnfl2z4is68kam      (g_cuqgaizsk_nq6fwir1_  ),
  .hl9x8gmcd9k2ttm0hui2j      (rrubg3ioxxvdto3bjmpfsy  ),
  .ioka849821_gx48yl9gk      (if5n6cmdrvnn2c0vt09  ),


  .cc7_9__0hrnupts              (onacehe6tcgr               ),     
  .pba2_zyealgm_jf64t          (pv44129rj0uy831j6           ), 
  .zpdph1sve               (jwbql4ta0c                ),      
  .o9d_zhwhmsph               (kmfvezt2                ),      
  .dte0cay394mhjhkr         (omler2igyskatx              ),
  .cmbn4qx1zcverw            (zcl5hta0nld             ),
  .r9098zakm9jc            (rdce2xlm_syu             ),
  .ye_x11o9y0je9god            (y3lf5lq_1tfm1iea             ),
  .tp46wehs200pll2qi           (x882ucszl6qqk9m7            ),
  .vyis_kjmkr7org4mer          (yd1xmujxb33j01a4c           ),
  .n20czkexgpbptzj5w          (i6yx610m2nd7razu           ),
  .uvysjueb4qilrx7           (luf9wadz1xvpbt            ),
  .qd0yrkr028oru_36lsp9       (ohftngf40mc7275vq        ),
  .zkhg8302rekq3           (r8b6cghj00gkt7            ),
  .yjox8n6veh2dfp4           (hv3n9x664ena            ),
  .xa_tll8bjyk6hu8         (zlp9p2qtwrt0ra6c7          ),
  .fwpoqfymdxr45bq2         (vqp0990pwh3u9u4f          ),
  .rnub9co3myzraj2l           (k_u427htf3nny            ),
  .azbeqtr4zo_xorty8           (snxyhe6q4j0ik6is            ),
  .fv_51fuukywshp7hm           (di_rao90w5qbjlfn9            ),
  .w20nxrvpdf716_           (r43_rk2c1l4t            ),
  .x2ypwv3n6g8jsweuweebmhq     (h41082ijgnoh480fx5t      ),
  .dwvp6uc1acommla           (lvamcxldxlbi7k3r              ),
  .p8to9sivjjwpc0pn2bvf21se3   (c_vdpq9m03rq493zpv2165d3      ),
  .x9t5ge71i97il9r8         (ja6yz91tkse7r9tt            ),
  .n7fla3l_dqx9jnxul4         (rcp57t3vlm6czu6            ),
  .vg7c1san7ef_              (ho405be3bp1ma                 ),                    
  .umwzm3ilav51kmk7r           (t4zsjo_uj3n_m5              ),                    
  .c8l2f5n1fhxm76kt3vlu6jp  (                          ),                    
  .hibevegtudxlh_nk6e8e         (ytygj4ti9khaqpbhp            ), 
  .y6lolb8cmealsn6ev          (d9hqn06qm44jqmxo             ), 
  .x2bck2rbbpoyqbz62ld0tg       (hpf6iii62xdb170ho7ax          ), 
  .abkeecplc6ueo97vo24tg       (ckkfhtew3eup3984z          ), 
  .b_fk_j1filrux_uod       (dved_rrjqsz_ib5rx8          ), 
  .oaedrllyjbu5y92f        (p_gj56fnt4qky4n6sxai           ), 
  .plgwduxqtms73miw0         (pjz1nevm60h9ihnmunx4        ), 
  .mf_okovo5c__xpv1x          (),
  .i1_2srs1sequ9t          (),
  .a4aa8t_dofc7_82w          (),

  .q6sud8b_vapga5ru5c           (ob602_qjqak28zc1l            ),                    
  .latkf6ie2l8fv5dg98qec         (hu2q59l06nvqg7i7f          ), 
  .azmawprujj_u7q6ofj          (                         ),
  .wigxwsu_39gcyutr_re          (                         ),
  .l0_j3191k35720flisiv          (                         ),
  .cf059q4pm79who8jb          (                  ),

  .pket_pq2m99ayix3fk5yps       (),
  .ty49bqt9pydf4fr50f89       (),

  .itofghyluwwiwmqnj_4imeao     (),
  .j47kiegbvv22z361yv9n5   (),
  .r75dlj23fr96kve4fzd8xpw2zn  (s2mopc8npltdcmohj94          ),
  .mx7juirxj661i6i9lns4hnnyw0ep(ab20niin2uxlfv9w5s5n7y        ),


  .frehkmd0xqj4qeyqqodmp0onx7 (                        ),
  .ms95k2pmbvtrb33p5oa2q      (                        ),
  .r928tvy6d88uh6s9qun65udol2   (                        ),
  .jtgchf8072p4v1h9xclp0t  (                        ),
  .jekm9yqqqogc7_czwax0r6an_f  (                        ),
  .vs9f2qtmvyxt6ycc5e_z47fnjr (                        ),
  .wvywyxp28r9wdwncg13zbc_6    (                        ),
  .suaktr_howpmkqxx3p5j4      (                        ),

  .mnym6ha4fxtg2oqq9hlac5s1      (                    ),
  .p6wfurur4eut85r8tktdi03zxb   (                    ),
  .xxr9qx83ggzl9q98ig_ys5w60a  (                    ),
  .lozr9fiy6p7y8rinc582m2bt2ha_xmf  (                    ),
  .u78ade2idh660umk_1m66fdlksb9b  (                    ),
  .z3j5lbdgqwmp5zmv4g_zn29fgvintdc (                    ),

  .ussyj508sxu9v0           (y9bk3uc02upz      ),
  .pdns51exd9ffhf5pykv42sq     (),  
  .k09nslb_nkoy4r0t34xu6    (),
  .crr9jljkvi3gsixv1_v8       (),
  .sca7p0942a6kocjqqvat       (),
  .go_m73qp_w0p7abohs24       (),
  .jm4ru1fdiqtw706w8        (fq4r9kho3s5rkyx  ),
  .j021ufdslrlb4m5c5h2      (b1_o25pwqim0zl2p159psk),



  .p1kjflyurzeuxj (),
  .yvjlu1e9eng5_5tme (),
  .hh8nc68zrpki2m9r (),
  .v8wv99vga5gkl8xhk7x9in (),
  .ahfx5rs9jkdyw3b8ztscfx (),
  .ts3_k4ergzh8upz7 (),
  .ktqya1x1mfi5j3q7 (),
  .z6njhanl_m_hv48x5i9y (),
  .dvm_h24fnflt11prmyvme (),
  .uvyubcp0tbk9yirhz (),
  .ivoui15mvw3de5ds44 (),

  .gf33atgy          (gf33atgy),
  .ru_wi        (ru_wi)
  ); 









  wire                     p8fm019vnx8ax_2_  ;
  wire [5-1:0]    i_17_dtjvzuo  ;




  wire                     olti9ndjvk_sohpa  ;

  wire                     nvpglpdnii1iho_rjkw8 ;
  wire                     h7szh92q4s7x6vx_   ; 
  wire                     zf3zgw37xlcc2o5eprc5k ;
  wire                     gzyfsm1lj5vk008   ;

  wire                     pjcdn7d17lcskz8qw3fi;
  wire                     c3edim0hxqlxh7ubn4hn;
  wire                     seyk3b__57tr0b_kv__y;
  wire [64-1:0] bymbiaovszt6x5okz      ;
  wire                     qb0v08s4r8feqekkzsn  ;
  wire                     uyh4zz3rdydme0z8m4r  ;


  wire                     zhmxkmggxfi_lkbi     ;
  wire                     qaa88tv5k9oc8zha     ;
  wire                     v3qougfmuenqjx1x5jpd5na;
  wire                     khxw8wn6dnz9n8jiacgq3i  ;
  wire                     ochxbfnjjoa52cv6jxvg3k  ;
  wire [64-1:0] rrf9cbyl53_nsr_sro      ;
  wire                     usdwk0yslx167lf9z58wa3;


  wire b1nlh4cxd_uoj3g   ;
  wire s0pkezm5eltk6mmh   ;
  wire nc7x0kfw1l45cj_qx   ;
  wire y7rwp45w4w_msnfk   ;

  wire ko3lr4ef3iromewayub;



  m0m7t4t8fpmv   #(
    .hcl69mdlw0ykna4ue4_t1(1) 
  ) zci1nbrhuad663ie9oe0kze(
      .w2h8uh3l463qbgqmv(1'b0),
      .tywculgjyor8ndw    (tywculgjyor8ndw   ),


      .pw3qcykea5ib_ieka(1'b1),
      .g6xvfy8tj0zmajl  (1'b0),

      .rvr30vvllni (rvr30vvllni),
      .z1cj655u31 (z1cj655u31),
      .lhu2z948o3n (lhu2z948o3n),









    .r0s7d8cr68i2qs1z     (r0s7d8cr68i2qs1z),
    .kakelc68be0x7tdm9b9o    (kakelc68be0x7tdm9b9o),
    .j3j1czgoam48vhs8auo    (j3j1czgoam48vhs8auo),
    .gm1r5itc44uxw_y0_msk    (gm1r5itc44uxw_y0_msk),
    .af5qc04tmn51e4u2h1z    (af5qc04tmn51e4u2h1z),
    .qwcb6hcmvfqmf032z    (qwcb6hcmvfqmf032z),

    .jjzotrbn             (o8rffdg1904azl0q),
    .hw1_k1jmu             (f0ziihie9il3138m),
    .i7vhyhns            (jvi2i2xkdm88aoes), 
    .lu44s70ub62            (hnsixpix0gzu), 
    .qbpmsk2              (omler2igyskatx   ),

    .tc88s6cm5b               (oajzut537ryb591kzk    ),
    .c3sszdooylrw               (qos_22gbinvor4    ),
    .e19iv2rqeu5          (ja6yz91tkse7r9tt),
    .m4y6v4ncsg          (rcp57t3vlm6czu6),
    .le3dqob2            (lvamcxldxlbi7k3r),
    .cpt0qfwiz            (5'h0),
    .j_rvclhfbeig5cqeb3_   (1'b0),
    .qpyjufa5h7y               ({64{1'b0}}    ),
    .hvv94pmafz               ({64{1'b0}}    ),
    .sjunepbdn               (aucihtckush    ),
    .yocn4o2zav           (64'b0),

    .veibgbyke             (1'b0    ), 




    .zawjtr32pktig            (t4zsjo_uj3n_m5),
    .vc529nuu             (3'b0),
    .xh52jycxcjs         (1'b0),
    .aziir_r1p           (d9hqn06qm44jqmxo    ),        
    .rnx27onf2lbe          (1'b0), 
    .ya8t4ev_aidf0t0x4or    (),
    .scadliwzjp0l78srd9p  (1'b0              ),
    .l6s_gf8go82fwn           ({64{1'b0}}),
    .afifdv1w9           ({64{1'b0}}),
    .u2bhabgcppcy           ({64{1'b0}}),

    .cj2osby26qlape         (ob602_qjqak28zc1l),



    .ojbpo5z6urt             (xyq4s_ubn1sx2s),
    .fhhe7189lmum             (5'h0),



    .t9b41sw5vpr  (k_u427htf3nny),
    .bfo1il0du_  (snxyhe6q4j0ik6is),
    .gnb98c7tbqat  (di_rao90w5qbjlfn9),
    .w4kjodkdva03q  (r43_rk2c1l4t),


    .hy14_6z7grvldvw(vqp0990pwh3u9u4f),

    .nrebzehsuam    (b7fov0er1gnx   ),
    .bvzc7t76o17 (pv44129rj0uy831j6),

    .begxws3d6mwhnm        (64'h0 ),
    .z1nw2lilgog_        (64'h0 ),
    .x6ywulzbb7jp        (64'h0 ),
    .b9mfhl8am_whqquz         (fq4r9kho3s5rkyx  ),
    .bqen_oh1ujvq9lj4       (b1_o25pwqim0zl2p159psk),


    .bwjyqadn                (jwbql4ta0c    ),
    .ipht6ss_sh6h            (yh8eetxf0xs392),
    .k0xug5g             (kmfvezt2    ),
    .b_sdf8               (onacehe6tcgr   ),

    .n1rp2mggtiknd88         (32'b0),

    .b7ilo27jne5k           (yd1xmujxb33j01a4c     ),
    .piwiqvrjoq           (i6yx610m2nd7razu     ),
    .al4xeg8mukgfg            (luf9wadz1xvpbt      ),
    .ryc6z1c7rmzrnlno        (ohftngf40mc7275vq  ),
    .rhufxsnopy0n            (r8b6cghj00gkt7      ),
    .wbhvg_1r9435            (hv3n9x664ena      ),
    .s1woka0byzgo          (zlp9p2qtwrt0ra6c7    ),
    .q8977k41y4             (bwd5a_yj_liikyo       ),
    .ciiwo7qhifea         (piiqrjby8_d9dndhct   ),

    .binjv97px9r7dt04h0       (ksgamvgvgr9n02_txmv     ),
    .ajl4tppx98ihuirj_mxih   (lgs2ndps7oi98rleg8tshcz ),
    .o_d157fc5_l           (kxcwjr8ri3x86f         ),

    .u2k4dyp52s_m             (rdce2xlm_syu  ),
    .djvj1e_             (y3lf5lq_1tfm1iea  ),
    .bktu0z1mk56             (zcl5hta0nld  ),
    .l6z1pzhjg5az            (x882ucszl6qqk9m7 ),
    .phofig8d5zd_8v9g8       (phofig8d5zd_8v9g8),
    .js0ml55dtie8qenb4eoj2 (js0ml55dtie8qenb4eoj2),
    .p343qo1j             (ticm3jrqt6tjtf6),
    .h8m3g7a             (hpaul9bznamp4qkl),
    .r9ix0zzks6zej       (vq7jwn83uus_ac4s4ghf),
    .l8xeqkc               (gzh3us4_ux10aey),


    .v35y3qnk7mx3l1695     (v35y3qnk7mx3l1695    ),

    .gqe6zqljzhgt5wz98      (qfspmfi47b5jx99i0     ),
    .tisftwun8guh8lnibary2gz (pjcdn7d17lcskz8qw3fi),
    .wdgj6jexv3_u8sb4gnsv5 (c3edim0hxqlxh7ubn4hn),
    .c_qlgbc7oqwu9as946yqls (seyk3b__57tr0b_kv__y),
    .nc5hf3a4mwl257q       (bymbiaovszt6x5okz      ),
    .cqq719hbl6kax00mwmrhj   (qb0v08s4r8feqekkzsn  ),
    .a_x852mvzp7z5occs1   (uyh4zz3rdydme0z8m4r  ),

    .v3e6l1k7eo9k3        (khxw8wn6dnz9n8jiacgq3i ),
    .hxrmt706n071lic0f7       (ochxbfnjjoa52cv6jxvg3k),

    .lrhkvgg4x13sq245     (                   ),
    .y45254ns5fjfjnwjiwr1_quk(rrf9cbyl53_nsr_sro                   ),
    .sshjsyphxbyaqk3kr    (                   ),
    .zu8yygom_ioh         (                   ),
    .od8eje0yjk8         (1'b1                   ),
    .l_km9bow2ubqs5dtd        (                   ),
    .cv8rkirz            (                   ),
    .mbnh9clp6pd3t         (                   ),
    .z091v3i7q4_rty4       (                   ),
    .tsml_wqqwnty         (                   ),
    .pdz01l48nt          (                   ),
    .l5zrepfg8it           (                   ),
    .aq4b6s94dp0f          (                   ),
    .dmg1a5xdc9           (                   ),
    .v1j50zesdgxioc           (                   ),
    .tkhm63y407b          (                   ),
    .qhkm8drwygkskh_          (                   ),
    .nh1gz4628x89          (                   ),
    .l4anyablbw3gt          (                   ),
    .vn5b662w76_a3npe         (                   ),
    .wigtf10_bybfdpp_x        (                   ),
    .w2gbqib7zable3o        (                   ),
    .zp24wdce6ufxkpbs        (                   ),
    .xxee65tc1tureck      (                   ),
    .wr1tfb0_sg9           (                   ),
    .enhpakthwj3e65vldt   (                   ),
    .mz47ksy6nekv1cbaq75    (                   ),
    .egplp36i1ttcggdv2b0xo2e(                   ),
    .rbsutocgtudusq3v    (                   ),
    .sgy1x259o9ltvsfe    (                   ),
    .tr2dgjt2yqfzjaos9o  (                   ),
    .o8m475rdcb4y71zte3fbd30(                  ),
    .nzm80hh72kwblbx4fcg   (                ),
    .l9wonwtwviy4i8w6s     (zhmxkmggxfi_lkbi), 
    .wuw4k4dyuslqkjap     (qaa88tv5k9oc8zha    ), 
    .s4o6xx8w0dylrebxlqmia79t5 (v3qougfmuenqjx1x5jpd5na), 
    .isvwkofue95j9ud7p3nrgntc(q97rqfy8n7ixfm2a5wev4nd5sylpcq3j),
    .mf10lk374lxu341vp3kpfl6(lln3b7iev7jpvogh964ro_9bc_3y),
    .nkemiexuw_o6b34go    (hujgg6hjnhtbspbkekuz5_u ),
    .bnnsit7f_1yqs20xcxk3l     (v3pnt81kfrgbaanm1mhh51w  ),
    .c2vqeph9snojapvdushbj    (i08eq60d_snxeq8si_ezod ),
    .w8wwz5822d7298zis7      (usdwk0yslx167lf9z58wa3   ),
    .br6lhce3u3l01blvxzrqphj5svlum(              ),
    .zq261z2pygzc0_h44fo     (                   ),
    .g_w5s5kg5qk2w1gyo7odo2nubrxo0(               ),
    .b1iduhkyfb7xynn3btxh6lhgev7_(               ),
    .ndtc71v47ribx6u_eqsx8tdk0  (               ),
    .efp001u9ffq4ypu8uk4l8tbblt8  (               ),
    .fce921hmrlbrv4qdu4cb0pee  (               ),
    .twjiv2hewisn6o      (                   ),
    .l4i6kd5vs494chi      (                   ),

    .d7kpxfpyhil_2nt     (                 ),



    .jugi02ecegnos3        (r9hdxtws4mibgldl     ), 
    .rxjuugktc38un        (olti9ndjvk_sohpa     ),
    .h8wu7unf_ixmxfeh         (rwtwoy92pmk4i       ),
    .b84l246u4jmnu        (i_17_dtjvzuo     ),
    .kdpgigzs75vcc1d         (nlbav8h239dt2a      ),
    .uh251o1pav          (p8fm019vnx8ax_2_     ), 


    .suxmggt9hea4ao3r        (b1nlh4cxd_uoj3g   ),
    .kwn45x5pjj_5mi        (s0pkezm5eltk6mmh   ),
    .lp9c9xlhbpjow4k        (nc7x0kfw1l45cj_qx   ),
    .ts1jnweqrdhomp        (y7rwp45w4w_msnfk   ),
    .ze26d9sog9r3thx     (ko3lr4ef3iromewayub),

   .vjkz8n6i44pc7o        (),     
   .cwmxezrc3jv6hzxcfc (),
   .uig3ujuyq0_61kqb (1'b0),
   .xc2becmsn4fcniw6ks (),
   .nb3w1rq_ny95rvrt (),
   .p_yx415so7q1vohijb (),


    .rb050tnl             (       ),
    .e1go3iu             (       ),
    .el7_p8jit09           (         ),
    .a94vd35etec4           (    ),
    .l9erxxpnphqd26vg9        (64'h0),
    .guuvp01vkcryglsu1p3   (                 ),
    .hig2gwwbeuhnt65xrp       (64'h0),
    .vf5xcr67bqhzlo43_        (            ),
    .bj7h5jqg66r51jxki6emra   (                 ),
    .zmfo8cca_77pc       (64'h0),

    .vmx1fh4kmh4c             (       ),

    .v657dksgaz1cki9         (),
    .qzz1jhwf_vd0r8g       (),
    .dwn42a1uvd9x3myec       (1'b0),
    .uiojikf9vcnz        (),
    .x1_k6oouttg7m3f         (),
    .fcvvhg9v3mx         (),
    .l_v5xmhbzqc         (),
    .i7iq7ecm_d9pi6uw6       (),
    .p5fn_ooo9rctbxkgm_jui    (1'b0),
    .a5z_23_ryr_m29hhia_p (1'b0),




    .isz7jw04u7k3s7b398   (                ), 
    .q4_7fnx90rztwn6_8dybi   ( 1'b1           ),
    .zq2e9j_emlri_qjtg    (                ),
    .gw6s_h2ymbn1ds50q8    (                ),
    .qv749hsiom75nyn49v     (                ), 
    .vo_fj58ip6ok0srq7t5   (                ), 
    .qq819v1yyh8derngk15k1   (1'b1            ),
    .o_q0qt9vjpibgshm714a    (                ),
    .iqx3cqyh7_mpvu_9om    (                ),
    .melkey3fxhhc3e649p     (                ), 

    .gf33atgy                 (gf33atgy          ),
    .ru_wi               (ru_wi        ) 
  );


  assign n3zlo14nquu5l7zf3 = ngy4ipxc1vxym69lu; 

















  wire [64-1:0]          fyeewgjh0ejxrrn        ;
  wire [64-1:0]          zpg071p8a094ze4        ;
  wire [64-1:0]          odgaqp3aclcfht_i7t        ;

  wire                           pjybabc2ndhp9w15      ;
  wire                           r8n4jj_yqo_psdycdpf      ;
  wire                           rc1qjhv_cq1wdp4lltk8      ;
  wire                           nw1d2c3l16ufwicfgjc     ;
  wire                           gtuyw8lwe5vig3whpwia     ;
  wire                           bepi9gxgibkbsjimgygx     ;

  wire                           mgtrw760fgm5m362j      ;
  wire                           id6e2963yn91s9_9_5on      ;
  wire                           kmw5zvgvlfxa11v33    ;
  wire                           sb8c9xuda2cis65y1ho    ;
  wire                           llejtcklcswz9nau7td0r     ;
  wire                           og_162hdl7wzfuaufz03z ;
  wire                           oy6he9jrp6z3la4aonl     ;
  wire                           w6j6nqqawzzgqlkzfpnm3     ;
  wire                           e8ek1pn7po43ud9g42t   ;
  wire                           o60e9qmmyfyb4lr      ;
  wire                           ymf9djwm1ss4fvtr68bfi  ;
  wire                           cgok74_0s8wxk7wiu3hnx3w9l  ;
  wire                           vqixsqz3vz_o2ze5ovcwp577;
  wire                           erx90sfzu891aujxq      ;
  wire [64-1:0]          qtfwu64s5lqiyyqles        ;
  wire [64-1:0]          y4so7d4uu1lfqzpbgq    ;
  wire [48-1:0] gyxiq3yqdnanuqt16bh7r0h   ;
  wire                           ie4dehipkb3b8__y5dt     ;
  wire                           zv7y8twrabykb59a8a4629;
  wire                           p1xbmu6wvqhuu3rp2xt     ;
  wire                           aq9__1ut60olwyc0dv_x     ;
  wire                           vynn8pxcf1uhro7e;
  wire                           p6pm4fdt9wqk___preo3g4ppz;
  wire [50-1:0] gc_pvwtyrxrfkd4sh3xn;
  wire [105-1:0] ynb8hbtopto1okekngx8;
  wire sfrkf5j74_e8qi;
  wire qryqhxq_uj5viaeq_tql;
  
  wire j09fc8frtaff7iig7zoft;
  wire [48-1:0] iecuqnis03sogixkg5at529;  
  wire [64-1:0] w9gp9paa_nei_cgq5;
  wire vtx1v5trwp6v5uo05kirprri;
  wire nvvhnw32pu5ftxhzv6ycffp;
  wire kfooiskivym4ubj3utuxjy451;
  wire ihlsip_az_gbdtb7cn43tr8wy;

  wire                                   pt8li1mpvd04qujh4o;
  wire [48-1:0]  kgd8co1m3ta9_sciodf;
  wire                           l_h0z16ew816k0kc59fz  ;
  wire [19-1:0] v1_i1c87etnhn8gl6t64rr;
  wire                           x967n2unm25k5336wf2 ;
  wire                           x2uw3xkpg8k47k8i ;
  wire                           po0i9bzsw2yj9tv ;
  wire                           ucybeaa15_qx208e ;
  wire                           pl1e1zu0kmorvnh8dd1yd_7mi  ;
  wire                           uh0wfy2udciats10exk7gx  ;
  wire                           da476r5mk9l38ofvakaxk118t7 ;
  wire                           n1vkvib_j_0t8v7t7pjy3uio26 ;
  wire                           r01knk1me0t4m3ue2ok4t6m ;
  wire [4-1:0]       q3ob282pxl36b1j5u1cpl5ets3r;
  wire [4-1:0]       yrg9fg2dzj0h1004qftims1;
  wire                           imk1vol1t7hn6gevzps7ze  ;
  wire [4-1:0]       voug2bdbrmjvpkny8ect9r;


  wire [64-1:0]       cvvsn7xc8qg5uk;
  wire [32-1:0]    xnf360j941m2n;
  wire [64-1:0]       phiz5ah_lfipt6fb6lfzws    ;
  wire                           eih6zsu_r0tzn0s9udfs5ie1mxg;

  wire                           jpplkccgktsmzedro78tuuvm8    ; 
  wire                           hnq2agjqmp3jnfvc02q9vn   ;
  wire                           b04f0gnze13bj90dolndjwsij1e  ;
  wire                           ga193bfpsqosp5on_bftetcu19  ;
  wire [64-1:0]       kzmdmorjvnpxc87jh5yawhk    ;
  wire                           dibc8pgq7tvu40lvceswojwq;
  wire                           rqprsakhpq9fka9os5knx7kiw;
  wire [64-1:0]       vmspdud3fb2xydastwgm95;
  wire                           bzjveslpnkrl4_vnqp01r2;

b0gv4gv3sqckul0vbemwxr#(
  .gdctpuyrfi_b (0),
  .l_7qc0w_2x6i(0),
  .t5462hhws9i6ynbxi(1)
  ) shxbj388mfwfn7(
  .cu1owrury8wsed               ({4{1'b0}}   ),
  .mt1z8r_sz               (pc67uztpd_zg6bsal       ),
  .uc9k3lw_iehx               (fs6jojwsl0l32t7brm38vh   ),
  .radwr7skyhm3jqso5         (ydtm1yuxqj7fmxvqc    ),
  .zdid44qi3bv7q4phl         ({4{1'b0}}  ),
  .x4owqbu74zh_xxr         (eo5skx1ygvzuasbjgnyl    ),

  .b43m7n67rav8he           (1'b0      ),
  .qcutfgh43gov5u4urt           (jf9ko0etxomcrj25  ),
  .s73raoa0ilom1wyi           (qd5sbh8mupp_n4y95vo  ),
  .dnwb40nhmse7rcj0epzjo     (vz63qkw5s3m8urb9       ),
  .omeribg0gbgvpn78urilv_a     (1'b0),
  .jxogr1vy8jotyh8ivd2u     (p1jdw9loxkz60taq_vkp_3       ),

  .kl8zh4diafqs                ({64{1'b0}}    ), 
  .jiartjoiycj2                (mne0dg23_1aal06pio        ), 
  .dtypmpwq1q2j                (s7vgjm2azmcc3uzzdc_7   ), 
  .uwl7jm0d1lv0xpo            (1'b0 ), 
  .u2l80pdclhyu1bl            (1'b0 ), 
  .uamf3ccv7ouhi18            (1'b1        ), 

  .pkw60eo867gghh          (iojqlhtwx45_siz         ), 
  .strg8286lgex8p4_0m          ( {64{1'b0}}), 
  .avpvrch0prpui67          (jwwku_el5h5h2lx6e0kyi ), 

  .e7nqb0p7cffw4lrkd      (d9_s5e6qdqa7haet4s),
  .dorqi70cvs05s     (o99cbvjf8lyjdj),
  .pgfbjdj832ly_     (y6tqh4z7ck7gj),
  .z0yti764_a15nwanb     (kzdc2z8f1n1qrac7),
  .k5yu5na0oo41y     (qw6ymq0u4qknlwh),
  .n8g2a10i7cbowtvjhc     (td_th3xz1iyqn_w),
  .pzlsmt96uolwfb47           (e25k01aox4_               ),
  .uzn8ik3rkkwib6p           ({5{1'b0}}       ),
  .kh00jq7wde_slaj     (tyvyxz0mf), 
  .rezwnhzl7vmkg     (iaejzw1j2jb5i), 
  .nq_d1dxi6n86s      (aucihtckush), 
  .z8xxe17sssy8tr8q219   (omler2igyskatx),
  .mn8sk0gr9oh54zn_o   (gjfmlxjpnnka6o8odi  ),
  .oetzq1g528ymdza0maph   (mbwb4j_f4iygi4phniwt  ),
  .x11xtpe4e78unv1ahgzinz4n (a6eyass0uv3sh81xwu),
  .ialrcyi5grz5o0hc0jyjuwv (zhaca_k1wq3sy5wznci2pu),
  .bwsazwvhtn9in7lpyjssdk    (t8qh_jt867ifbzdy0  ),
  .wfpum3du8gc8hr_xuerx  (l276zv1sj136kk9s9_unb3),
  .aly0oms0x8r1kmmdgyob   (g_cuqgaizsk_nq6fwir1_  ),
  .vckb4tc8r10z7n621obxkju   (rrubg3ioxxvdto3bjmpfsy  ),
  .f3lw5s13_0u5q6o4ep   (if5n6cmdrvnn2c0vt09  ),
  .u4k7uyzg9lp3zlf       (x882ucszl6qqk9m7  ),

  .cvqaktep17ac      (r9hdxtws4mibgldl),
  .h91pmjbyad1itr37      (olti9ndjvk_sohpa),
  .plk8ixck4wj7c        (rwtwoy92pmk4i),

  .mtsy6_whdwum2fu      (xyq4s_ubn1sx2s), 
  .k_igx5_oeq1ag3m      (bwd5a_yj_liikyo     ),
  .th3snuy_v19o06eanj  (piiqrjby8_d9dndhct ),
  .xxggjmznfu9b_       (b7fov0er1gnx   ),
  .t9kvx890cyg        (onacehe6tcgr     ),
  .i984chc2gxtcivks    (pv44129rj0uy831j6 ),
  .cyudxl51e         (jwbql4ta0c),
  .nv33gk9s6_         (kmfvezt2),
  .rtjejhmafpq7db     (b1nlh4cxd_uoj3g),   
  .vnc88f08k1s0obtnvb     (s0pkezm5eltk6mmh),   
  .u5pfnkzvz6fsvmgw4     (nc7x0kfw1l45cj_qx),   
  .zlk2yur1jgjwg     (y7rwp45w4w_msnfk),   
  .ow91ik9ily4bugcc43pp(h41082ijgnoh480fx5t),   
  .bf8iyrsqp4a2s         (lvamcxldxlbi7k3r              ),
  .pu764metopn524rq4hg2c24 (c_vdpq9m03rq493zpv2165d3      ),
  .j7l4qmkctu4k_1q6c       (ja6yz91tkse7r9tt            ),
  .x6t2ufv1z2uufogo       (rcp57t3vlm6czu6            ),
  .q5_q35rctah_              (ho405be3bp1ma                 ),                    
  .hm3iwty3s1d4si2p4           (t4zsjo_uj3n_m5              ),                    
  .txcys7e9ezk6xikpy2hu987  (1'b0              ),                    
  .eph11j28sez0oftr7b         (ytygj4ti9khaqpbhp            ), 
  .lq6932o27hlk9v4f1m          (d9hqn06qm44jqmxo             ), 
  .sll07sleuwo2fkitj       (hpf6iii62xdb170ho7ax          ), 
  .v2e4q5r07qxd6fxruqia3f       (ckkfhtew3eup3984z          ), 
  .e5nqx8gg2u3gxy0y4c       (dved_rrjqsz_ib5rx8          ), 
  .ajka24wmafrwpta96cf2        (p_gj56fnt4qky4n6sxai           ), 
  .bod813pzaejozw9p1         (pjz1nevm60h9ihnmunx4 ),
  .z1et08p41uxcl76          (ob602_qjqak28zc1l  ),
  .jymdjzitd0hv0e9uhul        (hu2q59l06nvqg7i7f),
  .juyjh9cdf4vvzhq   (vqp0990pwh3u9u4f),
  .w37tf6nz0oty_z89xv1    (yd1xmujxb33j01a4c),
  .pfeci7n4c83yiwln58    (i6yx610m2nd7razu),
  .mzu7xfmjf4mwa0b     (luf9wadz1xvpbt ),
  .g3t8ql0mi58ddizau_8t3 (ohftngf40mc7275vq),
  .gg468ty1pm6_zgec     (r8b6cghj00gkt7 ),
  .jtvucg9wp5nxn     (hv3n9x664ena ),
  .ofe8xctslv6q5w48ky   (zlp9p2qtwrt0ra6c7),
  .tv7ak8mtfqswt      (zcl5hta0nld),
  .axbsuznhe7w6rrd      (rdce2xlm_syu),
  .j49by1lxo4ie9_ho      (y3lf5lq_1tfm1iea),
  .vh0cb71_xnjsewqur3 (gkfhdl1lvs93nq2q),
  .gbgabhg8e_ul0e24r6jq (a6qybr3pioqo0),
  .pwppbjb8emt8vd9_w        (ko3lr4ef3iromewayub),
  .z69pfny03ofcxvjyygmo6      (b1_o25pwqim0zl2p159psk),

  .rgip60bn9st8htirgmhnohyj     (1'b0    ),
  .duo6acmepph_0ahl_0ebyyjh   (1'b0    ),
  .mylxtynzir7dvcouvb5thi  (s2mopc8npltdcmohj94  )  ,
  .o5yttui8un64i2r3s3yxxxjc25iwv(ab20niin2uxlfv9w5s5n7y)  ,

  .fxsynukaasxx8lt57bwdodyn3cem (1'b0                    ),
  .oel93f4rkl6esczbag9yld      (1'b0                    ),
  .vmp6zvyj46lrfmg3bl_kecu59   (1'b0                    ),
  .gj_lc7e2uh1cdx5b2bmynhvw  (1'b0                    ),
  .b7ker79ak62g5qei_oa7kxdm0  (1'b0                    ),
  .i3rcr_tmnynzs9lr254bac9x2b (64'h0      ),
  .ti5a3yv8_m3rzzigzeuzrt1 (1'b0      ),
  .cb86_62ddnv8i2whbc   (1'b0      ),

  .i_2lk2qupeba0sjgw6sdnbedc (1'b0                    ),
  .a46z1a4rlrucmwj5ju3o83orp8jx2e (1'b0                    ),
  .ti9h9knu4vrm6k3vqry9vfxbc4b (1'b0                    ),
  .p8zi9oi86dxmkaq4uqhu8j1hl0e (1'b0                    ),
  .plmzz80_s0_tb0kwjjgu5p7uktpi2 (1'b0                    ),
  .z_r1pp7wjooqw6n7rnoyv7nka81o (64'h0  ),

  .kr13pzf9ml9ic_vbl            (1'b0      ),
  .wkixlev_tj12x_lfp6p04t      (khxw8wn6dnz9n8jiacgq3i      ),
  .jzx45r8bb79aj5ddz7h_565f     (ochxbfnjjoa52cv6jxvg3k     ),

  .lot9xvzuqrd5jm0scdx5t       (qrodgqtao6oexta13898),
  .mn3tic51ckga0gc           (s4ec4uwf6ke9r_tpu    ),
  .k0be3wres3xocvs9tpkn4fu      (o8s3z5xdvprqa0193p0),  
  .akk0_n8kvb1w0wxrz            (kxcwjr8ri3x86f     ),
  .s6in6vliinq9udhsofa         (qaa88tv5k9oc8zha        ),
  .cuxay1hemfm214cwu1513x         (zhmxkmggxfi_lkbi        ),
  .ephp7dpea6ymyg0eucjv0        (crpiujipdzd_h3djv_bjup ),
  .w42z5c2wv916u4df79p            (sh7px5ghy0tmin8 ),
  .ej5tfrzf8ad7noezo8gdkb1xg4   (qwcb6hcmvfqmf032z        ), 
  .ekmvur7r4qz7ea7htd             (alu_cmt_wfi             ),
  .ndvqmbwgzq08mbdaxnn4          (j39tby_g7kqga33w_m           ),
  .rx4zxlit4v_5k4fclu        (ksgamvgvgr9n02_txmv     ),
  .vq3a19my9wldb5hug_nnbu0    (lgs2ndps7oi98rleg8tshcz ),
  .imj0glh0tzynz             (yh8eetxf0xs392          ),
  .k_7iagb48feg9b3wj         (rrf9cbyl53_nsr_sro),
  .cnp1c4afdljmpemgot3sa     (v3qougfmuenqjx1x5jpd5na),
  .wsh7h1p7b0zifvs0kwabih        (hujgg6hjnhtbspbkekuz5_u),
  .qhk0gez3kmex8twzly7mxn         (v3pnt81kfrgbaanm1mhh51w),
  .rafwujb8lw59lcbn9vsz8o        (i08eq60d_snxeq8si_ezod),
  .dqpwtmmizdh6bvzsx6          (usdwk0yslx167lf9z58wa3),

  .pysgbgu5mzucuewf1             (tb198r6lzk1sr77g4         ),
  .r26sxdceh7f2t6xroiyejiud7e    (eih6zsu_r0tzn0s9udfs5ie1mxg),
  .h_4gbwx46f8brur_wc        (phiz5ah_lfipt6fb6lfzws    ),
  .nabilb10azux1hnithsys       (q7iyngsmbckvi2tht2wb5nh),
  .pcmvrs0wuwr_x06ql           (mq09q0m1l74z182ajkt2udd    ),
  .du9lzthd93rvmfcw7rz0wap      (xsziw9gaor0xrlm1hvlpjr),
  .q2vmic6hc_08xqnvwhw            (reu5ooijp0czeggc974     ),
  .v175vi3kjhjhl37_p         (b6p6azv95fkv2o7od5rkww9t  ),
  .vir1r5sxmryfghdpp_u82bq6     (ga193bfpsqosp5on_bftetcu19  ),
  .soumhrmo71_bkr9v6s5         (b81kg80kxviv6w2l2dt8qq     ),
  .fqx1jny69kgy_gimut        (m5mjr032v1z_erq3mxi07t3v ),
  .sd2su0k2v13e1jhtkwj            (kccav9va65o92d7d9d),
  .ruzuip2lmd_5bjdch         (kzmdmorjvnpxc87jh5yawhk),
  .t7xboey2yuqaq15sxya1b5        (dibc8pgq7tvu40lvceswojwq),
  .v4icsnfwb3y76_4utq         (rqprsakhpq9fka9os5knx7kiw),
  .u4560ic2z4t9ft8jb0rvw        (vmspdud3fb2xydastwgm95),
  .de7s4aih29brxnb18p          (bzjveslpnkrl4_vnqp01r2),

  .dckyl_qt92wqvghtw3            (                         ),
  .vyug4w9rb9kj6bmwwu            (                         ),

  .v8zi5h4rj36jt             (fyeewgjh0ejxrrn        ),
  .livvja2ywo91o8v             (zpg071p8a094ze4        ),
  .t5p9q190fm              (odgaqp3aclcfht_i7t), 
  .jdngc81st67hk8p           (pjybabc2ndhp9w15      ),
  .u4t194j1c9najq           (r8n4jj_yqo_psdycdpf      ),
  .gkzjw6iff1idxo            (rc1qjhv_cq1wdp4lltk8      ),
  .jcj76rmi3pqujm3v           (                    ),
  .ptu54kun7juh0          (nw1d2c3l16ufwicfgjc     ), 
  .tsns5phts_z2fnf          (gtuyw8lwe5vig3whpwia     ),
  .rsdyvyptjiksvewu          (bepi9gxgibkbsjimgygx    ),
  .fw_dplmj46w6             (mne0dg23_1aal06pio        ),
  .g65q46nnz7gip0zyo         (                        ),   
  .akdv8vv97zk549v           (jf9ko0etxomcrj25      ),   
  .k_wnu24cz94zwh8           (mgtrw760fgm5m362j      ),   
  .zf1w750jg2mtdij           (id6e2963yn91s9_9_5on      ),   
  .pw6i533r0oou6ub           (o60e9qmmyfyb4lr      ),   
  .getq71b86zu18ri7x       (ymf9djwm1ss4fvtr68bfi  ),   
  .iouqv7uynzgvde_v            (erx90sfzu891aujxq             ),    
  .hb36pq8e0n24raht15      (pl1e1zu0kmorvnh8dd1yd_7mi       ),  
  .xphk4z06widyipxfcjr      (uh0wfy2udciats10exk7gx       ),  
  .j9fcegru44_r74xlm2sbp    (q3ob282pxl36b1j5u1cpl5ets3r     ),  
  .uw1jajj_fvu9278tlptmv_    (yrg9fg2dzj0h1004qftims1     ),   
  .xcu8n5tos13pfc6jhw22      (imk1vol1t7hn6gevzps7ze       ),  
  .tdwhghf609ku2jek72pn3    (voug2bdbrmjvpkny8ect9r     ),   
  .lbx9pnfl2z4is68kam     ( da476r5mk9l38ofvakaxk118t7 ),
  .hl9x8gmcd9k2ttm0hui2j     ( n1vkvib_j_0t8v7t7pjy3uio26 ),
  .ioka849821_gx48yl9gk     ( r01knk1me0t4m3ue2ok4t6m ),
  .cc7_9__0hrnupts        (qtfwu64s5lqiyyqles        ),     
  .pba2_zyealgm_jf64t    (y4so7d4uu1lfqzpbgq    ), 
  .zpdph1sve         (cvvsn7xc8qg5uk         ),      
  .o9d_zhwhmsph         (xnf360j941m2n         ),      
  .dte0cay394mhjhkr   (pc67uztpd_zg6bsal       ),
  .vyis_kjmkr7org4mer    (kmw5zvgvlfxa11v33    ),
  .n20czkexgpbptzj5w    (sb8c9xuda2cis65y1ho    ),
  .uvysjueb4qilrx7     (llejtcklcswz9nau7td0r     ),
  .qd0yrkr028oru_36lsp9 (og_162hdl7wzfuaufz03z ),
  .zkhg8302rekq3     (oy6he9jrp6z3la4aonl     ),
  .yjox8n6veh2dfp4     (w6j6nqqawzzgqlkzfpnm3     ),
  .xa_tll8bjyk6hu8   (e8ek1pn7po43ud9g42t   ),
  .cmbn4qx1zcverw      (x967n2unm25k5336wf2      ),
  .r9098zakm9jc      (x2uw3xkpg8k47k8i      ),
  .ye_x11o9y0je9god      (po0i9bzsw2yj9tv      ),
  .tp46wehs200pll2qi     (ucybeaa15_qx208e),
  .fwpoqfymdxr45bq2   (gyxiq3yqdnanuqt16bh7r0h   ),
  .rnub9co3myzraj2l     (icczfaorqi6bmvsm5c4h     ),
  .azbeqtr4zo_xorty8     (ie4dehipkb3b8__y5dt     ),
  .fv_51fuukywshp7hm     (p1xbmu6wvqhuu3rp2xt     ),
  .w20nxrvpdf716_     (aq9__1ut60olwyc0dv_x     ),
  .x2ypwv3n6g8jsweuweebmhq(e0xd37xbhk4bxmxa9_93qr    ),
  .dwvp6uc1acommla           (vynn8pxcf1uhro7e              ),
  .p8to9sivjjwpc0pn2bvf21se3   (p6pm4fdt9wqk___preo3g4ppz      ),
  .x9t5ge71i97il9r8         (ynb8hbtopto1okekngx8            ),
  .n7fla3l_dqx9jnxul4         (gc_pvwtyrxrfkd4sh3xn            ),
  .h40f1u8xaz57o3c          (),
  .bv8rdomgcr9w6r2z          (),
  .ujgn98iv8k5xidjk          (),
  .vg7c1san7ef_              (sfrkf5j74_e8qi                 ),                    
  .umwzm3ilav51kmk7r           (qryqhxq_uj5viaeq_tql              ),                    
  .c8l2f5n1fhxm76kt3vlu6jp  (                               ),                    
  .hibevegtudxlh_nk6e8e         (iecuqnis03sogixkg5at529            ), 
  .y6lolb8cmealsn6ev          (w9gp9paa_nei_cgq5             ), 
  .x2bck2rbbpoyqbz62ld0tg       (vtx1v5trwp6v5uo05kirprri          ), 
  .abkeecplc6ueo97vo24tg       (nvvhnw32pu5ftxhzv6ycffp          ), 
  .b_fk_j1filrux_uod       (kfooiskivym4ubj3utuxjy451          ), 
  .oaedrllyjbu5y92f        (j09fc8frtaff7iig7zoft           ), 
  .plgwduxqtms73miw0         (ihlsip_az_gbdtb7cn43tr8wy     ),
  .mf_okovo5c__xpv1x          (),
  .i1_2srs1sequ9t          (),
  .a4aa8t_dofc7_82w          (),

  .q6sud8b_vapga5ru5c           (pt8li1mpvd04qujh4o              ),                    
  .latkf6ie2l8fv5dg98qec         (kgd8co1m3ta9_sciodf            ), 
  .azmawprujj_u7q6ofj          (                  ),
  .wigxwsu_39gcyutr_re          (                  ),
  .l0_j3191k35720flisiv          (                  ),
  .cf059q4pm79who8jb          (                  ),
  .pket_pq2m99ayix3fk5yps (w0p_8cae4cqs_1hdeoydtp ),
  .ty49bqt9pydf4fr50f89 (hncm6yp50zjrhz9dcp1t1q ),

  .itofghyluwwiwmqnj_4imeao     (                        ),
  .j47kiegbvv22z361yv9n5   (                        ),
  .r75dlj23fr96kve4fzd8xpw2zn  (cgok74_0s8wxk7wiu3hnx3w9l    ), 
  .mx7juirxj661i6i9lns4hnnyw0ep(vqixsqz3vz_o2ze5ovcwp577  ),

  .frehkmd0xqj4qeyqqodmp0onx7 (                        ),
  .ms95k2pmbvtrb33p5oa2q      (                        ),
  .r928tvy6d88uh6s9qun65udol2   (                        ),
  .jtgchf8072p4v1h9xclp0t  (                        ),
  .jekm9yqqqogc7_czwax0r6an_f  (                        ),
  .vs9f2qtmvyxt6ycc5e_z47fnjr (                        ),
  .wvywyxp28r9wdwncg13zbc_6    (                        ),
  .suaktr_howpmkqxx3p5j4      (                        ),

  .mnym6ha4fxtg2oqq9hlac5s1      (                    ),
  .p6wfurur4eut85r8tktdi03zxb   (                    ),
  .xxr9qx83ggzl9q98ig_ys5w60a  (                    ),
  .lozr9fiy6p7y8rinc582m2bt2ha_xmf  (                    ),
  .u78ade2idh660umk_1m66fdlksb9b  (                    ),
  .z3j5lbdgqwmp5zmv4g_zn29fgvintdc (                    ),

  .ussyj508sxu9v0           (jpplkccgktsmzedro78tuuvm8  ),
  .pdns51exd9ffhf5pykv42sq     (hnq2agjqmp3jnfvc02q9vn ),  
  .k09nslb_nkoy4r0t34xu6    (b04f0gnze13bj90dolndjwsij1e),
  .crr9jljkvi3gsixv1_v8       (),
  .sca7p0942a6kocjqqvat       (),
  .go_m73qp_w0p7abohs24       (),
  .jm4ru1fdiqtw706w8        (l_h0z16ew816k0kc59fz),
  .j021ufdslrlb4m5c5h2      (v1_i1c87etnhn8gl6t64rr),



  .p1kjflyurzeuxj (p1kjflyurzeuxj),
  .yvjlu1e9eng5_5tme (yvjlu1e9eng5_5tme),
  .hh8nc68zrpki2m9r (hh8nc68zrpki2m9r),
  .v8wv99vga5gkl8xhk7x9in (v8wv99vga5gkl8xhk7x9in),
  .ahfx5rs9jkdyw3b8ztscfx (ahfx5rs9jkdyw3b8ztscfx),
  .ts3_k4ergzh8upz7 (ts3_k4ergzh8upz7),
  .ktqya1x1mfi5j3q7 (ktqya1x1mfi5j3q7),
  .z6njhanl_m_hv48x5i9y (z6njhanl_m_hv48x5i9y),
  .dvm_h24fnflt11prmyvme (dvm_h24fnflt11prmyvme),
  .uvyubcp0tbk9yirhz (uvyubcp0tbk9yirhz),
  .ivoui15mvw3de5ds44 (ivoui15mvw3de5ds44),

  .gf33atgy          (gf33atgy),
  .ru_wi        (ru_wi)
  ); 


  wire y86fvwjf6k22ahfluzpt9; 
  wire q4gz66g470k0a1u_kk; 

  wire hraqlcavq96j53yrbyif;
  wire bf5ypgqi4grkg506x  ;

  wire flv4ybjx_fxnt8ahli; 
  wire mp50sb0x32pr82qg; 
  wire r1mbz1476mmd6eb_2gb;
  wire omlfl4p9_5zoeeas3; 
  wire p0e6oiwfprzmn8yx9hsoby9;
  wire [64-1:0] ue5tzeds4j8o5wx5zkx;
  wire i3fga9mifalr9g_siehz7127f4; 
  wire sd8rqg0mey7v6mthfjratzooccvk9;
  wire e0srj1jifo6i8ocnkw8xqhp  ; 
  wire ckrr5bi6ad3t5_60gouyjr9vvpfr;



  wire                       ypn14jlxvbvoxkesp;
  wire                       w70wabyhluyk3s21d4kaq;
  assign mgtrw760fgm5m362j     =  ie4dehipkb3b8__y5dt ? ypn14jlxvbvoxkesp : w70wabyhluyk3s21d4kaq;
  wire   x8j7zqt_iteyb74s7eq4w =  ie4dehipkb3b8__y5dt ? 1'b0         : jf9ko0etxomcrj25;
  wire   fl5uzx8oymfa        =  ie4dehipkb3b8__y5dt ? jf9ko0etxomcrj25 : 1'b0; 
  wire   q9d7ens0ettrow       =  ie4dehipkb3b8__y5dt ? tb198r6lzk1sr77g4 : 1'b0;
  wire [48-1:0] gyb1vfnsiaxnp  = {48{ie4dehipkb3b8__y5dt}} & gyxiq3yqdnanuqt16bh7r0h;



  wire f29yand0_mv30jc6grvj6;

  wire jgah5jfw;


tkyketfhrvq0gmush9p8_myoe xyckjo2h15upilfiwvu_jtc3q (


  .exltui35irvvmodu205vw(exltui35irvvmodu205vw),

  .vyxop00ua6vr(vyxop00ua6vr   ),  
  .p6rw9no76a3m  (p6rw9no76a3m   ),  
  .zowrmckfhx7k5    (pldoasxyzlvx2),
  .tvh1llq2i3_y  (tvh1llq2i3_y   ),  
  .hfsmpma3    (bde41te346q515l),

  .sxvvsxtbhyvt(sxvvsxtbhyvt),
  .azll7rq5fab5ou(azll7rq5fab5ou),
  .n6a0r_0zddzrme8(n6a0r_0zddzrme8),

  .pcr4upio7_tx37   (pcr4upio7_tx37   ), 
  .uzklqlncpqqm1rav(uzklqlncpqqm1rav),
  .ortueunvnkx_l5m_j(ortueunvnkx_l5m_j),
  .hwuhtb7ucto_utk56(hwuhtb7ucto_utk56),
  .i1env2kmns7qvvuuc(i1env2kmns7qvvuuc),
  .g3s3vpafvy3i(g3s3vpafvy3i),

  .rm1dxjejhq7dh3q5m(rm1dxjejhq7dh3q5m),
  .rvr30vvllni  (rvr30vvllni),
  .z1cj655u31  (z1cj655u31),



  .f29yand0_mv30jc6grvj6(f29yand0_mv30jc6grvj6), 



  .ibc9r3db5iet7          (zpg071p8a094ze4),
  .h7pglrrhtu6x34l5a21ern   (uh0wfy2udciats10exk7gx),

  
  
  
  
  
  
  
  
  
  
  
  
  
  

  
  
  
  
  

  
  
  
  
  .vs6ryzcr0bwqs5so          (vs6ryzcr0bwqs5so          ),
  .j25ub196dc_agl8oovaex4         (j25ub196dc_agl8oovaex4         ),
  .pi2nokcm8qf7och7l4g         (pi2nokcm8qf7och7l4g         ),
  .c0i0hs5tz64_ce5f0z        (c0i0hs5tz64_ce5f0z        ),
  .dmzdczrqcueolg3dzufj_by5rmf   (dmzdczrqcueolg3dzufj_by5rmf   ),
  .a1sqko6fok9qzpbtyuw0        (a1sqko6fok9qzpbtyuw0        ),
  .bquohubxiv2rsayn62v        (bquohubxiv2rsayn62v        ),
  .kqyojh1maxy0x834htg       (kqyojh1maxy0x834htg       ),


  
  
  
  
  .oa95jvzldxkjxnka5         (oa95jvzldxkjxnka5         ),
  .hjbzyjew4g2fmth4l66ng8        (hjbzyjew4g2fmth4l66ng8        ),
  .dl59edtk0_9k5jd65gxp        (dl59edtk0_9k5jd65gxp        ),
  .unzbnfwje52jxr_9yt38_bmn       (unzbnfwje52jxr_9yt38_bmn       ),
  .qtcuhd18j5hjtx41o9tjmv0cm434  (qtcuhd18j5hjtx41o9tjmv0cm434  ),
  .srphqbnx3w67orxkuwvoz       (srphqbnx3w67orxkuwvoz       ),
  .jbju6a9hecf_f8kg2bsz4       (jbju6a9hecf_f8kg2bsz4       ),
  .w66c528fqa9qnfz1btjnm      (w66c528fqa9qnfz1btjnm      ),






  .q9d7ens0ettrow(q9d7ens0ettrow), 
  .fl5uzx8oymfa(fl5uzx8oymfa), 
  .ypn14jlxvbvoxkesp(ypn14jlxvbvoxkesp), 

  .gyb1vfnsiaxnp(gyb1vfnsiaxnp),
  .elf4ijc6zyn02ua(pc67uztpd_zg6bsal),
  .ijrke0oayz6k (x2uw3xkpg8k47k8i ),
  .in937eccpoct (po0i9bzsw2yj9tv ),
  .kc2beprm1o1chr7jv (x967n2unm25k5336wf2 ),
  .zhfmvvqqyhe6l74(ucybeaa15_qx208e),

  .e28x1bh5rb6(cvvsn7xc8qg5uk),

  .scadliwzjp0l78srd9p    (ihlsip_az_gbdtb7cn43tr8wy),

  .o0gxucmy66th1ly2om5p      (jfnkyxema4_sqj5v2v),
  .wzqcq7ug3_gv3tuf0o       (j9pnp242pb8iiimxe87y),

  .hr0gt1i5t2qzoifxdtx3  (cgok74_0s8wxk7wiu3hnx3w9l  ), 
  .tnr82i_e_q5p_n4o9w2cp5(vqixsqz3vz_o2ze5ovcwp577),

  .n3zlo14nquu5l7zf3 (n3zlo14nquu5l7zf3),
  .a_1o1o8345o28hui    (a_1o1o8345o28hui  ),
  .t8p1kh0tvb2ej56s  (t8p1kh0tvb2ej56s),

  .y86fvwjf6k22ahfluzpt9 (y86fvwjf6k22ahfluzpt9), 
  .q4gz66g470k0a1u_kk (q4gz66g470k0a1u_kk), 

  .hraqlcavq96j53yrbyif(hraqlcavq96j53yrbyif),
  .bf5ypgqi4grkg506x  (bf5ypgqi4grkg506x  ),

  .flv4ybjx_fxnt8ahli(flv4ybjx_fxnt8ahli),
  .mp50sb0x32pr82qg     (mp50sb0x32pr82qg     ),
  .r1mbz1476mmd6eb_2gb  (r1mbz1476mmd6eb_2gb  ),
  .omlfl4p9_5zoeeas3 (omlfl4p9_5zoeeas3 ),
  .p0e6oiwfprzmn8yx9hsoby9(p0e6oiwfprzmn8yx9hsoby9),
  .ue5tzeds4j8o5wx5zkx (ue5tzeds4j8o5wx5zkx ),
  .i3fga9mifalr9g_siehz7127f4  (i3fga9mifalr9g_siehz7127f4  ), 
  .sd8rqg0mey7v6mthfjratzooccvk9(sd8rqg0mey7v6mthfjratzooccvk9),
  .e0srj1jifo6i8ocnkw8xqhp  (e0srj1jifo6i8ocnkw8xqhp  ), 
  .ckrr5bi6ad3t5_60gouyjr9vvpfr(ckrr5bi6ad3t5_60gouyjr9vvpfr),

  .an6zohwqn5kwj_tsi4_pczkvu (vdtkg4_jnsbu0p8wqnasmncdouhwmk),
  .bvvlopjoczq9r7vemdrzz3xd (dll7vburbug9zho0oh3rpr0pnjnnh),
  .yuloizdmigr7b94rp         (wqbvx_uqjrfzj8cjke712tpq),
  .c9k79dqw2z4f63_8lcp4w   (c9k79dqw2z4f63_8lcp4w),
  .u6f8hwzstewuo7nl0iywamw     (u6f8hwzstewuo7nl0iywamw),
  .o_4mw1alrjmdzl           (s47txxhzt1zertcfln5),
  .nkjxsm02z2_q5_0_         (w0s0l3_vvnnjgr_7cg2),








  .o21b8ypt1xiu5ml63d        (eyvp_wq1ero7byc8pxubqtg   ),
  .badsf4ksbp3k6p_p5hnj2i      (g0gwombfdn5ycvw4m1vh7f95 ),
  .ed4kcy8s9nrisftgx_q      (umtp4mg0svcx_tzytl9f2gx_9qa ),
  .bdqo1tgw2_bpi2e8alini       (ave0oxjdt4lz6czd61woyw2yb  ), 
  .jp5nha2l14e7kx2jzpke       (hc665sbb0domfwj0scqo_bhyan0  ), 
  .a4a48egkdkec8d9b_9      (ehzuy3rj6cnownydmlhhqorz ), 
  .xwfmltfzahuj4qfn4qf2      (a8hb7l400suw5vjdy40x_cjbtdzv ), 
  .ggxoqcj7ytp1a4pjf7ee       (rn2r2g1hhe3zfa2usi0x_mw  ),
  .oq9b5zfhza9yvdoj       (fcfcmwdw40u0wskca41p_6qb7m3  ),
  .l3c127qdc9a2mfc13      (gy3d5ed4dpwebmbht825jpu ),
  .zdpamqgv7ddf1n3x5t2q      (evt2fcz8mh_y8u4scgguyq287kcm ),
  .wpsukhyqhl92dzoam7cm      (wrqq_2zdqd0x7l_8uyy75putmx ),
  .v3oo69y614hgiemyyld      (f9gyp2oa2mz_rqxqxrizc1l ),
  .vy1zc0f0lrbzkonj3v     (srz_pttv795yabd3rlohv25jpcoj),
  .uxlldm0w_h7kicit8gvhqv2     (w9feuue3j76drwahit30vtv396w),
  .yvu98r_7ji4o250r_u         (caj02kz7j7ejw81vsf0fla    ),
  
  .szrgf24or2mbt7w_yleh_vt(szrgf24or2mbt7w_yleh_vt),





























  .l_giy79jkzkxy7j        (l_giy79jkzkxy7j ),
  .cw9xa748nw          (cw9xa748nw   ),
  .x1huhi29x9mco         (x1huhi29x9mco  ),
  .fpo04urqz74           (fpo04urqz74    ),
  .a2i6e7_7          (a2i6e7_7   ),
  .cque110xwd150_       (cque110xwd150_),
  .m705cbtazx7y        (m705cbtazx7y ),
  .etp831o_vh94        (etp831o_vh94 ),
  .w3p1po3pu         (w3p1po3pu  ),
  .nxy2oljfg0lssc        (nxy2oljfg0lssc ),
  .n2s7mr_zvl9k        (n2s7mr_zvl9k ),
  .mzwwsw0h6m1        (mzwwsw0h6m1 ),
  .lydg_n0cr655       (lydg_n0cr655),
  .tb62wswspbytv       (tb62wswspbytv),
  .jttn_e63nm4n4lm9       (jttn_e63nm4n4lm9), 

  .yixt0a_xmh    (yixt0a_xmh), 
  .ej7frm_ut9j6y(ej7frm_ut9j6y), 
  .izjeme5aukvcc(izjeme5aukvcc), 
  .x5nbgu5ggtet3   (jgah5jfw     ), 

  .ttgsydregi0kgoj_z(mne0dg23_1aal06pio[64-1:0]), 

  .dw0ku_p4sgs3627wdlt6 (tcveomov4rt0zai5ns),
  .ygvgcd3cyi2ipiz53hbsp   (ygvgcd3cyi2ipiz53hbsp),

  .gf33atgy  (gf33atgy  ),
  .ru_wi(ru_wi)

);








xqy0kx72ozzh4s06ej rfbxpg_a_jvq33y4tma8b4k (

  .sxvvsxtbhyvt  (sxvvsxtbhyvt),

  
  
  
  
  
  
                            
  .rm1dxjejhq7dh3q5m              (rm1dxjejhq7dh3q5m              ),
  .rvr30vvllni                (rvr30vvllni                ),
  .oa95jvzldxkjxnka5         (oa95jvzldxkjxnka5         ),
  .hjbzyjew4g2fmth4l66ng8        (hjbzyjew4g2fmth4l66ng8        ),
  .dl59edtk0_9k5jd65gxp        (dl59edtk0_9k5jd65gxp        ),
  .unzbnfwje52jxr_9yt38_bmn       (unzbnfwje52jxr_9yt38_bmn       ),
  .qtcuhd18j5hjtx41o9tjmv0cm434  (qtcuhd18j5hjtx41o9tjmv0cm434  ),
  .srphqbnx3w67orxkuwvoz       (srphqbnx3w67orxkuwvoz       ),
  .jbju6a9hecf_f8kg2bsz4       (jbju6a9hecf_f8kg2bsz4       ),
  .w66c528fqa9qnfz1btjnm      (w66c528fqa9qnfz1btjnm      ),
  
  
  
  


  .st2zalpx0uf (st2zalpx0uf), 
  .ni01kj42oob2x (ni01kj42oob2x), 
  .ah8kjlmvnaxzbi (ah8kjlmvnaxzbi), 
  .w30ye15yns15    (w30ye15yns15),
  .vdtkg4_jnsbu0p8wqnasmncdouhwmk       (vdtkg4_jnsbu0p8wqnasmncdouhwmk),
  .wqbvx_uqjrfzj8cjke712tpq               (wqbvx_uqjrfzj8cjke712tpq), 
  .dll7vburbug9zho0oh3rpr0pnjnnh       (dll7vburbug9zho0oh3rpr0pnjnnh),
  .evji0n54bi8hm_n24uk853qw9c         (evji0n54bi8hm_n24uk853qw9c       ),       
  .s9psy03yyyxh7qrmosmb1                (s9psy03yyyxh7qrmosmb1              ),               
  .sqkbogq1h4psprgoosl2lmrpj9_         (sqkbogq1h4psprgoosl2lmrpj9_       ),
  .n5gj_lxl9078ky9b2zawd0             (n5gj_lxl9078ky9b2zawd0           ),
  .b0fkq6hghv6az5l_j1j2c12imdd6          (b0fkq6hghv6az5l_j1j2c12imdd6        ),         
  .argq10f3h723e0jtlrdbu53               (argq10f3h723e0jtlrdbu53             ),              
  .e7iar94ylidlt25a9g9n               (e7iar94ylidlt25a9g9n             ),              
  .qj6kqe1holct34gfb0q9p9a04_alrzg         (qj6kqe1holct34gfb0q9p9a04_alrzg       ),                        
  .bmkssziw1_8am7ea6dv                 (bmkssziw1_8am7ea6dv               ),
  .xefc2nul9m648jueckdrui_l             (xefc2nul9m648jueckdrui_l           ),
  .woq47beoqkpu1um82nv58l1u_hyj4         (woq47beoqkpu1um82nv58l1u_hyj4       ),       
  .a1r66jlym5w100htq8lfn_o0rapdf5s      (a1r66jlym5w100htq8lfn_o0rapdf5s    ),    
  .trt0bnwhmoe0r7apy2x_p9hltd           (trt0bnwhmoe0r7apy2x_p9hltd         ),         
  .wqjorkypks0nndgahingvyvil3dvqo          (wqjorkypks0nndgahingvyvil3dvqo        ),        
  .obokll126527kg6wlw1t6vfh8          (obokll126527kg6wlw1t6vfh8        ),        
  .msh4030y2dhqf78kyckys0c2ue0ic          (msh4030y2dhqf78kyckys0c2ue0ic        ),        
  .oebo4piph5o2byr1030bgmb0ye31c6          (oebo4piph5o2byr1030bgmb0ye31c6        ),        
  .tlmtrlht_1gsijvzms1twiewyym          (tlmtrlht_1gsijvzms1twiewyym        ),        
  .ez_fxjs3_wlsve__62ua9tqsfa6k89twfir    (ez_fxjs3_wlsve__62ua9tqsfa6k89twfir  ),  
  .p3nsxkqv6seglstz4ge77tdjcngbig0w30rq  (p3nsxkqv6seglstz4ge77tdjcngbig0w30rq),


    .xhpc6eofokpbnya1h3s117_2  (umtp4mg0svcx_tzytl9f2gx_9qa ),
    .badsf4ksbp3k6p_p5hnj2i      (g0gwombfdn5ycvw4m1vh7f95 ),
    .ed4kcy8s9nrisftgx_q      (umtp4mg0svcx_tzytl9f2gx_9qa ),
    .bdqo1tgw2_bpi2e8alini       (ave0oxjdt4lz6czd61woyw2yb  ), 
    .jp5nha2l14e7kx2jzpke       (hc665sbb0domfwj0scqo_bhyan0  ), 
    .a4a48egkdkec8d9b_9      (ehzuy3rj6cnownydmlhhqorz ), 
    .xwfmltfzahuj4qfn4qf2      (a8hb7l400suw5vjdy40x_cjbtdzv ), 
    .ggxoqcj7ytp1a4pjf7ee       (rn2r2g1hhe3zfa2usi0x_mw  ),
    .oq9b5zfhza9yvdoj       (fcfcmwdw40u0wskca41p_6qb7m3  ),
    .l3c127qdc9a2mfc13      (gy3d5ed4dpwebmbht825jpu ),
    .zdpamqgv7ddf1n3x5t2q      (evt2fcz8mh_y8u4scgguyq287kcm ),
    .wpsukhyqhl92dzoam7cm      (wrqq_2zdqd0x7l_8uyy75putmx ),
    .v3oo69y614hgiemyyld      (f9gyp2oa2mz_rqxqxrizc1l ),
    .vy1zc0f0lrbzkonj3v     (srz_pttv795yabd3rlohv25jpcoj),
    .uxlldm0w_h7kicit8gvhqv2     (w9feuue3j76drwahit30vtv396w),
    .yvu98r_7ji4o250r_u         (caj02kz7j7ejw81vsf0fla    ),
    .o21b8ypt1xiu5ml63d        (eyvp_wq1ero7byc8pxubqtg   ),

    .l_giy79jkzkxy7j        (l_giy79jkzkxy7j ),
    .cw9xa748nw          (cw9xa748nw   ),
    .x1huhi29x9mco         (x1huhi29x9mco  ),
    .fpo04urqz74           (fpo04urqz74    ),
    .a2i6e7_7          (a2i6e7_7   ),
    .cque110xwd150_       (cque110xwd150_),
    .m705cbtazx7y        (m705cbtazx7y ),
    .etp831o_vh94        (etp831o_vh94 ),
    .w3p1po3pu         (w3p1po3pu  ),
    .nxy2oljfg0lssc        (nxy2oljfg0lssc ),
    .n2s7mr_zvl9k        (n2s7mr_zvl9k ),
    .mzwwsw0h6m1        (mzwwsw0h6m1 ),
    .lydg_n0cr655       (lydg_n0cr655),
    .tb62wswspbytv       (tb62wswspbytv),
    .jttn_e63nm4n4lm9       (jttn_e63nm4n4lm9),

    .jgah5jfw           (jgah5jfw    ), 

    .xmbe_e4vm6ofjbn7lq    (xmbe_e4vm6ofjbn7lq),

    .aht5xalx865dt9ymg6t4    (badsf4ksbp3k6p_p5hnj2i   ),
    .zjmbnwsbyle24ayly67    (ed4kcy8s9nrisftgx_q   ),
    .icfwo5l56zab795f     (bdqo1tgw2_bpi2e8alini    ), 
    .n78yvkhg0miifi58     (jp5nha2l14e7kx2jzpke    ), 
    .wu02k99r_ok2kjj4u119us    (a4a48egkdkec8d9b_9   ), 
    .ccwk4o03vlem_hqcccf1g6    (xwfmltfzahuj4qfn4qf2   ), 
    .yx2bhxvyxmxjggxrsrr833 (p648zxn2luyxy8mt992a), 
    .qe64ftxd03f_vqrd2sd     (za9xg3zsqni_aeqmke    ),
    .b36sriu021vdo_ujif8     (c1gmncmorg16sachdas    ),
    .ltx9lurd9p2ivmnufrgrw     (ggxoqcj7ytp1a4pjf7ee    ),
    .o1gawztvzi0onzitk     (oq9b5zfhza9yvdoj    ),
    .lr02cqs6anj9gvr45kv    (l3c127qdc9a2mfc13   ),
    .z6ncd60zcel8m99zg6v    (zdpamqgv7ddf1n3x5t2q   ),
    .st9_is6howar7iysonyyhk    (wpsukhyqhl92dzoam7cm   ),
    .o8407eu9fhzcuymr2a4    (v3oo69y614hgiemyyld   ),
    .t3ubula_wguy1a2tut1_e   (),
    .ukl6eat4ng6xala4y597l2i   (uxlldm0w_h7kicit8gvhqv2  ),
    .w3yoivbzacxwr95dw       (yvu98r_7ji4o250r_u  ),
    .qsw59ks9jxcsmmh      (o21b8ypt1xiu5ml63d     ),
                          
    .s4dz24kz7cxir4hxtt   (flcopog5zzpohfautwy   ),
    .epoc75xqnuvcqziu_9i55h   (gtb8f_h0g28itdr8k   ),
    .w0vagcfu1v7wkym9f     (wf15djwi2hw25nz_     ),
    .sjx2nupt4_7eb6_metse (t1q5qmk9jzpf6glng4y ),
    .gxo5tf4bea2gsq4yyn   (xsmx4zoewhbt07jxq   ),

    .jugi02ecegnos3        (qhvzepznvxpv9_wyiu767h7      ),    
    .rxjuugktc38un        (lwjhzma3f8s38cp0iw7a471x      ),
    .h8wu7unf_ixmxfeh         (kcliouozy4gzxf4ji1d_1ug       ),
    .kdpgigzs75vcc1d         (t208_ksfx0p48awxbbi41vdc6k       ),   
    .coohnlu_ri          (p6887dnv76xwdpql2ru4c        ),   
    .x6uy7s6mcepqq2j527jtxk   (lkdi90h27rm6bstdc_lv43xs9hw ),   
    .igo49dpz9ealh4h13a   (p1todm057e8_laqnquniw6y0rw6 ),   
    .ks33bi5hojtg0te9bl7   (uvbcza18x9h661vyy9t1uik595c ),   
    .dwet7q3ucodidho7qxlw  (ff37q45o11p27pc_tlfpgr8yspb0w),  
    .p_p6yt19xmgqbfsn0y       (bv8onmahmkg35l9opjmw5v1axpaj),   
    .k5h5ux92dlz_nn0       (d_arhdx13m6c57bz_fusjchynkad     ),   
    .e6uinbhqc8o7iylg7d    (vx75xcy7pymxftm_8zyk4pytv9kuyd     ),  

    .j2_lz0mpsxf4xotgqf1ngx   (j2_lz0mpsxf4xotgqf1ngx),
    .hcugdkhp9szims1nk8rhakn(hcugdkhp9szims1nk8rhakn),
    .dw2ygdedledlm7ps830qgbwonu(dw2ygdedledlm7ps830qgbwonu), 

    .ygvgcd3cyi2ipiz53hbsp   (ygvgcd3cyi2ipiz53hbsp),

    .gf33atgy                 (gf33atgy),
    .ru_wi               (ru_wi)

);


assign sg33s7pt45jp_ = hcugdkhp9szims1nk8rhakn;


  wire no7xdtjyy1_rzn5 = af5qc04tmn51e4u2h1z 
                          & jgah5jfw & jp5nha2l14e7kx2jzpke
                          & (badsf4ksbp3k6p_p5hnj2i & ed4kcy8s9nrisftgx_q)
                          ;











assign hey6uxy22wzzlom6mekyg2y = {1'b0,y3lf5lq_1tfm1iea};
assign qerr94cedlotaj08239y = zcl5hta0nld; 
wire   hhx3zl7wc_kiw7l = d9_s5e6qdqa7haet4s & zh907qs92c1ixb_97gmdepk;   

  kho7cvkwdsu6ed90f6_18aax2 #(
    .xio4kx7ep1ojwa_r     (55),
    .cmnocc9r2aiw8za      (8 ),
    .xholqktr732apzsv8d0 (3 )
  ) rdmhx1mfymki4grjbn1w3eqc0 (
    .es6_9ffb14edb7t                     (hhx3zl7wc_kiw7l                   ),  
    .mv5to8v6                          (kvpemhoim1tq5y8mzwvix5              ),  
    .zh907qs92c1ixb_97gmdepk             (zh907qs92c1ixb_97gmdepk             ),
    .phofig8d5zd_8v9g8                    (phofig8d5zd_8v9g8                    ),
    .hey6uxy22wzzlom6mekyg2y             (hey6uxy22wzzlom6mekyg2y             ),
    .qerr94cedlotaj08239y                 (qerr94cedlotaj08239y                 ),
    .js0ml55dtie8qenb4eoj2              (js0ml55dtie8qenb4eoj2              ),
    .ticm3jrqt6tjtf6                   (ticm3jrqt6tjtf6                   ),
    .hpaul9bznamp4qkl                   (hpaul9bznamp4qkl                   ),
    .vq7jwn83uus_ac4s4ghf             (vq7jwn83uus_ac4s4ghf             ),
    .gzh3us4_ux10aey                     (gzh3us4_ux10aey                     ),
    .np3fnkgbpsuf8nkgnf                 (np3fnkgbpsuf8nkgnf                 ),
    .evji0n54bi8hm_n24uk853qw9c       (evji0n54bi8hm_n24uk853qw9c       ),
    .s9psy03yyyxh7qrmosmb1              (s9psy03yyyxh7qrmosmb1              ),
    .sqkbogq1h4psprgoosl2lmrpj9_       (sqkbogq1h4psprgoosl2lmrpj9_       ),
    .n5gj_lxl9078ky9b2zawd0           (n5gj_lxl9078ky9b2zawd0           ),
    .b0fkq6hghv6az5l_j1j2c12imdd6        (b0fkq6hghv6az5l_j1j2c12imdd6        ),
    .argq10f3h723e0jtlrdbu53             (argq10f3h723e0jtlrdbu53             ),
    .e7iar94ylidlt25a9g9n             (e7iar94ylidlt25a9g9n             ),
    .qj6kqe1holct34gfb0q9p9a04_alrzg       (qj6kqe1holct34gfb0q9p9a04_alrzg       ),
    .bmkssziw1_8am7ea6dv               (bmkssziw1_8am7ea6dv               ),
    .xefc2nul9m648jueckdrui_l           (xefc2nul9m648jueckdrui_l           ),
    .hpk3eafyque5ubt_c62flnny            (hpk3eafyque5ubt_c62flnny            ),       
    .sfezv1xz2ghvo8pkt                   (sfezv1xz2ghvo8pkt                   ),               
    .vagaza053272juvmo59v8w20s            (vagaza053272juvmo59v8w20s            ),       
    .rzf45534z36ejq96260                (rzf45534z36ejq96260                ),       
    .frzfsbt7hp3n4aj3zvvumnh0s             (frzfsbt7hp3n4aj3zvvumnh0s             ),         
    .zkuxqezrmlhyyjjgx                  (zkuxqezrmlhyyjjgx                  ),              
    .u3h5tvu1g2q93141j9o                  (u3h5tvu1g2q93141j9o                  ),              
    .pjh0wad7t_5du3cync_0c            (pjh0wad7t_5du3cync_0c            ),                        
    .wmkgrgf631pbq                    (wmkgrgf631pbq                    ),
    .oyq1p3qa2iffjuqns0jkgg                (oyq1p3qa2iffjuqns0jkgg                ),
    .c9k79dqw2z4f63_8lcp4w             (c9k79dqw2z4f63_8lcp4w             ),
    .ly39gmn8_bufgxi162s47mj5md          (ly39gmn8_bufgxi162s47mj5md          ),
    .u6f8hwzstewuo7nl0iywamw               (u6f8hwzstewuo7nl0iywamw               ),
    .owio9cfz6lmpk7katn_gtlo9              (owio9cfz6lmpk7katn_gtlo9              ),
    .dna64e9sa3ona8c40stq              (dna64e9sa3ona8c40stq              ),
    .yqonk7rjhe328d_deg1              (yqonk7rjhe328d_deg1              ),
    .fvuwaqmgv_r72l8z4ys0lq59              (fvuwaqmgv_r72l8z4ys0lq59              ),
    .x5_495u23v2cqjqs7nx9m3s              (x5_495u23v2cqjqs7nx9m3s              ),
    .qvfjqeg7co1udtegoqx2t09jmc        (qvfjqeg7co1udtegoqx2t09jmc        ),
    .m6_yvtzjevmj_c4bel_9vu0kkk_t      (m6_yvtzjevmj_c4bel_9vu0kkk_t      ),
    .woq47beoqkpu1um82nv58l1u_hyj4       (woq47beoqkpu1um82nv58l1u_hyj4       ),
    .a1r66jlym5w100htq8lfn_o0rapdf5s    (a1r66jlym5w100htq8lfn_o0rapdf5s    ),
    .trt0bnwhmoe0r7apy2x_p9hltd         (trt0bnwhmoe0r7apy2x_p9hltd         ),
    .wqjorkypks0nndgahingvyvil3dvqo        (wqjorkypks0nndgahingvyvil3dvqo        ),
    .obokll126527kg6wlw1t6vfh8        (obokll126527kg6wlw1t6vfh8        ),
    .msh4030y2dhqf78kyckys0c2ue0ic        (msh4030y2dhqf78kyckys0c2ue0ic        ),
    .oebo4piph5o2byr1030bgmb0ye31c6        (oebo4piph5o2byr1030bgmb0ye31c6        ),
    .tlmtrlht_1gsijvzms1twiewyym        (tlmtrlht_1gsijvzms1twiewyym        ),
    .ez_fxjs3_wlsve__62ua9tqsfa6k89twfir  (ez_fxjs3_wlsve__62ua9tqsfa6k89twfir  ),
    .p3nsxkqv6seglstz4ge77tdjcngbig0w30rq(p3nsxkqv6seglstz4ge77tdjcngbig0w30rq),
    .qjw2q0j88rjr42lautsqnca            (qjw2q0j88rjr42lautsqnca            ),       
    .imkm56ujne9v4m6n08w1yf5622         (imkm56ujne9v4m6n08w1yf5622         ),     
    .txk1r9aiq_7l2nkw101w_              (txk1r9aiq_7l2nkw101w_              ),          
    .ih4hmwugasiodbx5da9_40kx             (ih4hmwugasiodbx5da9_40kx             ),        
    .x5vjq7mshfwr0h3q514t7mhdt             (x5vjq7mshfwr0h3q514t7mhdt             ),        
    .qrxtk7e03100_uwkx73sg7             (qrxtk7e03100_uwkx73sg7             ),        
    .i7qiq2q9c6hbeful9qu9lb             (i7qiq2q9c6hbeful9qu9lb             ),         
    .yr0s3skqk7cdqflsrbsxg9znu             (yr0s3skqk7cdqflsrbsxg9znu             ),         
    .adqieke11qo0elfz93hlouwjc0       (adqieke11qo0elfz93hlouwjc0       ),   
    .w93gdpnnxuydy53eu0s9nxw7xdct7     (w93gdpnnxuydy53eu0s9nxw7xdct7     ), 
    .v66ux9ovjkzt3jn                   (bz8qao4o4xqslni1d3               ),
    .cd3lo77nievm4v3                    (vpecdc5kos                       ),
    .rgnht1zljy67subvhyua_             (pccd7o463jfc_dpc5va                ),
    .uy22rssg5uc6vyiti9szp                 (deo3wn_907tw886r                  ),
    .h8djzt4zbmppcv2_ai                  (k5ovx8tintgvetip                     ),
    .nmlix317bu48vgct7x02m7vgn             (f97le_hyejv7saw9vslna                ),
    .s6zb15tq6xjiqgce5nwjcg7be4        (yruel3nusosm39gnmb9ev_               ),
    .ry0rypry86op3l_hqbwk8pe32ena3e      (oeux55k_cre0he7w7jip5b1             ),
    .h4zmq2srkdf5iaeagd8d7i87              (r8z2r_ud53zj8mrpk                ),
    .dzo70vq3_1_kyxyiurxy1d20ed            (bu1949pq_9946o1_e2q_uvr8p4          ),
    .b0c0o6unssb9h3tgqck870            (b4isf5u8b8pj34e09f72vxe38zg          ),
    .dlygovkaje808pt5_j                   (e2rgt3d7pxx8bv6_w1v7                  ),
    .c2_546oy8pb0vifo                  (refz65mt7g99f_cb9h                 ),
    .gf33atgy                              (gf33atgy                              ),
    .ru_wi                            (ru_wi                            ),
    .gc4b3kdcan6do88ta_                   (gc4b3kdcan6do88ta_                   )

);




wire   brjte07eirv05n2q      = yd1xmujxb33j01a4c;
assign d6ltnbdw_4ll2          = o8rffdg1904azl0q && f0ziihie9il3138m;
assign lmrvfbh6ipddvrrollz4_   = np3fnkgbpsuf8nkgnf || fa9nldm69zre__ccuu82h;
assign zh907qs92c1ixb_97gmdepk = snxyhe6q4j0ik6is && d6ltnbdw_4ll2 && !fa9nldm69zre__ccuu82h && !brjte07eirv05n2q;  
assign fa9nldm69zre__ccuu82h     =     ~fkuqlh34r                                                
                              || ( aw82i964do && !rm1dxjejhq7dh3q5m)                                 
                              || ( aw82i964do && (st2zalpx0uf == 2'b11))                        
                              || (zcl5hta0nld && !(sxvvsxtbhyvt && rm1dxjejhq7dh3q5m) )            
                              || (zcl5hta0nld && !(sxvvsxtbhyvt && (st2zalpx0uf == 2'b11)) )  
                              ;
ux607_gnrl_dfflr #(1) b31uig740s4bms8knt_r7b48 (d6ltnbdw_4ll2,fa9nldm69zre__ccuu82h,jfnkyxema4_sqj5v2v,gf33atgy,ru_wi);







  cqpjxz2qb247thego6htwvkw_aiu lpcbtkgnuc86ae4xr8g1d9jqhojv_j(
  .f_8ecse5wf0jrndlozy2070bja                       (c9k79dqw2z4f63_8lcp4w       ),        
  .e4sprh35cvfb6sw6lnskyaga91                    (ly39gmn8_bufgxi162s47mj5md    ),
  .qrvtg_49_dmoggu94orq0                        (owio9cfz6lmpk7katn_gtlo9        ),         
  .iocew24g1qos_gvi3_r3uoqfdf                        (dna64e9sa3ona8c40stq        ),         
  .qh_y92pv7dp1us9t5wxdmm57                        (yqonk7rjhe328d_deg1        ),         
  .cznjry8adajzgi6gkmyr830m_u                        (fvuwaqmgv_r72l8z4ys0lq59        ),         
  .ugixcggahb26m1glzpuqvpq                        (x5_495u23v2cqjqs7nx9m3s        ),         
  .vbpz6tidsg3o93kih6nmamlyg9wmr1zz                  (qvfjqeg7co1udtegoqx2t09jmc  ),   
  .j2dtuvq0m4iir947lery9tpxqwhjj2g3                (m6_yvtzjevmj_c4bel_9vu0kkk_t), 
  .wzqcq7ug3_gv3tuf0o                           (j9pnp242pb8iiimxe87y),
  .ng5gq72xr47fw8fztwfo8hw                         (rm1dxjejhq7dh3q5m ), 
  .cmyy3ooatm0bn2s6fv8_r                          (st2zalpx0uf ), 
  .ckgybqpbvuzwgxv1ixd_6rpf                          (ni01kj42oob2x ),
  .nguthky_k_yqsf8fa9btry1                          (ah8kjlmvnaxzbi ),
  .w30ye15yns15                                     (w30ye15yns15 ),
  .jyl_xsaj6z1u9wndwpi                               (sxvvsxtbhyvt ),
  .idg19n7mm21jtb                                  (x967n2unm25k5336wf2 ),
  .o_4mw1alrjmdzl                                 (s47txxhzt1zertcfln5),
  .nkjxsm02z2_q5_0_                               (w0s0l3_vvnnjgr_7cg2),
  .gf33atgy                                          (gf33atgy),
  .ru_wi                                        (ru_wi)
);








  wire [64-1:0]          v_t46_oqiae0c4es9uht        ;
  wire [64-1:0]          xw9obr7t22kfov7grph7        ;

  wire                           apf9b6zz11802cqi      ;
  wire                           trff4kgfudc86mj      ;
  wire                           ooadt7528tbax93myw      ;
  wire                           qx67s81zzlmp_0y3     ;
  wire                           hmu_zk66odn2umlzrf0     ;
  wire                           z9601_tn67y_68ndtufn9     ;

  wire                           aykpj7s87z_wdrbcx0hx  ;
  wire                           f1k1tltm39p_5uxhp5l80q4  ;
  wire                           vztmqpg2g1jegcsjy       ;
  wire                           ztrmt5hqf4t_572v6d0p      ;
  wire [64-1:0]          mhwy3r0_oj3dwbbkxci        ;
  wire [64-1:0]          ktexyfhmd3f6j0oghmg        ;
  wire [64-1:0]          imkdfcjp0n3752tqx        ;
  wire                           o88kin60h043_xvw1jjqkq    ;
  wire                           mg3fx2urlykksnscs_7t0    ;
  wire                           clqozm1jbmldowubnqirw     ;
  wire                           yhtdgk1ljckfa3gybu4ofkrm9 ;
  wire                           ysh2g3tr4jy_ogbn47v1     ;
  wire                           kf_d85407aznl0ii     ;
  wire                           dm23tkdzwq_nstqh7q   ;
  wire                           r1upbgyfw2ogtmd_      ;
  wire                           c_2htc3ogchp6l1b_ocaywwd  ;
  wire [64-1:0]          mq4z316n9yhcwtvfe        ;
  wire [64-1:0]          hiqrrqluaq93akcapxdylg    ;
  wire [48-1:0] pa6s_tjxpy4gq16f7iur7   ;
  wire                           ix1bi23f1mg6sekjqzl     ;
  wire                           jwsf_7nftft_w24ca     ;
  wire                           mqkvwvl8pflc9cluk      ;
  wire                           seo11tmtq27hed2p      ;
  wire                           mtuge6clzfy0w9er3      ;
  wire                           lvi1vea5zurx7sli3iif74  ;
  wire                           tbuth82v2mm2g7uok_hiph  ;
  wire    [4-1:0]    anj5c56sztftipab3_sfkos7yi;
  wire    [4-1:0]    l0z8mly9ui8x1u5ulfb4walt6;

  wire [64-1:0]       j3zy8mipfns_ki;
  wire [32-1:0]    xls7sq397kcp2;
  wire [64-1:0]       eemxwz9vo25r4djt76yzhab1ue;
  wire                           gsmurqtk28c99urfc3mhf1804;

  wire [64-1:0]       oungyftsa5o1qeiq0zbvzw5f;
  wire                           xckbb1f5bxl8d6iqjh7et8uce;
  wire                           b39373uuxt1fwwvp8c2yhm;
  wire  [64-1:0]      qm7esy9r83ecuoam3onh6tm;
  wire                           dclg9gzyeu9de8scca2r66;

  wire                           ak3_rgqx75eo7s2jfbhemwqz8ng ; 
  wire                           hbinkk7e8nmokz2d2dm9gq2j82r;
  wire                           y6zepdb9e4svr2kxsxig3dej9  ;
  wire                           leq1ne49igptrh__p_5kz23048rjzm ;
  wire                           ipj0pyjf76qkv519em1jiaiutbhsr ;
  wire                           szaorjzmus1ssgjq7e30bdssuadwt0 ;
  wire                           yi0r5xirgktqhr99j3jz345g11t51 ;
  wire                           ogkluwmj9mmpgtmicjnh6_yya46ukkp2s;
  wire [64 -1:0]         d250junaig195xflrdmkjjl5pxtaf4;
  wire                           unntlrmfpzgdq8rnz3ug3_8 = vx75xcy7pymxftm_8zyk4pytv9kuyd;
  wire                           gkjb6c98b5j1zsgbv26  = d_arhdx13m6c57bz_fusjchynkad;
  wire                           n9q1kib2q28tfyzyue2j2or = lkdi90h27rm6bstdc_lv43xs9hw & ygvgcd3cyi2ipiz53hbsp;
  wire                           asxvrob6s2_85u99em22 = p1todm057e8_laqnquniw6y0rw6 & ygvgcd3cyi2ipiz53hbsp;
  wire                           bva3_s2oj2hgomj0eyrk = uvbcza18x9h661vyy9t1uik595c & ygvgcd3cyi2ipiz53hbsp;
  wire [64 -1:0]         fbgda1d6z8gr725snyc2ylc = ff37q45o11p27pc_tlfpgr8yspb0w;



  wire lhs982qsuxsw7i76wzs9;
  wire er1ax0dpgq0b7g6i = y86fvwjf6k22ahfluzpt9 | x8j7zqt_iteyb74s7eq4w;
  wire [64-1:0] s27lb72llmh3g7i6uu = qhvzepznvxpv9_wyiu767h7 ? kcliouozy4gzxf4ji1d_1ug : mne0dg23_1aal06pio;

  assign w70wabyhluyk3s21d4kaq = lhs982qsuxsw7i76wzs9; 


  assign q4gz66g470k0a1u_kk  = lhs982qsuxsw7i76wzs9;
  assign lwjhzma3f8s38cp0iw7a471x = lhs982qsuxsw7i76wzs9;

  wire tpd5fcgyg_240nz8md69oj  ;
  wire npkoy9e2dsczayfq7h6cko59;
  wire kmlf0ops49wvgcz2howfob59khsqir  ;
  wire kw590mop2ic8u619z7c_owrnv9t;

  wire                       oa_1ibjpvwpv6bg5ivcau2uo6z3s;
  wire                       noc4nf4qform41kyqw6m4     ;
  wire                       ktqyocabrct3iqhlj18u9fhnz6f3d  ;
  wire                       ihbxqlci_5lmn6uyuoxv158n18bua ;
  wire                       xv9g6nf92837e31mav06v03y2t ;
  wire [64-1:0] ppwfzi9r2pfdu5oiww3x5a9g94u6ut0;
  wire                       by0pbwftr5xjmht8u5rapxeyd1g ;
  wire                       z3m510kw9uow1_jbl0xi6lrg   ;



  wire                                   woqfe5v065k3eom51g4h1jq;
  wire [19-1:0]  x6s44jsh488qbnj6v9ppkpceb;
  wire [64-1:0]                  d228vs4sizjmlag0hkfk;
  wire [64-1:0]                  wz4he34y3_e1ieaudx5sv;
  wire [64-1:0]                  r2mcos1t0vvp47i3ka_vsc_;

  wire sdil6s1uzxtjt_viwt;
  wire ik7kganikfrfc8z_c;
  wire v9o_kfa70i0fkql780cet087h389;
  
  wire z492i2r2osjb1wm_z8kg_vzs;
  wire svrztr5zqc119uyafi4qw0w8e;
  wire [64-1:0]  vlpn6saddwb42teg;
  wire [64-1:0]  m3kk01rml527m1oq0v;
  wire [64-1:0]  d0g9hx2h2bufn9qst9s;



  assign zv7y8twrabykb59a8a4629 = ie4dehipkb3b8__y5dt  && !ygvgcd3cyi2ipiz53hbsp; 

  wire  zhfhfu89sj5v_ci5gp96ysg = icczfaorqi6bmvsm5c4h | (ie4dehipkb3b8__y5dt && ygvgcd3cyi2ipiz53hbsp); 
  
  
  wire  f09gaw2v2ppnj18jqy1n_ = (ie4dehipkb3b8__y5dt & ygvgcd3cyi2ipiz53hbsp) ? (sfrkf5j74_e8qi ? (hc665sbb0domfwj0scqo_bhyan0 & ~p6887dnv76xwdpql2ru4c) : (id6e2963yn91s9_9_5on & ~p6887dnv76xwdpql2ru4c)) : id6e2963yn91s9_9_5on; 


 assign nb2chelz4_ijwumv9murokla = qx67s81zzlmp_0y3;
 assign bcrcin74qehflgu36ch9ghyv = hmu_zk66odn2umlzrf0;
 assign fbzipldpa3ewvv31mgr = z9601_tn67y_68ndtufn9;



b0gv4gv3sqckul0vbemwxr#(
  .gdctpuyrfi_b (1),
  .l_7qc0w_2x6i(0),
  .t5462hhws9i6ynbxi(2)
  ) d6o_els12pvrpum2m(
  .cu1owrury8wsed               ({4{1'b0}}   ),
  .mt1z8r_sz               ({4{1'b0}}       ),
  .uc9k3lw_iehx               (fs6jojwsl0l32t7brm38vh   ),
  .radwr7skyhm3jqso5         (ydtm1yuxqj7fmxvqc    ),
  .zdid44qi3bv7q4phl         ({4{1'b0}}  ),
  .x4owqbu74zh_xxr         (eo5skx1ygvzuasbjgnyl    ),

  .b43m7n67rav8he           (1'b0      ),
  .qcutfgh43gov5u4urt           (1'b0  ),
  .s73raoa0ilom1wyi           (qd5sbh8mupp_n4y95vo  ),
  .dnwb40nhmse7rcj0epzjo     (vz63qkw5s3m8urb9       ),
  .omeribg0gbgvpn78urilv_a     (1'b0),
  .jxogr1vy8jotyh8ivd2u     (p1jdw9loxkz60taq_vkp_3       ),

  .kl8zh4diafqs                ({64{1'b0}}    ), 
  .jiartjoiycj2                ({64{1'b0}}   ), 
  .dtypmpwq1q2j                (s7vgjm2azmcc3uzzdc_7   ), 
  .uwl7jm0d1lv0xpo            (1'b0 ), 
  .u2l80pdclhyu1bl            (1'b0 ), 
  .uamf3ccv7ouhi18            (1'b1        ), 
  .pkw60eo867gghh          (iojqlhtwx45_siz         ), 
  .strg8286lgex8p4_0m          ( {64{1'b0}}), 
  .avpvrch0prpui67          (jwwku_el5h5h2lx6e0kyi ), 


  .plk8ixck4wj7c          (s27lb72llmh3g7i6uu ), 
  .e7nqb0p7cffw4lrkd        (bq9gnoi981qw397qkojrj),
  .dorqi70cvs05s       (nw1d2c3l16ufwicfgjc),
  .pgfbjdj832ly_       (gtuyw8lwe5vig3whpwia),
  .z0yti764_a15nwanb       (bepi9gxgibkbsjimgygx),
  .k5yu5na0oo41y       (pjybabc2ndhp9w15),
  .n8g2a10i7cbowtvjhc       (r8n4jj_yqo_psdycdpf),
  .pzlsmt96uolwfb47           (rc1qjhv_cq1wdp4lltk8               ),
  .uzn8ik3rkkwib6p           ({5{1'b0}}       ),
  .kh00jq7wde_slaj       (fyeewgjh0ejxrrn), 
  .rezwnhzl7vmkg       (zpg071p8a094ze4), 
  .nq_d1dxi6n86s        (odgaqp3aclcfht_i7t), 
  .z8xxe17sssy8tr8q219     (pc67uztpd_zg6bsal),
  .mn8sk0gr9oh54zn_o   (pl1e1zu0kmorvnh8dd1yd_7mi  ),
  .oetzq1g528ymdza0maph   (uh0wfy2udciats10exk7gx  ),
  .x11xtpe4e78unv1ahgzinz4n (q3ob282pxl36b1j5u1cpl5ets3r),
  .ialrcyi5grz5o0hc0jyjuwv (yrg9fg2dzj0h1004qftims1),
  .bwsazwvhtn9in7lpyjssdk    (imk1vol1t7hn6gevzps7ze  ),
  .wfpum3du8gc8hr_xuerx  (voug2bdbrmjvpkny8ect9r),
  .aly0oms0x8r1kmmdgyob   (da476r5mk9l38ofvakaxk118t7),
  .vckb4tc8r10z7n621obxkju   (n1vkvib_j_0t8v7t7pjy3uio26),
  .f3lw5s13_0u5q6o4ep   (r01knk1me0t4m3ue2ok4t6m),

  .u4k7uyzg9lp3zlf       (1'b0  ),
  .cvqaktep17ac      (er1ax0dpgq0b7g6i ),
  .h91pmjbyad1itr37      (lhs982qsuxsw7i76wzs9 ),
  .mtsy6_whdwum2fu      (f09gaw2v2ppnj18jqy1n_), 
  .k_igx5_oeq1ag3m      (o60e9qmmyfyb4lr     ),
  .th3snuy_v19o06eanj  (ymf9djwm1ss4fvtr68bfi ),
  .xxggjmznfu9b_       (erx90sfzu891aujxq   ),
  .t9kvx890cyg        (qtfwu64s5lqiyyqles     ),
  .i984chc2gxtcivks    (y4so7d4uu1lfqzpbgq ),
  .cyudxl51e         (cvvsn7xc8qg5uk        ),      
  .nv33gk9s6_         (xnf360j941m2n        ),   
  .w37tf6nz0oty_z89xv1    (kmw5zvgvlfxa11v33),
  .pfeci7n4c83yiwln58    (sb8c9xuda2cis65y1ho),
  .mzu7xfmjf4mwa0b     (llejtcklcswz9nau7td0r ),
  .g3t8ql0mi58ddizau_8t3 (og_162hdl7wzfuaufz03z),
  .gg468ty1pm6_zgec     (oy6he9jrp6z3la4aonl ),
  .jtvucg9wp5nxn     (w6j6nqqawzzgqlkzfpnm3 ),
  .ofe8xctslv6q5w48ky   (e8ek1pn7po43ud9g42t),
  .tv7ak8mtfqswt      (x967n2unm25k5336wf2),
  .axbsuznhe7w6rrd      (x2uw3xkpg8k47k8i),
  .j49by1lxo4ie9_ho      (po0i9bzsw2yj9tv),
  .rtjejhmafpq7db     (zhfhfu89sj5v_ci5gp96ysg ),
  .vnc88f08k1s0obtnvb     (zv7y8twrabykb59a8a4629),
  .u5pfnkzvz6fsvmgw4     (p1xbmu6wvqhuu3rp2xt    ),
  .zlk2yur1jgjwg     (aq9__1ut60olwyc0dv_x    ),
  .ow91ik9ily4bugcc43pp(e0xd37xbhk4bxmxa9_93qr),
  .bf8iyrsqp4a2s           (vynn8pxcf1uhro7e              ),
  .pu764metopn524rq4hg2c24   (p6pm4fdt9wqk___preo3g4ppz      ),
  .j7l4qmkctu4k_1q6c         (ynb8hbtopto1okekngx8            ),
  .x6t2ufv1z2uufogo         (gc_pvwtyrxrfkd4sh3xn            ),
  .q5_q35rctah_              (sfrkf5j74_e8qi                 ),                    
  .hm3iwty3s1d4si2p4           (qryqhxq_uj5viaeq_tql              ),                    
  .txcys7e9ezk6xikpy2hu987  (no7xdtjyy1_rzn5              ),                    
  .eph11j28sez0oftr7b         (iecuqnis03sogixkg5at529            ), 
  .lq6932o27hlk9v4f1m          (w9gp9paa_nei_cgq5             ), 
  .sll07sleuwo2fkitj       (vtx1v5trwp6v5uo05kirprri          ), 
  .v2e4q5r07qxd6fxruqia3f       (nvvhnw32pu5ftxhzv6ycffp          ), 
  .e5nqx8gg2u3gxy0y4c       (kfooiskivym4ubj3utuxjy451          ), 
  .ajka24wmafrwpta96cf2        (j09fc8frtaff7iig7zoft           ), 
  .bod813pzaejozw9p1         (ihlsip_az_gbdtb7cn43tr8wy           ), 
  .z1et08p41uxcl76          (pt8li1mpvd04qujh4o  ),
  .jymdjzitd0hv0e9uhul        (kgd8co1m3ta9_sciodf),
  .juyjh9cdf4vvzhq   (gyxiq3yqdnanuqt16bh7r0h),
  .pwppbjb8emt8vd9_w        (l_h0z16ew816k0kc59fz),
  .z69pfny03ofcxvjyygmo6      (v1_i1c87etnhn8gl6t64rr),
  .vh0cb71_xnjsewqur3 (w0p_8cae4cqs_1hdeoydtp),
  .gbgabhg8e_ul0e24r6jq (hncm6yp50zjrhz9dcp1t1q),

  .lot9xvzuqrd5jm0scdx5t       (q7iyngsmbckvi2tht2wb5nh),
  .mn3tic51ckga0gc           (mq09q0m1l74z182ajkt2udd    ),
  .k0be3wres3xocvs9tpkn4fu      (xsziw9gaor0xrlm1hvlpjr),  
  .akk0_n8kvb1w0wxrz            (reu5ooijp0czeggc974     ),
  .s6in6vliinq9udhsofa         (b81kg80kxviv6w2l2dt8qq     ),
  .cuxay1hemfm214cwu1513x         (b6p6azv95fkv2o7od5rkww9t  ),
  .ephp7dpea6ymyg0eucjv0        (m5mjr032v1z_erq3mxi07t3v ),
  .w42z5c2wv916u4df79p            (kccav9va65o92d7d9d),
  .ej5tfrzf8ad7noezo8gdkb1xg4   (qwcb6hcmvfqmf032z        ), 
  .ekmvur7r4qz7ea7htd             (alu_cmt_wfi             ),
  .ndvqmbwgzq08mbdaxnn4          (abn9qjx8er38bt0stedss),
  .rx4zxlit4v_5k4fclu        (phiz5ah_lfipt6fb6lfzws       ),
  .vq3a19my9wldb5hug_nnbu0    (eih6zsu_r0tzn0s9udfs5ie1mxg   ),
  .imj0glh0tzynz             (tb198r6lzk1sr77g4             ),
  .k_7iagb48feg9b3wj         (kzmdmorjvnpxc87jh5yawhk),
  .cnp1c4afdljmpemgot3sa     (ga193bfpsqosp5on_bftetcu19),
  .wsh7h1p7b0zifvs0kwabih        (dibc8pgq7tvu40lvceswojwq),
  .qhk0gez3kmex8twzly7mxn         (rqprsakhpq9fka9os5knx7kiw),
  .rafwujb8lw59lcbn9vsz8o        (vmspdud3fb2xydastwgm95),
  .dqpwtmmizdh6bvzsx6          (bzjveslpnkrl4_vnqp01r2),



  .rgip60bn9st8htirgmhnohyj     (i3fga9mifalr9g_siehz7127f4  ),
  .duo6acmepph_0ahl_0ebyyjh   (sd8rqg0mey7v6mthfjratzooccvk9),
  .mylxtynzir7dvcouvb5thi  (e0srj1jifo6i8ocnkw8xqhp  )  ,
  .o5yttui8un64i2r3s3yxxxjc25iwv(ckrr5bi6ad3t5_60gouyjr9vvpfr)  ,

  .fxsynukaasxx8lt57bwdodyn3cem (flv4ybjx_fxnt8ahli      ),
  .oel93f4rkl6esczbag9yld      (mp50sb0x32pr82qg           ),
  .vmp6zvyj46lrfmg3bl_kecu59   (r1mbz1476mmd6eb_2gb        ),
  .gj_lc7e2uh1cdx5b2bmynhvw  (omlfl4p9_5zoeeas3       ),
  .b7ker79ak62g5qei_oa7kxdm0  (p0e6oiwfprzmn8yx9hsoby9       ),
  .i3rcr_tmnynzs9lr254bac9x2b (ue5tzeds4j8o5wx5zkx      ),
  .ti5a3yv8_m3rzzigzeuzrt1 (hraqlcavq96j53yrbyif      ),
  .cb86_62ddnv8i2whbc   (bf5ypgqi4grkg506x        ),

  .i_2lk2qupeba0sjgw6sdnbedc      (gkjb6c98b5j1zsgbv26  ),
  .a46z1a4rlrucmwj5ju3o83orp8jx2e   (unntlrmfpzgdq8rnz3ug3_8  ),
  .p8zi9oi86dxmkaq4uqhu8j1hl0e  (asxvrob6s2_85u99em22  ),
  .plmzz80_s0_tb0kwjjgu5p7uktpi2  (bva3_s2oj2hgomj0eyrk  ),
  .ti9h9knu4vrm6k3vqry9vfxbc4b  (n9q1kib2q28tfyzyue2j2or  ),
  .z_r1pp7wjooqw6n7rnoyv7nka81o (fbgda1d6z8gr725snyc2ylc),



  .kr13pzf9ml9ic_vbl            (1'b0      ),
  .wkixlev_tj12x_lfp6p04t      (hnq2agjqmp3jnfvc02q9vn      ),
  .jzx45r8bb79aj5ddz7h_565f     (b04f0gnze13bj90dolndjwsij1e     ),



  .pysgbgu5mzucuewf1                (abn9qjx8er38bt0stedss         ),
  .h_4gbwx46f8brur_wc           (eemxwz9vo25r4djt76yzhab1ue     ),
  .r26sxdceh7f2t6xroiyejiud7e       (gsmurqtk28c99urfc3mhf1804),
  .nabilb10azux1hnithsys          (elfo368_wilpagxfb_udyc10aej),
  .pcmvrs0wuwr_x06ql              (h33etngddojmz59z88a1yv3    ),
  .du9lzthd93rvmfcw7rz0wap         (qbwq6loiooi7x8oz3mm),  
  .q2vmic6hc_08xqnvwhw               (qcs_9_0j844qh49kucr_8     ),
  .v175vi3kjhjhl37_p            (blw41o7zqxmgmztc9cwl593q4  ),
  .vir1r5sxmryfghdpp_u82bq6        (y6zepdb9e4svr2kxsxig3dej9  ),
  .fqx1jny69kgy_gimut           (vmcutkgts6eafpyi257frl0pq ),
  .soumhrmo71_bkr9v6s5            (jxknblho9wokk6irza7q48k6h     ),
  .sd2su0k2v13e1jhtkwj               (nmn1jadde_4_xom6aqb),
  .ruzuip2lmd_5bjdch            (oungyftsa5o1qeiq0zbvzw5f),
  .t7xboey2yuqaq15sxya1b5           (xckbb1f5bxl8d6iqjh7et8uce),
  .v4icsnfwb3y76_4utq            (b39373uuxt1fwwvp8c2yhm),
  .u4560ic2z4t9ft8jb0rvw           (qm7esy9r83ecuoam3onh6tm),
  .de7s4aih29brxnb18p             (dclg9gzyeu9de8scca2r66),

  .dckyl_qt92wqvghtw3              (v_t46_oqiae0c4es9uht        ),
  .vyug4w9rb9kj6bmwwu              (xw9obr7t22kfov7grph7        ),

  .v8zi5h4rj36jt              (),
  .livvja2ywo91o8v              (),
  .t5p9q190fm              (),
  .jdngc81st67hk8p            (apf9b6zz11802cqi      ),
  .u4t194j1c9najq            (trff4kgfudc86mj      ),
  .ptu54kun7juh0           (qx67s81zzlmp_0y3     ),
  .tsns5phts_z2fnf           (hmu_zk66odn2umlzrf0     ),
  .rsdyvyptjiksvewu           (z9601_tn67y_68ndtufn9     ),
  .gkzjw6iff1idxo            (ooadt7528tbax93myw      ),
  .jcj76rmi3pqujm3v           (                    ),

  .fw_dplmj46w6              (em0guzjh3x0tokxd        ),
  .akdv8vv97zk549v            (i7qg9zxylz7rpfw286      ),   
  .k_wnu24cz94zwh8            (aykpj7s87z_wdrbcx0hx      ),   
  .g65q46nnz7gip0zyo          (tcveomov4rt0zai5ns    ),   
  .zf1w750jg2mtdij           (ztrmt5hqf4t_572v6d0p      ),   
  .pw6i533r0oou6ub            (r1upbgyfw2ogtmd_      ),   
  .getq71b86zu18ri7x        (c_2htc3ogchp6l1b_ocaywwd  ),   
  .iouqv7uynzgvde_v             (vztmqpg2g1jegcsjy             ),    
  .hb36pq8e0n24raht15       (lvi1vea5zurx7sli3iif74       ),  
  .xphk4z06widyipxfcjr       (tbuth82v2mm2g7uok_hiph       ),  
  .j9fcegru44_r74xlm2sbp     (anj5c56sztftipab3_sfkos7yi     ),  
  .uw1jajj_fvu9278tlptmv_     (l0z8mly9ui8x1u5ulfb4walt6     ),  
  .xcu8n5tos13pfc6jhw22       (),  
  .tdwhghf609ku2jek72pn3     (),  
  .lbx9pnfl2z4is68kam      (),
  .hl9x8gmcd9k2ttm0hui2j      (),
  .ioka849821_gx48yl9gk      (),
  .cc7_9__0hrnupts              (mq4z316n9yhcwtvfe        ),     
  .pba2_zyealgm_jf64t          (hiqrrqluaq93akcapxdylg    ), 
  .zpdph1sve               (j3zy8mipfns_ki             ),      
  .o9d_zhwhmsph               (xls7sq397kcp2             ),      
  .dte0cay394mhjhkr         (hno6u0yd_gjy_1t     ),
  .vyis_kjmkr7org4mer          (o88kin60h043_xvw1jjqkq ),
  .n20czkexgpbptzj5w          (mg3fx2urlykksnscs_7t0 ),
  .uvysjueb4qilrx7           (clqozm1jbmldowubnqirw  ),
  .qd0yrkr028oru_36lsp9       (yhtdgk1ljckfa3gybu4ofkrm9 ),
  .zkhg8302rekq3           (ysh2g3tr4jy_ogbn47v1  ),
  .yjox8n6veh2dfp4           (kf_d85407aznl0ii  ),
  .xa_tll8bjyk6hu8         (dm23tkdzwq_nstqh7q),
  .cmbn4qx1zcverw            (mqkvwvl8pflc9cluk),
  .r9098zakm9jc            (seo11tmtq27hed2p),
  .ye_x11o9y0je9god            (mtuge6clzfy0w9er3),
  .tp46wehs200pll2qi           (),
  .fwpoqfymdxr45bq2   (pa6s_tjxpy4gq16f7iur7   ),
  .rnub9co3myzraj2l     (o_adoo65svxjvftm_rm3     ),
  .azbeqtr4zo_xorty8     (ix1bi23f1mg6sekjqzl     ),
  .fv_51fuukywshp7hm     (jwsf_7nftft_w24ca     ),
  .w20nxrvpdf716_     (evh7l6yf2zeh1opg8dw     ),
  .x2ypwv3n6g8jsweuweebmhq(gsbir68u7ok8gu2xesw0zek ),
  .dwvp6uc1acommla           (lbuuy3oqfy7m98dnu6x6              ),
  .p8to9sivjjwpc0pn2bvf21se3   (k48o66po4ld1pl217myx5me3      ),
  .x9t5ge71i97il9r8         (ai272s0_wt92lhlok1_j2            ),
  .n7fla3l_dqx9jnxul4         (rj9754hija256ughfk96zd            ),
  .h40f1u8xaz57o3c          (mhwy3r0_oj3dwbbkxci),
  .bv8rdomgcr9w6r2z          (ktexyfhmd3f6j0oghmg),
  .ujgn98iv8k5xidjk          (imkdfcjp0n3752tqx),

  .vg7c1san7ef_              (sdil6s1uzxtjt_viwt                 ),                    
  .umwzm3ilav51kmk7r           (ik7kganikfrfc8z_c              ),                    
  .c8l2f5n1fhxm76kt3vlu6jp  (v9o_kfa70i0fkql780cet087h389      ),                    
  .hibevegtudxlh_nk6e8e         (zscjnjl4ffiey84zel2            ), 
  .y6lolb8cmealsn6ev          (qy0ycb_z4ngy2ll8pqo             ), 
  .x2bck2rbbpoyqbz62ld0tg       (nlptjpg_zybrljgsnky1iwvhf          ), 
  .abkeecplc6ueo97vo24tg       (zgv8w7jqb5wr6l2elow5znmm          ), 
  .b_fk_j1filrux_uod       (rpceina94e3bcz2ov7g1t_iom          ), 
  .oaedrllyjbu5y92f        (z492i2r2osjb1wm_z8kg_vzs           ), 
  .plgwduxqtms73miw0         (svrztr5zqc119uyafi4qw0w8e     ),
  .mf_okovo5c__xpv1x          (vlpn6saddwb42teg),
  .i1_2srs1sequ9t          (m3kk01rml527m1oq0v),
  .a4aa8t_dofc7_82w          (d0g9hx2h2bufn9qst9s),

  .q6sud8b_vapga5ru5c           (c4i0yanuek7va0ztp  ),                    
  .latkf6ie2l8fv5dg98qec         (n5x33q1l9ewebt6692qaofd8), 
  .azmawprujj_u7q6ofj          (eqhoch739wo4sqhno2u),
  .wigxwsu_39gcyutr_re          (qj1fn7kk041c_7kez4t2fkt),
  .l0_j3191k35720flisiv          (q2qa0la3s98x10a2aqsb73g),
  .cf059q4pm79who8jb          (ajk1fk4kecwsdaeiybv),

  .pket_pq2m99ayix3fk5yps (g7rjoc9tw3_k7r1i21ghnsfcv ),
  .ty49bqt9pydf4fr50f89 (g_wqbz93wfi5bmx7bczdub7 ),
  .itofghyluwwiwmqnj_4imeao     (tpd5fcgyg_240nz8md69oj  ),
  .j47kiegbvv22z361yv9n5   (npkoy9e2dsczayfq7h6cko59),
  .r75dlj23fr96kve4fzd8xpw2zn  (kmlf0ops49wvgcz2howfob59khsqir  ), 
  .mx7juirxj661i6i9lns4hnnyw0ep(kw590mop2ic8u619z7c_owrnv9t),


  .frehkmd0xqj4qeyqqodmp0onx7 (oa_1ibjpvwpv6bg5ivcau2uo6z3s),
  .ms95k2pmbvtrb33p5oa2q      (noc4nf4qform41kyqw6m4     ),
  .r928tvy6d88uh6s9qun65udol2   (ktqyocabrct3iqhlj18u9fhnz6f3d  ),
  .jtgchf8072p4v1h9xclp0t  (ihbxqlci_5lmn6uyuoxv158n18bua ),
  .jekm9yqqqogc7_czwax0r6an_f  (xv9g6nf92837e31mav06v03y2t ),
  .vs9f2qtmvyxt6ycc5e_z47fnjr (ppwfzi9r2pfdu5oiww3x5a9g94u6ut0),

  .wvywyxp28r9wdwncg13zbc_6(by0pbwftr5xjmht8u5rapxeyd1g),
  .suaktr_howpmkqxx3p5j4  (z3m510kw9uow1_jbl0xi6lrg   ),

  .mnym6ha4fxtg2oqq9hlac5s1      (leq1ne49igptrh__p_5kz23048rjzm    ),
  .p6wfurur4eut85r8tktdi03zxb   (ipj0pyjf76qkv519em1jiaiutbhsr ),
  .u78ade2idh660umk_1m66fdlksb9b  (szaorjzmus1ssgjq7e30bdssuadwt0),
  .xxr9qx83ggzl9q98ig_ys5w60a  (yi0r5xirgktqhr99j3jz345g11t51),
  .lozr9fiy6p7y8rinc582m2bt2ha_xmf  (ogkluwmj9mmpgtmicjnh6_yya46ukkp2s),
  .z3j5lbdgqwmp5zmv4g_zn29fgvintdc (d250junaig195xflrdmkjjl5pxtaf4 ),

  .ussyj508sxu9v0           (h_iyw8puc0v6p12hca799v99  ),
  .pdns51exd9ffhf5pykv42sq     (ak3_rgqx75eo7s2jfbhemwqz8ng ),  
  .k09nslb_nkoy4r0t34xu6    (hbinkk7e8nmokz2d2dm9gq2j82r),
  .crr9jljkvi3gsixv1_v8       (d228vs4sizjmlag0hkfk ),
  .sca7p0942a6kocjqqvat       (wz4he34y3_e1ieaudx5sv ),
  .go_m73qp_w0p7abohs24       (r2mcos1t0vvp47i3ka_vsc_ ),
  .jm4ru1fdiqtw706w8        (woqfe5v065k3eom51g4h1jq  ),
  .j021ufdslrlb4m5c5h2      (x6s44jsh488qbnj6v9ppkpceb),



  .p1kjflyurzeuxj (),
  .yvjlu1e9eng5_5tme (),
  .hh8nc68zrpki2m9r (),
  .v8wv99vga5gkl8xhk7x9in (),
  .ahfx5rs9jkdyw3b8ztscfx (),
  .ts3_k4ergzh8upz7 (),
  .ktqya1x1mfi5j3q7 (),
  .z6njhanl_m_hv48x5i9y (),
  .dvm_h24fnflt11prmyvme (),
  .uvyubcp0tbk9yirhz (),
  .ivoui15mvw3de5ds44 (),


  .gf33atgy          (gf33atgy),
  .ru_wi        (ru_wi)
  ); 





  wire                       qwcdw99v1uotvc5emiry7z  ; 
  wire                       p1k8b_ul5r4iaqvma4l ;
  wire                       ctgxr_wil90tj1ur64;
  wire                       gqxkhqynd510udp0tpbr   ;
  wire                       u_hs70f19eo9kuxrncia;
  wire [64-1:0]   sp1w3gxueck6hge7wiki;
  wire                       akig71_dnhvxrc3d3u_de;
  wire                       w9z2kr44j8w6w3w1zqa;
  wire [64-1:0]   q94xtoze0utbz_anbev; 
  wire                       e43glfkwrdo0_s; 

  wire                       gbzetyyhf8hyf9t; 
  assign gbzetyyhf8hyf9t          = jwsf_7nftft_w24ca && pa6s_tjxpy4gq16f7iur7[9:9];
  assign hwpkcsh2atrq            = hxrmt706n071lic0f7 ^ gbzetyyhf8hyf9t;
  wire   ppz7pt801h8fopmz2r6        = i7qg9zxylz7rpfw286 & aykpj7s87z_wdrbcx0hx; 
  wire   yt8ni4mv3z6738d0cjg       = g_wqbz93wfi5bmx7bczdub7 ? qwcdw99v1uotvc5emiry7z : ak3_rgqx75eo7s2jfbhemwqz8ng;
  assign v3e6l1k7eo9k3           = yt8ni4mv3z6738d0cjg & ppz7pt801h8fopmz2r6;
  wire   l7syduiu9_pn9k_8llfwh      = g_wqbz93wfi5bmx7bczdub7 ? p1k8b_ul5r4iaqvma4l : hbinkk7e8nmokz2d2dm9gq2j82r;
  assign hxrmt706n071lic0f7          = l7syduiu9_pn9k_8llfwh & ppz7pt801h8fopmz2r6;
  wire   xk32a7aw5px7i4ned2         =  g_wqbz93wfi5bmx7bczdub7 ? ctgxr_wil90tj1ur64 : blw41o7zqxmgmztc9cwl593q4;
  assign texy7g6tpvcgwtyd           = xk32a7aw5px7i4ned2 & ppz7pt801h8fopmz2r6;
  wire   zmkqqbcgacufp_na86275hfye = g_wqbz93wfi5bmx7bczdub7 ? u_hs70f19eo9kuxrncia : y6zepdb9e4svr2kxsxig3dej9;
  assign gfod0nmy6eta29jeeg6mr2     = zmkqqbcgacufp_na86275hfye & ppz7pt801h8fopmz2r6;
  wire   pls1_s6_92julifn5xbq    = g_wqbz93wfi5bmx7bczdub7 ? gqxkhqynd510udp0tpbr : jxknblho9wokk6irza7q48k6h;
  assign n4soswat5yihd74b        = pls1_s6_92julifn5xbq & ppz7pt801h8fopmz2r6;
  assign if0fog4bug_zkykpi         = g_wqbz93wfi5bmx7bczdub7 ? sp1w3gxueck6hge7wiki : oungyftsa5o1qeiq0zbvzw5f;
  wire   rppmitoogp3uvxw2trfk    = g_wqbz93wfi5bmx7bczdub7 ? akig71_dnhvxrc3d3u_de : xckbb1f5bxl8d6iqjh7et8uce;
  assign a3xib90kwk4_hm1        = rppmitoogp3uvxw2trfk & ppz7pt801h8fopmz2r6;
  wire   nb8cugitmn43ebp7pirfn14     = g_wqbz93wfi5bmx7bczdub7 ? w9z2kr44j8w6w3w1zqa : b39373uuxt1fwwvp8c2yhm;
  assign nfzexr8q9g893gi         = nb8cugitmn43ebp7pirfn14 & ppz7pt801h8fopmz2r6;
  assign opkkwp3eg8g3448t        = g_wqbz93wfi5bmx7bczdub7 ? q94xtoze0utbz_anbev : qm7esy9r83ecuoam3onh6tm;
  assign tv3_4qrynvnaoy4riz          = g_wqbz93wfi5bmx7bczdub7 ? e43glfkwrdo0_s : dclg9gzyeu9de8scca2r66;

  assign w7uciar2_6p9xc5mc = elfo368_wilpagxfb_udyc10aej;
  assign ex6ixmgf331     = h33etngddojmz59z88a1yv3;
  assign vfu1cc_k9n55lt38g_vii =  qbwq6loiooi7x8oz3mm;   
  assign gkps1gyqdwgzcvr0c  = vmcutkgts6eafpyi257frl0pq;
  assign q52oeddgdt76b      = nmn1jadde_4_xom6aqb;



  wire kbyvllfhv4g65k60,baeb5atyeipjmjtwdx66m;
  wire [4-1:0] kud4a7p3c8pym85u6, w6xoq8do9qo8kitx8e;



  wire ihuhf6fv7o59qgws8zewd;

  assign ya8t4ev_aidf0t0x4or = v9o_kfa70i0fkql780cet087h389 | ihuhf6fv7o59qgws8zewd;

  wire mkdazd4f_aukad6x = z492i2r2osjb1wm_z8kg_vzs & ztrmt5hqf4t_572v6d0p;




  m0m7t4t8fpmv   #(
    .hcl69mdlw0ykna4ue4_t1(0) 
  ) wlpgzbimzzjy6k_xw3vv(

      .w2h8uh3l463qbgqmv(umnrzb6pv8dzc),
      .tywculgjyor8ndw        (tywculgjyor8ndw   ),

      .pw3qcykea5ib_ieka(by0pbwftr5xjmht8u5rapxeyd1g),
      .g6xvfy8tj0zmajl  (z3m510kw9uow1_jbl0xi6lrg  ),

      .rvr30vvllni (rvr30vvllni),
      .z1cj655u31 (z1cj655u31),
      .lhu2z948o3n (lhu2z948o3n),










    .r0s7d8cr68i2qs1z     (r0s7d8cr68i2qs1z),
    .kakelc68be0x7tdm9b9o    (kakelc68be0x7tdm9b9o),
    .j3j1czgoam48vhs8auo    (j3j1czgoam48vhs8auo),
    .gm1r5itc44uxw_y0_msk    (gm1r5itc44uxw_y0_msk),
    .af5qc04tmn51e4u2h1z    (af5qc04tmn51e4u2h1z),
    .qwcb6hcmvfqmf032z    (1'b0),

    .veibgbyke             (1'b0                ),
    .jjzotrbn             (i7qg9zxylz7rpfw286),
    .hw1_k1jmu             (f1k1tltm39p_5uxhp5l80q4),
    .qbpmsk2              (hno6u0yd_gjy_1t    ),
    .tc88s6cm5b           (v_t46_oqiae0c4es9uht ), 
    .c3sszdooylrw           (xw9obr7t22kfov7grph7 ),
    .qpyjufa5h7y           (mhwy3r0_oj3dwbbkxci    ),
    .hvv94pmafz           (ktexyfhmd3f6j0oghmg    ),
    .e19iv2rqeu5          (ai272s0_wt92lhlok1_j2),
    .m4y6v4ncsg          (rj9754hija256ughfk96zd),
    .le3dqob2            (lbuuy3oqfy7m98dnu6x6),
    .j_rvclhfbeig5cqeb3_   (k48o66po4ld1pl217myx5me3),
    .cpt0qfwiz            (5'h0),
      .sjunepbdn               (imkdfcjp0n3752tqx    ),
    .i7vhyhns            (g7rjoc9tw3_k7r1i21ghnsfcv), 
    .lu44s70ub62            (g_wqbz93wfi5bmx7bczdub7), 
    .yocn4o2zav           (em0guzjh3x0tokxd ),
    .ojbpo5z6urt             (ztrmt5hqf4t_572v6d0p     ),

    .t9b41sw5vpr            (o_adoo65svxjvftm_rm3    ),
    .hy14_6z7grvldvw          (pa6s_tjxpy4gq16f7iur7  ),
    .nrebzehsuam              (vztmqpg2g1jegcsjy      ),
    .b_sdf8               (mq4z316n9yhcwtvfe       ),




    .cj2osby26qlape              (c4i0yanuek7va0ztp), 
    .zawjtr32pktig               (ik7kganikfrfc8z_c), 
    .vc529nuu                (phk590vi2   ),
    .xh52jycxcjs            (mkdazd4f_aukad6x),
    .rnx27onf2lbe             (rnx27onf2lbe), 
    .aziir_r1p              ({64{1'b0}} ),        
    .ya8t4ev_aidf0t0x4or       (ihuhf6fv7o59qgws8zewd               ),
    .scadliwzjp0l78srd9p     (svrztr5zqc119uyafi4qw0w8e),
    
    .l6s_gf8go82fwn             (vlpn6saddwb42teg),
    .afifdv1w9             (m3kk01rml527m1oq0v),
    .u2bhabgcppcy             (d0g9hx2h2bufn9qst9s),



    .fhhe7189lmum             (5'h0          ), 



    .bfo1il0du_  (ix1bi23f1mg6sekjqzl ),
    .gnb98c7tbqat  (jwsf_7nftft_w24ca ),
    .w4kjodkdva03q  (evh7l6yf2zeh1opg8dw ),

    .bvzc7t76o17 (hiqrrqluaq93akcapxdylg         ),
    .begxws3d6mwhnm        (d228vs4sizjmlag0hkfk ),
    .z1nw2lilgog_        (wz4he34y3_e1ieaudx5sv ),
    .x6ywulzbb7jp        (r2mcos1t0vvp47i3ka_vsc_ ),
    .b9mfhl8am_whqquz         (woqfe5v065k3eom51g4h1jq  ),
    .bqen_oh1ujvq9lj4       (x6s44jsh488qbnj6v9ppkpceb),

    .bwjyqadn                (j3zy8mipfns_ki    ),
    .k0xug5g             (xls7sq397kcp2    ),
    .ipht6ss_sh6h            (abn9qjx8er38bt0stedss),


    .binjv97px9r7dt04h0       (eemxwz9vo25r4djt76yzhab1ue),
    .ajl4tppx98ihuirj_mxih   (gsmurqtk28c99urfc3mhf1804),
    .o_d157fc5_l           (qcs_9_0j844qh49kucr_8),

    .n1rp2mggtiknd88         (32'b0),

    .b7ilo27jne5k           (o88kin60h043_xvw1jjqkq),
    .piwiqvrjoq           (mg3fx2urlykksnscs_7t0),
    .al4xeg8mukgfg            (clqozm1jbmldowubnqirw),
    .ryc6z1c7rmzrnlno        (yhtdgk1ljckfa3gybu4ofkrm9),
    .rhufxsnopy0n            (ysh2g3tr4jy_ogbn47v1),
    .wbhvg_1r9435            (kf_d85407aznl0ii),
    .s1woka0byzgo          (dm23tkdzwq_nstqh7q),
    .q8977k41y4             (r1upbgyfw2ogtmd_    ),
    .ciiwo7qhifea         (c_2htc3ogchp6l1b_ocaywwd),

    .u2k4dyp52s_m             (seo11tmtq27hed2p),
    .djvj1e_             (mtuge6clzfy0w9er3),
    .bktu0z1mk56             (mqkvwvl8pflc9cluk),
    .l6z1pzhjg5az            (1'b0),
    .phofig8d5zd_8v9g8       (),
    .js0ml55dtie8qenb4eoj2 (),
    .p343qo1j             (),
    .h8m3g7a             (),
    .r9ix0zzks6zej       (),
    .l8xeqkc               (),

    .v35y3qnk7mx3l1695     (1'b0   ),


    .gqe6zqljzhgt5wz98      (                    ),
    .tisftwun8guh8lnibary2gz (                    ),
    .wdgj6jexv3_u8sb4gnsv5 (                    ),
    .c_qlgbc7oqwu9as946yqls (                    ),
    .nc5hf3a4mwl257q       (                    ),
    .cqq719hbl6kax00mwmrhj   (                    ),
    .a_x852mvzp7z5occs1   (                    ),





















    .v3e6l1k7eo9k3 (qwcdw99v1uotvc5emiry7z  ) ,
    .hxrmt706n071lic0f7(p1k8b_ul5r4iaqvma4l ) ,
    .lrhkvgg4x13sq245     (ap889z2q8jbzn4dhurkzl  ),
    .y45254ns5fjfjnwjiwr1_quk(sp1w3gxueck6hge7wiki  ),
    .sshjsyphxbyaqk3kr    (rnodgdrxyr_tulm0nnnign),
    .zu8yygom_ioh         (j39tby_g7kqga33w_m      ),
    .od8eje0yjk8         (t0o4cn_ndv2lmnp      ),
    .l_km9bow2ubqs5dtd        (aa5a1tnclwe351p5ujs     ),
    .cv8rkirz            (my5_v4hhb7oc51         ),
    .mbnh9clp6pd3t         (lmv45fhtl015bg      ),
    .z091v3i7q4_rty4       (yd4wqg2e0i386ccq6y9    ),
    .tsml_wqqwnty         (uv_3uzx5ti04u5nd      ),
    .pdz01l48nt          (y_gvnr7uidhcof1       ),
    .l5zrepfg8it           (zh_0_4wrffapmbs        ),
    .aq4b6s94dp0f          (nrze6rcjz4m65z        ),
    .dmg1a5xdc9           (cjxy_cr6jzz17mr8         ),
    .v1j50zesdgxioc           (g0ovdu1w9dcoqg         ),
    .tkhm63y407b          (uxdt29u4dd96ukc        ),
    .qhkm8drwygkskh_          (cmv9vkluc86swnlc        ),
    .nh1gz4628x89          (r_cdggxn_7syt0g        ),
    .l4anyablbw3gt          (uvw8h6lqr2ou0        ),
    .vn5b662w76_a3npe         (rwip45nhuhbz2jkd4      ),
    .wigtf10_bybfdpp_x        (x3r6u6q7ck5ud8wbii     ),
    .w2gbqib7zable3o        (p0ga7mahvd8zjma     ),
    .zp24wdce6ufxkpbs        (hlxcm16byj04fp0     ),
    .xxee65tc1tureck      (o4lqcf45nah3boccbw   ),
    .wr1tfb0_sg9           (alu_cmt_wfi        ),
    .enhpakthwj3e65vldt   (alu_cmt_ifu_misalgn),
    .mz47ksy6nekv1cbaq75    (qjg3a6detqucp4byrgs ),
    .egplp36i1ttcggdv2b0xo2e(qn6g68ul7q8pz3pvopdmh0m),
    .rbsutocgtudusq3v    (kxmzp6o3alj05dfq9d_e8ci ),
    .sgy1x259o9ltvsfe    (d2gcdo57ra3yxudimcwal0 ),
    .tr2dgjt2yqfzjaos9o  (ob__kc7kdtjxp74ajo7ql548o),
    .o8m475rdcb4y71zte3fbd30(co8g52huetu0l9justjw5wcy19yi ),
    .nzm80hh72kwblbx4fcg   (ihmezohdr7mg9_blli7  ),
    .l9wonwtwviy4i8w6s     (                    ), 
    .wuw4k4dyuslqkjap     (                    ), 
    .s4o6xx8w0dylrebxlqmia79t5 (                    ), 
    .br6lhce3u3l01blvxzrqphj5svlum(oozkxp7aywu4l0hz73uedbtyiad ),
    .isvwkofue95j9ud7p3nrgntc(),
    .mf10lk374lxu341vp3kpfl6 (),
    .nkemiexuw_o6b34go    (),
    .bnnsit7f_1yqs20xcxk3l     (),
    .c2vqeph9snojapvdushbj    (),
    .w8wwz5822d7298zis7      (),

    .zq261z2pygzc0_h44fo     (v85ovm_7gp20oi4vj  ),
    .g_w5s5kg5qk2w1gyo7odo2nubrxo0(j5wtbhk36xx9j2h1kgsniu9p0d9xzj),
    .b1iduhkyfb7xynn3btxh6lhgev7_(qh0m9d6yrl5kb_1vvecw1kb1wrbm),
    .ndtc71v47ribx6u_eqsx8tdk0  (kihyrfzcb87yz3qnxq7c0o11at5u  ),
    .efp001u9ffq4ypu8uk4l8tbblt8  (ho49hpl6ijpiop4thzf8rh6apio4u  ),
    .fce921hmrlbrv4qdu4cb0pee  (wk2sssl74c1xyhbm7pf29qtbpws1  ),
    .twjiv2hewisn6o      (vxcgun4z0ztx7nmvm   ),
    .l4i6kd5vs494chi      (fq2y4oplmud5drf9s   ),

    .d7kpxfpyhil_2nt     (ne5matgyfjvw3elazxt7p),

    .jugi02ecegnos3        (e45zjh64jxwnli64ak ), 
    .rxjuugktc38un        (ka4_ngr35vo6rrkp72 ),
    .h8wu7unf_ixmxfeh         (jz2qz87howt08ld8lq  ),
    .b84l246u4jmnu        (jhes_c10xw065fcx ),
    .kdpgigzs75vcc1d         (dg8pvkc6n2uz2w2f  ),
    .uh251o1pav          (ngiuqj2j6rsgfaeu27   ), 
    .vjkz8n6i44pc7o          (zc9t_vib9_fw44d     ),
    .cwmxezrc3jv6hzxcfc (cwmxezrc3jv6hzxcfc),
    .uig3ujuyq0_61kqb (uig3ujuyq0_61kqb),
    .nb3w1rq_ny95rvrt  (nb3w1rq_ny95rvrt),
    .xc2becmsn4fcniw6ks   (xc2becmsn4fcniw6ks),
    .p_yx415so7q1vohijb (p_yx415so7q1vohijb),

    .suxmggt9hea4ao3r        (               ),
    .kwn45x5pjj_5mi        (               ),
    .lp9c9xlhbpjow4k        (               ),
    .ts1jnweqrdhomp        (               ),
    .ze26d9sog9r3thx     (               ),


    .rb050tnl             (rb050tnl          ),
    .e1go3iu             (e1go3iu          ),
    .el7_p8jit09           (el7_p8jit09        ),
    .a94vd35etec4           (a94vd35etec4        ),
    .l9erxxpnphqd26vg9        (l9erxxpnphqd26vg9     ),
    .guuvp01vkcryglsu1p3   (guuvp01vkcryglsu1p3),
    .hig2gwwbeuhnt65xrp       (hig2gwwbeuhnt65xrp    ),
    .vf5xcr67bqhzlo43_        (vf5xcr67bqhzlo43_     ),
    .vmx1fh4kmh4c             (vmx1fh4kmh4c          ),
    .bj7h5jqg66r51jxki6emra   (bj7h5jqg66r51jxki6emra),
    .zmfo8cca_77pc       (zmfo8cca_77pc    ),


    .v657dksgaz1cki9         (dkmuhc79d2wm0wubp  ),
    .qzz1jhwf_vd0r8g       (u2demhkod_er3kf6b),
    .dwn42a1uvd9x3myec       (uz7pt71lvqit85od),
    .uiojikf9vcnz        (v3uvhtx7e5vbtvie ),
    .x1_k6oouttg7m3f         (tmqkgmlzi018 ),
    .fcvvhg9v3mx         (lx_olubu7t8h ),
    .l_v5xmhbzqc         (dd1p3tnenmm9r ),
    .i7iq7ecm_d9pi6uw6       (l60zv02z95hlayri ),
    .p5fn_ooo9rctbxkgm_jui    (l1xzyldaa9dr2q7mla ),
    .a5z_23_ryr_m29hhia_p (a5z_23_ryr_m29hhia_p),





    .isz7jw04u7k3s7b398   (kbyvllfhv4g65k60), 
    .q4_7fnx90rztwn6_8dybi   (nvpglpdnii1iho_rjkw8),
    .zq2e9j_emlri_qjtg    (du9nxa6qo7knx2et1gw6 ),
    .gw6s_h2ymbn1ds50q8    (kud4a7p3c8pym85u6 ),
    .qv749hsiom75nyn49v     (h7szh92q4s7x6vx_  ), 
    .vo_fj58ip6ok0srq7t5   (baeb5atyeipjmjtwdx66m), 
    .qq819v1yyh8derngk15k1   (zf3zgw37xlcc2o5eprc5k),
    .o_q0qt9vjpibgshm714a    (a9rvmf7a9nbie6nd923 ),
    .iqx3cqyh7_mpvu_9om    (w6xoq8do9qo8kitx8e ),
    .melkey3fxhhc3e649p     (gzyfsm1lj5vk008  ), 

    .gf33atgy                 (gf33atgy          ),
    .ru_wi               (ru_wi        ) 
  );




  wire gccap1c6hft7o1z7esm;
  wire ar7xgugq1a_pz7b82ds;
  wire [5-1:0] vjhpkmep8g_u_cizhsw;
  wire v19st7vd9_bi485e6ak0;
  wire [4:0] zt19omidnr_zyp2gc3bywfb;



  wire pbtolkl953sk14id0iy;
  wire z2qyay491938ppnlxuc;
  wire zeseql2htbxpugyu5_j;
  wire al3t866kz4po45vfuyjy;
  wire xutsaulafh4onxtthm8n ;
  wire me7unt7fapqqhtc6epso ;
  wire[64-1:0]m2as3qe7miuhj662j1zvt;

  sdt_3ftsvyvhysb2f7uduiazuiu hjkbz6gw9d1awyb7gp1ssmb3bnrvc(


    .y40x_uwnqs6f       (s_7qgktcx5l9b  ),
    .qlykdb48c89hfbq5l3v     (eru3qosawo7xqc6t999),
    .ejlcmcywa2ghgwvj     (ybf0zo9v_845pqb_jh),
    .fk7qm80i_py_6       (swk0us69_ctq2k  ),
    .utfce4yxn08kh9t     (j29miwazgbxlk8),
    .gof9x1lyu2n5rnf     (cw3uprz8e2rwau3z7),
    .f7t_bak0dfaq3       (zcqvodebks4c  ),
    .oy1tzeyrsbr3bg7dr9u     (wsvr7r5n5ep12y),
    .rpnvo9xxx6nke515     (i6zt9kqe09i5ky),
    .v2fkznl9m7dtfymx     (bsnlk54ub6j_e7),

    .tdg7ccg5dltr5l9s   (q58rcdx67tyrer ),
    .z5s1cielsyyeza34h (c4juuyd55lxion9c ),
    .ggpqgd6b8zuelz8 (tk22_ghwl49rxxdnop ),



    .ret9emt0e4v60a6cwap10   (o4qff84vfbn      ),
    .l5447rrn286zsq9mt6k   (x74_jhmpouk      ),
    .fg4h6qs_th28xw7il0    (z5tnbveujliw633sxlb8  ),
    .q7ns1l4tc_kuf5az3u    (l8ng5e_pa1fg07__37  ),
    .h_ld26vo8tpdty     (erdoc9bbdnq8065yw   ),
    .pxbhqh6yl6hotx       (zqx1cj9lvt0e     ),
    .toib7p7z_deij2b       (zsxgccndqw2suf6     ),
    .vqldrx_4vk7av570m8fv  (y9389ymcyh2ia2082yx1_),
    .zhwwio_mprrvjud04       (uiu4_g7j41kz     ),
    .p_2daj_9kqsf0ekr101   (ro93aearv5754gz9w ),
    .djb42mrmnunfufgxzh   (rqy9v1_k_o74etonfc ),
    .dufpf9uw3i8khwmvb2h   (ytp8_jsqr2sjmu08gdn ),
    .p7ah58va5_2njbtv      (p7ah58va5_2njbtv), 
    .u981qrwkgi5h0e72b__gg19w (u981qrwkgi5h0e72b__gg19w),  
    .p0i2i3v3j1tclelx51     (p0i2i3v3j1tclelx51),

    .q89zlvtwzxkjd6h5k     (keta7gjvl7x   ), 
    .gjoru9khthrg8j6pfamu   (xg63_va9bynd285dre ), 
    .vf6etunsloifr12azv4he6   (no1k1_uyge8hlp ), 
    .f63hhh0gzajzsiyjd8cqb   (mwzhu7wrbq1rkp ),
    .v7f1q1_fp5fc8b_u     (s1j5549fqdsj5ad   ), 
    .mvneatl67xbzspkpyi1   (onnke16xcq5904dt ), 
    .ltzlg4gy4noc9555li   (msqwr_9vjwohg ), 
    .nfozodmnsmlv22fi3oe   (fy0rb852ky8dy1 ),
    .vmwegtj2c0zt7rilpw     (qgpl_3pohcjc3g   ), 
    .szgl0r6i254qax8jkjr   (w5151c0ak9j8c ), 
    .bp90ffmjkj3u4__poo   (kf18wkamz8k9bxuv2j ), 
    .nq8gzr65b3p_cdc52lshh   (u0oho0bfx9igpi ),

    .ju3gksnn2mup5h81eh28   (y7rd1k0an54clel_5q6 ), 
    .tymuflph4h7mej5umh86   (com03bquiktu249yb0 ), 
    .c5csn3nczo8zlvq621sy    (tzg0yjgx9bn98i  ),
    .g5gmidj6od8k58avl_h9y    (c2mipfm_6z5ef4p3aoz  ),
    .h5w2di84ketcahr4     (y3z8rf7c6hvsiux   ), 
    .rd0rvbiicactt4sbf   (x8_a2j7z3gz3l0tfjqp ), 

    .lanyt81iat_ws21fv   (xq0mj5mg2_512eu4 ), 
    .b1eabu9fa3jnjln5tc   (e11m1298jo38qcwq9er2 ), 
    .nt0ndhbk6x29ae8da95    (ec94_mk193di7tj  ),
    .u7vn3gjmd4owzsi7tk    (m2sw40fca0wvnmy  ),
    .ik4ulvmx89l0u0ko     (ywhfwlbfro2dmuvf   ), 
    .ri8f9g_paihffhz9_8qgu   (nodrapn01yl1vxle30p ), 
                         
    .nz5iij5cadsnx4fokudqbo   (ex_g_cnadtiu1r9u ),
    .bz1hc72g_22hgoqs8   (orzasugx5h5pio22_ ),
    .wctv6a1mmq6dtwsg9n    (dxwtzud_wfj8jqk0  ),
    .zakjetcb_4mzmn_bchz    (gi8o690aydhqi8  ),
    .ys8dsx5hx_injk9b     (zl1r9cfvuhltjq   ),
    .onijw658b2__et8fr1has   (dn074lh73rzchvrqzm8 ), 

    .o9vvv_q4ikz_2yp0w    (kbyvllfhv4g65k60), 
    .c1ilkc2r6es72c5h2vcc    (nvpglpdnii1iho_rjkw8),
    .l3sefagtx4ai4ljb     (du9nxa6qo7knx2et1gw6 ),
    .josyt39cvr3gignopao     (kud4a7p3c8pym85u6 ),
    .bjn5x3u7v4u3rm6d      (h7szh92q4s7x6vx_  ), 

    .ipq0f4_yvmml7o06891    (baeb5atyeipjmjtwdx66m), 
    .p4jgl36nmqe8ud7_g4i7    (zf3zgw37xlcc2o5eprc5k),
    .wyhg5n7dklr59dxgm_bs     (a9rvmf7a9nbie6nd923 ),
    .ubk6j4rwgfrf5ryn1ibp     (w6xoq8do9qo8kitx8e ),
    .cbr_upfu_0ywren54f      (gzyfsm1lj5vk008  ), 


    .ll0_hbknv5bc_8mxvx5c (cwmxezrc3jv6hzxcfc), 
    .qloskxsiztazdeq2ad95i (uig3ujuyq0_61kqb), 
    .px17v86p_7_1fdvm1w  (nb3w1rq_ny95rvrt), 
    .a3g162j6o30b4qdpd_z   (xc2becmsn4fcniw6ks), 
    .jb9locwfccqzb06jjon  (p_yx415so7q1vohijb), 



    .p1jdw9loxkz60taq_vkp_3   (p1jdw9loxkz60taq_vkp_3 ), 
    .ar7xgugq1a_pz7b82ds   (ar7xgugq1a_pz7b82ds ),
    .jwwku_el5h5h2lx6e0kyi    (jwwku_el5h5h2lx6e0kyi  ),
    .vjhpkmep8g_u_cizhsw   (vjhpkmep8g_u_cizhsw ),
    .v19st7vd9_bi485e6ak0   (v19st7vd9_bi485e6ak0 ),
    .zt19omidnr_zyp2gc3bywfb   (zt19omidnr_zyp2gc3bywfb ),
    .gccap1c6hft7o1z7esm     (gccap1c6hft7o1z7esm   ), 
    .eo5skx1ygvzuasbjgnyl    (eo5skx1ygvzuasbjgnyl  ), 






    .z2qyay491938ppnlxuc   (z2qyay491938ppnlxuc  ),
    .pbtolkl953sk14id0iy   (pbtolkl953sk14id0iy  ),
    .zeseql2htbxpugyu5_j      (zeseql2htbxpugyu5_j     ),
    .al3t866kz4po45vfuyjy      (al3t866kz4po45vfuyjy     ),
    .xutsaulafh4onxtthm8n  (xutsaulafh4onxtthm8n ),
    .me7unt7fapqqhtc6epso  (me7unt7fapqqhtc6epso ),
    .m2as3qe7miuhj662j1zvt (m2as3qe7miuhj662j1zvt),



    .gqat5ctwgmxi8n_5z03tivvpgqx6j5kb(m631c388smkc86tlvjo8cy0euyc), 
    .zmotzlbzlmuf2isjtqn2h8beel09 (hl8tx_5fn5baqsm5i614qe_ ),
    .vi7663z7hxlc4ngkh1_yfoxfpvbiq(gose7syxzsxbsjpxu9gf46ryn), 
    .ql2r_7apgocbap5k7ucf5a673x7v (ydctapy4pueuwk6n3mwwodl2o ),
    .bm0yhprev2rfpkaztktaxtnq7f8q0bp(xltf9w3ak66b70kftwbyhk8hfkvrk), 
    .i2kgxrwehfoyscnln10tc70_omph (v5654pk52c83hd4wif_iicjko ),


    .gkb40bm903wc32_2zjmb0l25g21p7(ua_r8723rm_0699y9ue0qself), 
    .yu_1foait_ukyv14b73xepo_1mj31mu (rlwzlq3wmb1t76we1pgot2d6_ ),
    .scom2gns1t5jrniqayb84g_h2a1zaxbv(boie2le90zg6moigey_xh5kjc6), 
    .xpvibysxiip4tytx5_ry26i78ce4j4 (jpa3mq_tg3w9jebkjw0qy4zhw ),
    .ky7mnv5l4jl0v17ox278fwktul3qti(vn7agcnzu58a7jbm9n9em4kadk_), 
    .a9_1a439ejmx35qe2g8yihj84g5 (ec2k88gmpr185bkl8ndglqu_p6l3 ),
    .rhx_hd60cwxftbqnr_uhlcmbab17eeue(yqlpqui4nfbe0t93srqmvngkzf4y1), 
    .l_w88r7i0zq6u0xtcywbwzu__s (n2nv4gollbb6vbo938tfa19gk ),

    .czyvvnzs3y3orktdmdfec8yla_1y    (kf2bfg0y804sefov7qwk95xq),
    .o_tztjh1zql5hzdma85okucmgxh     (u9jwgutri3owj857elesn ), 

    .gf33atgy                 (gf33atgy          ),
    .ru_wi               (ru_wi        ) 
  );


  wire[4:0] chezfp7x0va2ea9tdq;




  wire [4-1:0] xmi2_r3_mwq_b4a70u_m;
  wire                     u6xwpg4na3rdoy = ngy4ipxc1vxym69lu ;
  wire [4-1:0] pu89y6we99g  = xmi2_r3_mwq_b4a70u_m;

  fqo7x_ckpw9266xb2d57x8 nez96qqv3r1hdxrr37wae0y9fl_3(
    .mt0fxo7jph1jww9bml7   (),
    .katolbldvqgqsog94   (),
    .z22u8178eey1vl3   (),

    .cxkzjh6fduft16beuemi   (e45zjh64jxwnli64ak   ), 
    .uej0jzoacitho9mnzs   (ka4_ngr35vo6rrkp72   ),
    .hw1xobm2iv3kaij    (jz2qz87howt08ld8lq    ),


    .f12hi8g2fiznovp     (ngiuqj2j6rsgfaeu27     ), 
    .pupdpprs2srhv_sg    (dg8pvkc6n2uz2w2f    ),  
    .i68lo1vqlv0o48k7     (iy6jwb45n967lh       ), 
    .uwtwaa7c9764reokvm5   (z8h5zyhj54howg     ),
    .k7wz0kgj7f94f7hml   (f28m69gb9k8l_ic ), 
    .fkcyj1aq49159mfj    (1'b0   ), 

    .j26xb89a8xae2cmtqfby (p1jdw9loxkz60taq_vkp_3),  
    .mpl24r05br_tctrlxtx8d6p (ar7xgugq1a_pz7b82ds),  
    .k9ahcr_bj7e3lceyvmetj8  (jwwku_el5h5h2lx6e0kyi ),  
    .qil8zvwqkkfkcj8129d (vjhpkmep8g_u_cizhsw),  
    .x5ug4xxlpdw8ph_oo7x_m (v19st7vd9_bi485e6ak0),  
    .axktcwwx1l7erym3mvldq (zt19omidnr_zyp2gc3bywfb),  
    .fctsirgaydqowic465q   (gccap1c6hft7o1z7esm  ),  
    .u6gfx2g2h7t88vvhusrs5j  (eo5skx1ygvzuasbjgnyl ),  





    .mcnqahf70rz3wm2ilvhef  (1'b0   ), 

    .v1kvt26zg5d2p1i3      (u2a25670eeoaaxpdc   ),
    .z6cksoto8caeb0w8461f     (dl2wnjpp4e2270jy  ),
    .v5l563s9x82qkxwsx    (fy1at1kp6l7l_r5w__q ),

    .r7sap4hhn2lpgz_5t1t      (nruhqt4v8aa4ul498   ),
    .safx984k5yjm7fd8b3i     (sf3mcfi86e2vz   ),
    .pvrou_4d1woq_z6q    (j5zkfgic67jhz8  ),

    .hvxtf10aywneycg3      (aw3rv1bswmks   ),
    .qs405gb8afw52z6eyxi     (etusjysf1bvjmp5   ),
    .e_277pojqob91detq806    (u3fyvcviv3tk65gmcth  ),

    .owijmnymkyht7li_w68  (u6xwpg4na3rdoy), 
    .a3ns4toutens4xm0pf6a  (), 
    .i_2sypygf_zqo5p_t7fy   (pu89y6we99g ),

    .seccdclbkfl          (a42c0ps3vi3       ),
    .g6hr2opjly0         (p7165rjkv      ),
    .l9193amyxxm9g          (h5i09w3ul0070       ),
    .gehkicmawq02an4         (il76519zb__bx      ),
    .fcl5ybv5a2t4y          (srr68v2d6ti       ),
    .ukjsioluzl5t         (a2q31s2sx9u1      ),



    .vpzy7702dz4cc20ajy      (vejdvgqormu727s    ),
    .nwd_h3lrfk59xijt4s7qh1     (ar9ro1ql86jzmq_p   ),
    .s0n0jneoy6ez4dfj5y_9eq    (chezfp7x0va2ea9tdq ),
    .sta4f_rkbcr520sb707nff    (qz1gqv6vh5qturw6v1mz  ),
    .ptyuk4efbbdu9asp0b8cmreeh   (ptyuk4efbbdu9asp0b8cmreeh),
    .f71k3zhdtjavw19c52g45       (f71k3zhdtjavw19c52g45),


    .uy7dkgcktef73e762sbkgdq2teb(qd5sbh8mupp_n4y95vo), 
    .wsnaf53u3elqrc9oym2gh69u5 (fs6jojwsl0l32t7brm38vh ),
    .e49tm9dpy3o9o2w9ac5yowmx (s7vgjm2azmcc3uzzdc_7 ),

    .gf33atgy                 (gf33atgy          ),
    .ru_wi               (ru_wi        ) 
  );



  wire [64-1:0] wtd_nuaeb_mpye;
  wire x7eg618xaszd4f21cl_g;
  wire [64-1:0] cmt_epc;
  wire jlud6jeuxe0espga;







  wire [64-1:0] xd66pm611ai1dg;
  wire r9uxubpl2h2alj1q;
  wire ftp0juzjm2b587cyw5;

  wire sf0uuehfhfa;
  wire hvy2cpsp75f3;
  wire k3z202os;
  wire z35xlcc6bt4;
  wire [64-1:0] ew08uu2kn2p9e11s;
  wire xv08lot3vi9dag4vs0;
  wire [64-1:0] mtc04rctrfyb;
  wire if5jz8qk0aqefy3v35o;


  wire                      rrujrlc85mhm;




  wire                      cmt_dret_ena;
  wire                      s_m3pbf5m2tr6v;



  wire [64-1:0]     unbt3q05xijb;
  wire [64-1:0]     hawbmpz6j7pzibqr;

  wire o7hoht1pqz01v7;
  wire [64-1:0] kbv2bs_lxmvu;

  wire nmi_mode;

  wire status_mie_r;


  wire  x6eltyshbu5;
  wire  lt3v_fm0ipu;
  wire  v3ne7glf8d8;
  wire  v9dnbgjy6c0vf;
  wire  hmzw4exmjn8k921c;


  wire  siifnhwgancn8;
  wire  mfzl2fqml69hx;
  wire  aw0hbwfkx3f63s;
  wire  u83p4flbuvkqt26z;
  wire  tvglhc8o_izdq;

  wire   [64-1:0]     r4bs4k_53n5wp;
  wire   [64-1:0]     i7lgezdqu4bmka;

  wire   [64-1:0]  d3hccrck1fl7jjf6;
  wire                        vkyge0q4mfc5;
  wire   [64-1:0]     cppkd01vpwwnlfy;
  wire   [64-1:0]     h_qwsgi7nk2;
  wire                        w632tcbtqncn6;

  wire                        ai169tbqp4seb3;
  wire                        b0zz_ornhz010;
  wire                        yw4o4kdms07_32;
  wire                        ezl3jzeqhltgj7h;
  wire                        w529wbj853;
  wire                        i9xvsmm45fp0f58;

  wire   [64-1:0]     u25pqekq4df;
  wire                        dhjwho76fa8hqc;
  wire   [64-1:0]     xel6gw173w5x0;
  wire                        icauf4l_12_c2xkj53lf;
  wire   [64-1:0]     v8ydjtlz16x9tx;
  wire                        e_z6d7r9kxqg32te;
  wire   [64-1:0]  p5jpgn4rvarpo;
  wire                        z2g63deibg1b1quqr;
  wire   [64-1:0]     tlgcdv86voe9;
  wire                        u_ufp_wg29ieoklxxz1;


  wire [31:0] xq63jpu81drai3h0;

  wire btwmhh91h50d5flgwx4o6pwu;

  wire xsekawjaoeqedkdymhz6h;
  wire vsrfdna3ksbt8a__05sjdxr;  
  wire uttwdi1xwyv_l7uzt3x2ea;  
  wire d14swmczjaws9gr8uvx;  
  wire fg6gtaxnx8a0anercx;  
  wire [64-1:0] b0cs5n_1_q64sumeg;  

  wire bisaqpu86vneunhkqtg  ;  
  wire m3ar1m0lklmpw4oek2yjd3ev;  
  wire zk19lxmoqrzcdjx6rxuvc36;  
  wire a5_uct872oszxvfp4kn_;  
  wire pl2up5ze0wczfdx0ga70d;  
  wire [64-1:0] jathu3ui07hzkaq4g2z39;  

  wire psx330qmvh5so1to4iq;
  wire sefocn4wjn2k2f_zvlvnz;  
  wire qknomh2kbth19r1osddvzly;  
  wire bzz8x0np0dpmdjt1d0w7uf;  
  wire rl9a96pgy3troiao05jel;  
  wire [64-1:0] hzsp_nydab9ghw59v;  

  wire                     nnk16ophnwar6xhv2v31hjf35p3;  
  wire                     y4lca_o1ofuy216a413i3o;  
  wire                     x_ektinbtzel627cr45gbyrqye;  
  wire                     oi5vxgfcm0z4x5dvik_u6e_io;  
  wire [64-1:0] v37l93ums3fsmtje07   ;  
  wire                     y1cnmq2kze7nro8ev4b35agzl   ;  
  wire                     qufcxlv4zuihmld54ekoij4_e   ;  
  wire                     k3agjwljluupidx6jwin4j65e3j;
  wire                     ytbj92pm9mu_dvm2az0_iv0_72b8i6;
  wire [27-1:0] l_ttwmgineb0ow0w2l5m45r;
  wire [16-1:0] dt6wrpownw18rsx92vw6c1s_9s77; 


  wire                     u645al8bk5q7om05gqugh9ax6_;  
  wire                     zkhpxi7xn6l41mew4wcpsx;  
  wire                     ok06ota43enqbwt1an9er8;  
  wire                     u5hcem386u3f10aew2x9gw9uo5;  
  wire [64-1:0] q17cphsh8955gz9080   ;  
  wire                     dkrri4x05hgshzt6j031fbuc4   ;  
  wire                     c4e63_80r2ix7iqdtrhc   ;  
  wire                     ddzf4jp_h1sxj5bmo1niv6h85uu;
  wire                     qakv1ubh3s9rh1m7l0326d6y2ht7ji73d;
  wire [27-1:0] ks_o8hwsw7nutxfs49acle9i_;
  wire [16-1:0] zi809wzkq9pzbrt3xizvo9uld; 



  assign y_jjs1fut37ilha91qtxkacsoxy = g_wqbz93wfi5bmx7bczdub7 ? sp1w3gxueck6hge7wiki : oungyftsa5o1qeiq0zbvzw5f;

  wire [11:0] k3cmpuswk7in0u4;

  wire w2fpnf5fg1byp6;

  wire apid0ys34zyekptw7un;

  wire [64-1:0] lovkp0eqfnxtb7;

  wire cuxedtph_mmf5zt;
  wire axp009bfo575n9sjnnf;
  wire [5-1:0] brl3pfi8fhhizf3u;
  wire [64-1:0]          zcfxekf7ptrviima;

  ycwy7frvptowq59s2 u_ux607_exu_commit(
      .se2buoxmq91dbic3y2m5hu (se2buoxmq91dbic3y2m5hu),
      .e9u0rtvt8jrygyc8s     (e9u0rtvt8jrygyc8s),
      .lovkp0eqfnxtb7     (lovkp0eqfnxtb7),

    .a02zzbowpjn06h   (a02zzbowpjn06h),

    .feq1g7m2cy1erl     (feq1g7m2cy1erl),

    .k3cmpuswk7in0u4     (k3cmpuswk7in0u4),

    .av1w8ld09cfofn     (av1w8ld09cfofn    ),
    .im2b5l0h98avl6t4sj (im2b5l0h98avl6t4sj),
    .bw65wl7fvekfymd8vqx  (bw65wl7fvekfymd8vqx ),
    .pecbpcoa04vq      (pecbpcoa04vq     ),
    .tb_snaxyfs       (tb_snaxyfs      ),
    .zc4mldgm25r      (zc4mldgm25r     ),
    .d23wb5yh1iyvf      (d23wb5yh1iyvf     ),
    .srim3bfnzhve       (srim3bfnzhve      ),
    .fvqwdz2hdbb      (fvqwdz2hdbb     ),
    .cy3nuhzm_v2p73mt  (cy3nuhzm_v2p73mt ),  

    .btwmhh91h50d5flgwx4o6pwu(btwmhh91h50d5flgwx4o6pwu),
    .tywculgjyor8ndw    (tywculgjyor8ndw   ),
    .xq63jpu81drai3h0 (xq63jpu81drai3h0),
    .r21i4by0bu3ks             (r21i4by0bu3ks),


    .tw5xnp59d8x            (tw5xnp59d8x        ),
    .af5qc04tmn51e4u2h1z    (af5qc04tmn51e4u2h1z),

    .qo5p9t6s74zxpo         (qo5p9t6s74zxpo),

    .w2fpnf5fg1byp6      (w2fpnf5fg1byp6),


    .h7fseh5_df0hbx         (h7fseh5_df0hbx),

    .uc5qxb4d2b28ye5          (uc5qxb4d2b28ye5),
    .o2qkf90r783          (o2qkf90r783),

    .apid0ys34zyekptw7un       (apid0ys34zyekptw7un),
    .um8zsjyxn_4p             (um8zsjyxn_4p      ),  


    .qwcb6hcmvfqmf032z    (qwcb6hcmvfqmf032z),
    .woon4h3ivznl_qiu7i_9    (woon4h3ivznl_qiu7i_9),
    .y_0q8d40rrzolo1y6    (y_0q8d40rrzolo1y6),
    .ao17frh5wnr0wddz3    (ao17frh5wnr0wddz3),
    .p25dd0cxz7nmi6w9ebukmr   (hno6u0yd_gjy_1t),
    .uvgy9al0j8prciqsh      (ppx8euepv0evvizd),
    .f8pn1x6gurodpy04d3j1ihn   (f1yknbdsst7yvsgvm210),
    .mmludd_fnt2yevok8a1a0    (mmludd_fnt2yevok8a1a0),
    .buwj9_8l8bwj80kkinq9p    (buwj9_8l8bwj80kkinq9p),

    .c5ewdqztjw9za (c5ewdqztjw9za),
    .rn2mt6nngsc9w5cz(rn2mt6nngsc9w5cz),
    .fcjh1nct4r (fcjh1nct4r),
    .b4lwcgm6l21pi(b4lwcgm6l21pi),
    .zwcbp7zqfei5xz(zwcbp7zqfei5xz),
    .dz0zrf512290tvcy4q(dz0zrf512290tvcy4q),
    .z0yhjfv_e0yaa2r(z0yhjfv_e0yaa2r),
    .dn8riluj40uunvq5(dn8riluj40uunvq5),
    .w632tcbtqncn6         (w632tcbtqncn6    ),
    .ai169tbqp4seb3            (ai169tbqp4seb3       ),
    .b0zz_ornhz010            (b0zz_ornhz010       ),
    .yw4o4kdms07_32            (yw4o4kdms07_32       ),
    .ezl3jzeqhltgj7h            (ezl3jzeqhltgj7h       ),
    .w529wbj853            (w529wbj853       ),
    .i9xvsmm45fp0f58            (i9xvsmm45fp0f58       ),
    .r4bs4k_53n5wp         (r4bs4k_53n5wp    ),
    .jqsukc5b5drcc1e78        (jqsukc5b5drcc1e78   ),
    .gnn46rd7vvofruqij        (gnn46rd7vvofruqij   ),
    .vkyge0q4mfc5          (vkyge0q4mfc5     ),
    .cppkd01vpwwnlfy           (cppkd01vpwwnlfy      ),
    .d3hccrck1fl7jjf6          (d3hccrck1fl7jjf6     ),
    .h_qwsgi7nk2           (h_qwsgi7nk2      ),
    .u25pqekq4df            (u25pqekq4df       ),
    .dhjwho76fa8hqc        (dhjwho76fa8hqc   ),
    .xel6gw173w5x0           (xel6gw173w5x0      ),
    .icauf4l_12_c2xkj53lf       (icauf4l_12_c2xkj53lf  ),
    .v8ydjtlz16x9tx          (v8ydjtlz16x9tx     ),
    .e_z6d7r9kxqg32te      (e_z6d7r9kxqg32te ),
    .p5jpgn4rvarpo              (p5jpgn4rvarpo         ),
    .z2g63deibg1b1quqr          (z2g63deibg1b1quqr     ),
    .tlgcdv86voe9          (tlgcdv86voe9     ),
    .u_ufp_wg29ieoklxxz1      (u_ufp_wg29ieoklxxz1 ),
    .rn1o3sl83              (rn1o3sl83),
    .z1l80uwh6vyyg34          (z1l80uwh6vyyg34),

    .s5f_36xvqrtq7          (status_mie_r),

    .x6eltyshbu5            (x6eltyshbu5        ),
    .lt3v_fm0ipu            (lt3v_fm0ipu        ),
    .v3ne7glf8d8            (v3ne7glf8d8        ),
    .v9dnbgjy6c0vf          (v9dnbgjy6c0vf      ),
    .hmzw4exmjn8k921c           (hmzw4exmjn8k921c       ),

    .siifnhwgancn8            (siifnhwgancn8        ),
    .mfzl2fqml69hx            (mfzl2fqml69hx        ),
    .aw0hbwfkx3f63s            (aw0hbwfkx3f63s        ),
    .u83p4flbuvkqt26z          (u83p4flbuvkqt26z      ),
    .tvglhc8o_izdq           (tvglhc8o_izdq       ),
    .gkjb6c98b5j1zsgbv26       (leq1ne49igptrh__p_5kz23048rjzm),
    .unntlrmfpzgdq8rnz3ug3_8    (ipj0pyjf76qkv519em1jiaiutbhsr),
    .n9q1kib2q28tfyzyue2j2or   (szaorjzmus1ssgjq7e30bdssuadwt0  ),
    .asxvrob6s2_85u99em22   (yi0r5xirgktqhr99j3jz345g11t51  ),
    .bva3_s2oj2hgomj0eyrk   (ogkluwmj9mmpgtmicjnh6_yya46ukkp2s  ),
    .fbgda1d6z8gr725snyc2ylc  (d250junaig195xflrdmkjjl5pxtaf4),

    .s_qow7tm_gendxgd          (yh8eetxf0xs392       ),
    .j_v6uy8_pdqb7w              (jwbql4ta0c           ),
    .t3xakjcvvthgm_v0            (omler2igyskatx         ),

    .tb198r6lzk1sr77g4        (tb198r6lzk1sr77g4   ),
    .cvvsn7xc8qg5uk            (cvvsn7xc8qg5uk       ),
    .pc67uztpd_zg6bsal          (pc67uztpd_zg6bsal     ),

    .q23hngbyy69cc9ci9sjr8g4     (ap889z2q8jbzn4dhurkzl  ),
    .vqv5qr4a5j6difuyllem3ur_ (y_jjs1fut37ilha91qtxkacsoxy),
    .rnodgdrxyr_tulm0nnnign     (rnodgdrxyr_tulm0nnnign),

    .d3n7pwgwcgze9cr4         (j39tby_g7kqga33w_m      ),
    .cphtk1_x8fwehad         (t0o4cn_ndv2lmnp      ),
    .amc4c8vcbecv1i            (my5_v4hhb7oc51         ),
    .qgp6cehpls743wtn0i         (lmv45fhtl015bg      ),
    .ama4p78xalq9j32         (uv_3uzx5ti04u5nd      ),
    .zcldu5wj7n47pd36vbj        (aa5a1tnclwe351p5ujs     ),
    .d0e2kztse3ur2dt22q       (yd4wqg2e0i386ccq6y9    ),
    .y4fasvbsps__6yzpqc7eymh     (tv3_4qrynvnaoy4riz  ),
    .k_5q95o2gjo1w_rk          (y_gvnr7uidhcof1       ),
    .f_4x5ty4man9f87i           (zh_0_4wrffapmbs        ),
    .uzhgx8hpcw0vcm6nfex          (nrze6rcjz4m65z        ),
    .ichypldcqgx_6hsv           (cjxy_cr6jzz17mr8         ),
    .mn3xo91xnxw486688t           (g0ovdu1w9dcoqg         ),
    .omxbj0blxqsqi9h          (uxdt29u4dd96ukc        ),
    .c4mm5jszl6uvumay          (r_cdggxn_7syt0g        ),
    .npbrk566oq0dkbf982i          (cmv9vkluc86swnlc        ),
    .wyutdg78_ykde5xhd          (uvw8h6lqr2ou0        ),
    .gqwf5n54sp4jlral         (rwip45nhuhbz2jkd4      ),
    .eo9f914sbhga72uw1z        (x3r6u6q7ck5ud8wbii     ),
    .qa04tbszp_crup1y4rvk        (p0ga7mahvd8zjma     ),
    .p38eaxsiobphopbri        (hlxcm16byj04fp0     ),
    .jw67do539fm4kvlowut9k62      (o4lqcf45nah3boccbw   ),
    .yhg7so3hz941h           (alu_cmt_wfi     ),
    .xi8b7jmwma99a4gxgmri9v74   (alu_cmt_ifu_misalgn),
    .g0esgcmgdknyveiq2t72xopfk    (qjg3a6detqucp4byrgs ),
    .v1vwaj41ljxavm9366uapnar1zrk5(qn6g68ul7q8pz3pvopdmh0m),
    .o4512597_0nxc_jrf287w8it    (kxmzp6o3alj05dfq9d_e8ci ),
    .l4km4217yp2p969cwda8    (d2gcdo57ra3yxudimcwal0 ),
    .ugimrlqwlbs5gblkxuymto1h4  (ob__kc7kdtjxp74ajo7ql548o),
    .xktv6472l59a_iqmuyhu     (v85ovm_7gp20oi4vj  ),

    .p27tnvqrliur1xjlr527b   (ihmezohdr7mg9_blli7),
    .rx_c151de4k7bbwnwrak    (ctgxr_wil90tj1ur64),
    .k3t4av4o2bjnmmpxdoqfumyxecc09u7q5h(oozkxp7aywu4l0hz73uedbtyiad ),
    .n3tpm7ps0ygbm4a_yr6ryn06egc1(j5wtbhk36xx9j2h1kgsniu9p0d9xzj),
    .bnta1_ctyuyz6f0cs2zpyuy2nmfjv4(qh0m9d6yrl5kb_1vvecw1kb1wrbm),
    .rgf8gwy5mb_doix8zdjh30tiklwj  (kihyrfzcb87yz3qnxq7c0o11at5u  ),
    .khjs1qtt_oec9bu6269tck93yo8gpdw  (ho49hpl6ijpiop4thzf8rh6apio4u  ),
    .k7nmctokgpx6dz4ugb1i3zr9q20f  (wk2sssl74c1xyhbm7pf29qtbpws1  ),
    .awq_rxiss6jp46gvm3g      (vxcgun4z0ztx7nmvm   ),
    .rgsv1cqeh7x_1ex_5tj      (fq2y4oplmud5drf9s   ),

    .kdofxulgpcpa9q310       (oa_1ibjpvwpv6bg5ivcau2uo6z3s),
    .e9g0sper1c9v_vmf            (noc4nf4qform41kyqw6m4     ),
    .xv88qbq7hr0lskm4cqrn         (ktqyocabrct3iqhlj18u9fhnz6f3d  ),
    .zjuaef59fqixf4nfbc        (ihbxqlci_5lmn6uyuoxv158n18bua ),
    .yy8cmh_xtnis7nqw_60        (xv9g6nf92837e31mav06v03y2t ),
    .t73hv26oh7wdnclcbf5b6j9  (cuxedtph_mmf5zt            ),
    .zi6t1yvku2qc168r2cv9b4v10vi6ee7(axp009bfo575n9sjnnf    ),
    .fuvqsp044l3a4fk69bkuvqopz0 (brl3pfi8fhhizf3u             ),
    .pji7j1gx57ht5kwknem7at7  (zcfxekf7ptrviima              ),
    .o09mrpo1o2k6w4jsat2_o       (ppwfzi9r2pfdu5oiww3x5a9g94u6ut0),

    .qqlnmd2zlr98m5mdjyk     (ne5matgyfjvw3elazxt7p),
    .dxvoc8nirjgo0by0yoex4l01a7  (tpd5fcgyg_240nz8md69oj  ), 
    .cqlsgy50_6bt6xavc02vpsg9p(npkoy9e2dsczayfq7h6cko59),
    .iby9hp5grzp4ouc82c61kxa    (kmlf0ops49wvgcz2howfob59khsqir  ), 
    .mpp5ftr3blzju24mrjjk4nv  (kw590mop2ic8u619z7c_owrnv9t), 



    .gkhcosyb6da4dfdhh3       (apf9b6zz11802cqi     ),
    .qgf355r7t8juyfmkx9g       (trff4kgfudc86mj     ),
    .troptfm3sc9gj8rb         (v_t46_oqiae0c4es9uht   ),
    .d_4gaf_5w4wygi9         (xw9obr7t22kfov7grph7   ),



    .i32x_jtt7bvmr9lu2p    (pbtolkl953sk14id0iy  ),
    .mxa77etukhs8o_5z6962l19    (z2qyay491938ppnlxuc  ),
    .cd4v4c_rw906kt5       (zeseql2htbxpugyu5_j     ),
    .idat72abxke4z9s       (al3t866kz4po45vfuyjy     ),
    .hv4wuttuo9jk_cqa8sxqwt   (xutsaulafh4onxtthm8n ),
    .ac8_dky9fhpbsxu0b9t88ag8   (me7unt7fapqqhtc6epso ),
    .r_8f7p3tznijza5y03ko  (m2as3qe7miuhj662j1zvt),

    .pydatzxqqi              (pydatzxqqi),

    .qeb3z0x5               (qeb3z0x5        ),
    .ibhfuwrztbm8p4gg           (ibhfuwrztbm8p4gg    ),
    .i8_5wt0vppx            (i8_5wt0vppx     ),
    .osv2437qj_3nuf        (osv2437qj_3nuf ),


    .b7g_vsn0zoewh6g1          (b7g_vsn0zoewh6g1),
    .onnv64ydiajl              (onnv64ydiajl    ),
    .t5trf35s8vy            (t5trf35s8vy),
    .zbac123pv78sbz3         (zbac123pv78sbz3),
    .z4e_m564fxae0kpbjr         (z4e_m564fxae0kpbjr),
    .hixy2y36a1pn0         (hixy2y36a1pn0),
    .ozwene1gdpatk6g            (ozwene1gdpatk6g   ),

    .azll7rq5fab5ou      (azll7rq5fab5ou      ),
    .n6a0r_0zddzrme8      (n6a0r_0zddzrme8      ),
    .ns0i7siujgkrghjpqv6(ns0i7siujgkrghjpqv6),

                           

    .c4ughu0qm5sfai          (c4ughu0qm5sfai),

    .um28jgd2x4mbs            (1'b0), 
    .aw82i964do                (aw82i964do),
    .cwwkpmk260lrt              (nmi_mode),
    .rvr30vvllni            (rvr30vvllni),
    .z1cj655u31            (z1cj655u31),
    .y8_gkxsfle                (y8_gkxsfle),
    .lhu2z948o3n            (lhu2z948o3n),


    .wtd_nuaeb_mpye           (wtd_nuaeb_mpye    ), 
    .x7eg618xaszd4f21cl_g       (x7eg618xaszd4f21cl_g),
    .elth4vimq_j               (cmt_epc        ),
    .jlud6jeuxe0espga           (jlud6jeuxe0espga    ),






    .xd66pm611ai1dg             (xd66pm611ai1dg      ),
    .r9uxubpl2h2alj1q         (r9uxubpl2h2alj1q  ),
    .ftp0juzjm2b587cyw5       (ftp0juzjm2b587cyw5  ),

    .sf0uuehfhfa              (sf0uuehfhfa       ),
    .hvy2cpsp75f3               (hvy2cpsp75f3        ),
    .k3z202os              (k3z202os       ),
    .z35xlcc6bt4               (z35xlcc6bt4        ),
    .ew08uu2kn2p9e11s           (ew08uu2kn2p9e11s    ),
    .xv08lot3vi9dag4vs0       (xv08lot3vi9dag4vs0),
    .mtc04rctrfyb          (mtc04rctrfyb    ),
    .if5jz8qk0aqefy3v35o      (if5jz8qk0aqefy3v35o),

    .jw4fsjecr0u919fr7            (cmt_dret_ena     ),
    .rrujrlc85mhm            (rrujrlc85mhm     ),
    .s_m3pbf5m2tr6v            (s_m3pbf5m2tr6v     ),
    .bde41te346q515l              (bde41te346q515l       ),
    .gfod0nmy6eta29jeeg6mr2      (u_hs70f19eo9kuxrncia   ),
    .n4soswat5yihd74b         (gqxkhqynd510udp0tpbr),      
    .y8wz7aud_fd6dfiakjtx2i0g   (y8wz7aud_fd6dfiakjtx2i0g),
    .dgnjyd9xs8efyxm0tdlsvfq4eop  (dgnjyd9xs8efyxm0tdlsvfq4eop),
    .a3xib90kwk4_hm1         (akig71_dnhvxrc3d3u_de),
    .nfzexr8q9g893gi          (w9z2kr44j8w6w3w1zqa),
    .opkkwp3eg8g3448t         (q94xtoze0utbz_anbev),
    .tv3_4qrynvnaoy4riz           (e43glfkwrdo0_s ),



    .pldoasxyzlvx2              (pldoasxyzlvx2       ),

    .hn85hkp2yav               (hn85hkp2yav       ),
    .o7hoht1pqz01v7            (o7hoht1pqz01v7),
    .kbv2bs_lxmvu             (kbv2bs_lxmvu ),
    .unbt3q05xijb             (unbt3q05xijb     ),
    .hawbmpz6j7pzibqr             (hawbmpz6j7pzibqr),

    .v35y3qnk7mx3l1695       (v35y3qnk7mx3l1695    ),

    .zsgl59ydqwjln          (zsgl59ydqwjln    ),
    .b9yq2alidby7zgom1          (lkvz9_caztnpkd5y1a    ),
    .tvqijouldcgiz2dxdco7     (nnk16ophnwar6xhv2v31hjf35p3),  
    .zkxlkidschdubxpkpm     (y4lca_o1ofuy216a413i3o),  
    .xmcrni1qngfvh9pil9j     (x_ektinbtzel627cr45gbyrqye),  
    .btkcf2uqr61gkiqhde0lai     (oi5vxgfcm0z4x5dvik_u6e_io),  
    .h01d94xsxbxe_req           (v37l93ums3fsmtje07),  
    .w1casjl7bz73brz       (y1cnmq2kze7nro8ev4b35agzl),  
    .hjri7cufo9ckntq         (qufcxlv4zuihmld54ekoij4_e),  
    .yghffofulqa77bd7aw07badta1a  (k3agjwljluupidx6jwin4j65e3j  ),
    .rrl7evvmayt1_vvp74iq9h6_cjf(ytbj92pm9mu_dvm2az0_iv0_72b8i6),
    .zddoxp22m1o11x30gbe      (l_ttwmgineb0ow0w2l5m45r      ),
    .hwfethpzkuauejcgtbl6o    (dt6wrpownw18rsx92vw6c1s_9s77    ),  

    .n3ak8l6cvn0s4            (n3ak8l6cvn0s4     ),
    .hsxh9536ho4bw8o            (dvloyy6lickuq8759jcfc6     ),
    .r_edve7v9jcr26q6zk       (u645al8bk5q7om05gqugh9ax6_),
    .vrqfzuog2k4pos133       (zkhpxi7xn6l41mew4wcpsx),
    .bmw2yi333716crywk       (ok06ota43enqbwt1an9er8),
    .k2sr7sw1plcmnki5ajtscw       (u5hcem386u3f10aew2x9gw9uo5),
    .jkzw_f9anx55             (q17cphsh8955gz9080      ),
    .t8muv9e6d7yk_whqa0         (dkrri4x05hgshzt6j031fbuc4),  
    .hzdfp71n6g3f5fsg5         (c4e63_80r2ix7iqdtrhc),  
    .lwdhmuzyvcvv14mjbl0h2a41z  (ddzf4jp_h1sxj5bmo1niv6h85uu  ),
    .xy48dugh009wtmazqug3kpy2a5h_(qakv1ubh3s9rh1m7l0326d6y2ht7ji73d),
    .l4ztejmt2__wxqm2rw      (ks_o8hwsw7nutxfs49acle9i_      ),
    .s3ujdp2a8n69bm6engxok    (zi809wzkq9pzbrt3xizvo9uld    ),  

    .xsekawjaoeqedkdymhz6h       (xsekawjaoeqedkdymhz6h  ),
    .vsrfdna3ksbt8a__05sjdxr     (vsrfdna3ksbt8a__05sjdxr),  
    .uttwdi1xwyv_l7uzt3x2ea     (uttwdi1xwyv_l7uzt3x2ea),  
    .d14swmczjaws9gr8uvx     (d14swmczjaws9gr8uvx),  
    .fg6gtaxnx8a0anercx     (fg6gtaxnx8a0anercx),  
    .b0cs5n_1_q64sumeg        (b0cs5n_1_q64sumeg   ),  

    .bisaqpu86vneunhkqtg       (bisaqpu86vneunhkqtg  ),
    .m3ar1m0lklmpw4oek2yjd3ev     (m3ar1m0lklmpw4oek2yjd3ev),  
    .zk19lxmoqrzcdjx6rxuvc36     (zk19lxmoqrzcdjx6rxuvc36),  
    .a5_uct872oszxvfp4kn_     (a5_uct872oszxvfp4kn_),  
    .pl2up5ze0wczfdx0ga70d     (pl2up5ze0wczfdx0ga70d),  
    .jathu3ui07hzkaq4g2z39        (jathu3ui07hzkaq4g2z39   ),  

    .psx330qmvh5so1to4iq       (psx330qmvh5so1to4iq  ),
    .sefocn4wjn2k2f_zvlvnz     (sefocn4wjn2k2f_zvlvnz),  
    .qknomh2kbth19r1osddvzly     (qknomh2kbth19r1osddvzly),  
    .bzz8x0np0dpmdjt1d0w7uf     (bzz8x0np0dpmdjt1d0w7uf),  
    .rl9a96pgy3troiao05jel     (rl9a96pgy3troiao05jel),  
    .hzsp_nydab9ghw59v        (hzsp_nydab9ghw59v   ),  

    .qk0jm7flfzap             (ngy4ipxc1vxym69lu),
    .fj4fje1ckitqjb_7        (xmi2_r3_mwq_b4a70u_m),
    .nes78rg61lk5t2            (bjqlln4lucs2dyr),

    .dk2xhkj77a                 (dk2xhkj77a      ),
    .gf33atgy                     (gf33atgy          ),
    .ru_wi                   (ru_wi        ) 
  );

    
    assign b9yq2alidby7zgom1       =  lkvz9_caztnpkd5y1a ;
    assign tvqijouldcgiz2dxdco7  =  lkvz9_caztnpkd5y1a ? nnk16ophnwar6xhv2v31hjf35p3 : 1'b0;  
    assign zkxlkidschdubxpkpm  =  lkvz9_caztnpkd5y1a ? y4lca_o1ofuy216a413i3o : 1'b0;  
    assign xmcrni1qngfvh9pil9j  =  lkvz9_caztnpkd5y1a ? x_ektinbtzel627cr45gbyrqye : 1'b0;  
    assign btkcf2uqr61gkiqhde0lai  =  lkvz9_caztnpkd5y1a ? oi5vxgfcm0z4x5dvik_u6e_io : 1'b0;  
      assign h01d94xsxbxe_req        =  lkvz9_caztnpkd5y1a ? v37l93ums3fsmtje07    : 64'h0    ;  
      assign w1casjl7bz73brz    =  lkvz9_caztnpkd5y1a ? y1cnmq2kze7nro8ev4b35agzl: 1'b0;  
      assign hjri7cufo9ckntq    =  lkvz9_caztnpkd5y1a ? qufcxlv4zuihmld54ekoij4_e: 1'b0;  
      assign yghffofulqa77bd7aw07badta1a    = lkvz9_caztnpkd5y1a ? k3agjwljluupidx6jwin4j65e3j   : 1'b0;
      assign rrl7evvmayt1_vvp74iq9h6_cjf  = lkvz9_caztnpkd5y1a ? ytbj92pm9mu_dvm2az0_iv0_72b8i6 : 1'b0;
      assign zddoxp22m1o11x30gbe        = lkvz9_caztnpkd5y1a ? l_ttwmgineb0ow0w2l5m45r       : {27{1'b0}};
      assign hwfethpzkuauejcgtbl6o      = lkvz9_caztnpkd5y1a ? dt6wrpownw18rsx92vw6c1s_9s77     : 16'b0;

    assign hsxh9536ho4bw8o       =  (dvloyy6lickuq8759jcfc6 | qfspmfi47b5jx99i0);
    assign r_edve7v9jcr26q6zk  =  dvloyy6lickuq8759jcfc6 ? u645al8bk5q7om05gqugh9ax6_ : pjcdn7d17lcskz8qw3fi;  
    assign vrqfzuog2k4pos133  =  dvloyy6lickuq8759jcfc6 ? zkhpxi7xn6l41mew4wcpsx : c3edim0hxqlxh7ubn4hn;  
    assign bmw2yi333716crywk  =  dvloyy6lickuq8759jcfc6 ? ok06ota43enqbwt1an9er8 : seyk3b__57tr0b_kv__y;  
    assign k2sr7sw1plcmnki5ajtscw  =  dvloyy6lickuq8759jcfc6 ? u5hcem386u3f10aew2x9gw9uo5 : 1'b0;  
      assign jkzw_f9anx55        =  dvloyy6lickuq8759jcfc6 ? q17cphsh8955gz9080    : bymbiaovszt6x5okz    ;  
      assign t8muv9e6d7yk_whqa0    =  dvloyy6lickuq8759jcfc6 ? dkrri4x05hgshzt6j031fbuc4: qb0v08s4r8feqekkzsn;  
      assign hzdfp71n6g3f5fsg5    =  dvloyy6lickuq8759jcfc6 ? c4e63_80r2ix7iqdtrhc: uyh4zz3rdydme0z8m4r;  
      assign lwdhmuzyvcvv14mjbl0h2a41z    = dvloyy6lickuq8759jcfc6 ? ddzf4jp_h1sxj5bmo1niv6h85uu   : 1'b0;
      assign xy48dugh009wtmazqug3kpy2a5h_  = dvloyy6lickuq8759jcfc6 ? qakv1ubh3s9rh1m7l0326d6y2ht7ji73d : 1'b0;
      assign l4ztejmt2__wxqm2rw        = dvloyy6lickuq8759jcfc6 ? ks_o8hwsw7nutxfs49acle9i_       : {27{1'b0}};
      assign s3ujdp2a8n69bm6engxok      = dvloyy6lickuq8759jcfc6 ? zi809wzkq9pzbrt3xizvo9uld     : 16'b0;


  assign d3n7pwgwcgze9cr4 = j39tby_g7kqga33w_m;
  assign amc4c8vcbecv1i    = my5_v4hhb7oc51   ;




  assign yhbtmo4kyz_ewog3  = gkx4s0wv_05dt7e ;
  assign cd4d2_i3rcc1_p = f9_w27gbcq__  ;
  assign wyu42gj62n994v0wo_ = lnwarwpyiph_rhx;
  assign lz3vnoxnz_z    = f_ljupvj_wh;



  wire elspwgn4qhqqwg31epb = (|chezfp7x0va2ea9tdq);

  assign st4f16aums5 = aw82i964do;
  assign p05ld2ghmwh = y8_gkxsfle;


  nrcp90w_wy4yo u_ux607_exu_csr(
      .pby60vfdze02     (pby60vfdze02),
      .vm3pyzc9nt95     (vm3pyzc9nt95),
      .vdr9fi9zwq         (y_gvnr7uidhcof1),
      .rbz4pv_atxqopdwt     (rbz4pv_atxqopdwt),
      .qs1xgat7r8xow     (qs1xgat7r8xow),
      .lovkp0eqfnxtb7     (lovkp0eqfnxtb7),
      .vyxop00ua6vr     (vyxop00ua6vr),
      .p6rw9no76a3m       (p6rw9no76a3m),
      .nchi0_6mu           (my5_v4hhb7oc51),
      .w92a5o09fp9dg6    (w92a5o09fp9dg6   ),
      .eglor15f7p2ivpny5dc    (eglor15f7p2ivpny5dc   ),
      .ous_emkpecrqhg5e7 (ous_emkpecrqhg5e7),
      .doh50j3p7c7yl7uk9 (doh50j3p7c7yl7uk9),
      .exltui35irvvmodu205vw (exltui35irvvmodu205vw ),
      .s7eq8f6z1uyi2in    (s7eq8f6z1uyi2in    ),
      .qbsr1jytrqtsbk4ttb8nz(qbsr1jytrqtsbk4ttb8nz),
      .btwmhh91h50d5flgwx4o6pwu(btwmhh91h50d5flgwx4o6pwu),
      .zz5wo47gw146x4        (zz5wo47gw146x4),
      .fgr486jx5kevbua        (fgr486jx5kevbua),
      .pvfk1_6o89lmby         (pvfk1_6o89lmby),
      .xx87vzbpchg         (xx87vzbpchg),

      .apid0ys34zyekptw7un   (apid0ys34zyekptw7un),

      .k3cmpuswk7in0u4     (k3cmpuswk7in0u4),

      .xsekawjaoeqedkdymhz6h   (xsekawjaoeqedkdymhz6h  ),
      .vsrfdna3ksbt8a__05sjdxr (vsrfdna3ksbt8a__05sjdxr),  
      .uttwdi1xwyv_l7uzt3x2ea (uttwdi1xwyv_l7uzt3x2ea),  
      .d14swmczjaws9gr8uvx (d14swmczjaws9gr8uvx),  
      .fg6gtaxnx8a0anercx (fg6gtaxnx8a0anercx),  
      .b0cs5n_1_q64sumeg    (b0cs5n_1_q64sumeg   ),  

      .bisaqpu86vneunhkqtg   (bisaqpu86vneunhkqtg  ),
      .m3ar1m0lklmpw4oek2yjd3ev (m3ar1m0lklmpw4oek2yjd3ev),  
      .zk19lxmoqrzcdjx6rxuvc36 (zk19lxmoqrzcdjx6rxuvc36),  
      .a5_uct872oszxvfp4kn_ (a5_uct872oszxvfp4kn_),  
      .pl2up5ze0wczfdx0ga70d (pl2up5ze0wczfdx0ga70d),  
      .jathu3ui07hzkaq4g2z39    (jathu3ui07hzkaq4g2z39   ),  

      .w2fpnf5fg1byp6(w2fpnf5fg1byp6),
      .x_cq40qmp6a  (x_cq40qmp6a), 

      .wd9dvepxj     (wd9dvepxj),

      .xq63jpu81drai3h0 (xq63jpu81drai3h0),


      .habgbg2jn3qi     (habgbg2jn3qi),
      .dg4hzu_          (dg4hzu_     ),
      .h7fseh5_df0hbx     (h7fseh5_df0hbx),
      .wj5ypo5k        (zc9t_vib9_fw44d),









      .ix299qulxi5            (ix299qulxi5    ),
      .jjj61w03m77lv           (jjj61w03m77lv    ),
      .enwn0u48p2_ls5az80          (enwn0u48p2_ls5az80),
      .f_i1959b4xizzq9jea           (f_i1959b4xizzq9jea),
      .b4lwcgm6l21pi          (b4lwcgm6l21pi),
      .hjrk_rwjkqj3zk_b         (hjrk_rwjkqj3zk_b),
      .zwcbp7zqfei5xz         (zwcbp7zqfei5xz),
      .znzjygllppv1s0a8cqub3c    (znzjygllppv1s0a8cqub3c), 
      .gfy3zost37aq8qmr          (gfy3zost37aq8qmr),
      .dxi_ue3gf5zqqqxwgq2a    (dxi_ue3gf5zqqqxwgq2a),
      .dn8riluj40uunvq5        (dn8riluj40uunvq5),
      .z0yhjfv_e0yaa2r          (z0yhjfv_e0yaa2r),
      .guuvp01vkcryglsu1p3    (guuvp01vkcryglsu1p3),
      .hig2gwwbeuhnt65xrp        (hig2gwwbeuhnt65xrp),


      .pcr4upio7_tx37     (pcr4upio7_tx37   ), 
      .uzklqlncpqqm1rav  (uzklqlncpqqm1rav),
      .ortueunvnkx_l5m_j  (ortueunvnkx_l5m_j),
      .hwuhtb7ucto_utk56  (hwuhtb7ucto_utk56),
      .i1env2kmns7qvvuuc  (i1env2kmns7qvvuuc),
      .g3s3vpafvy3i  (g3s3vpafvy3i),


      .rm1dxjejhq7dh3q5m  (rm1dxjejhq7dh3q5m ),

    .r0s7d8cr68i2qs1z     (r0s7d8cr68i2qs1z),
    .kakelc68be0x7tdm9b9o    (kakelc68be0x7tdm9b9o),
    .j3j1czgoam48vhs8auo    (j3j1czgoam48vhs8auo),
    .gm1r5itc44uxw_y0_msk    (gm1r5itc44uxw_y0_msk),

    .canacnkc7zibtkn418i                 (canacnkc7zibtkn418i                ), 
    .x8rpm78rvvycis                      (x8rpm78rvvycis                     ), 
    .bwbmafs1inesgjyn                      (h7lpiwlxyb79qyr06                     ), 
    .bkkiffh6ob85nh79doya_                 (bkkiffh6ob85nh79doya_                ), 
    .qhqqh0lyehgtfop1tc                 (qhqqh0lyehgtfop1tc                ), 
    .x03ux1utw4qem5kk3c                 (x03ux1utw4qem5kk3c                ), 
    .sxhicsqvufwfbnk0                      (sxhicsqvufwfbnk0                     ), 
    .ydydp69z03wvr97                      (c5wzn6bil69i9toc                     ), 
    .pjic5x84bqxpvdduy4r2s                 (pjic5x84bqxpvdduy4r2s                ), 
    .w5az87bw32r0tjbo0tdrv2ouvx            (w5az87bw32r0tjbo0tdrv2ouvx           ), 

    .vs6ryzcr0bwqs5so                   (vs6ryzcr0bwqs5so                  ), 
    .j25ub196dc_agl8oovaex4                  (j25ub196dc_agl8oovaex4                 ), 
    .pi2nokcm8qf7och7l4g                  (pi2nokcm8qf7och7l4g                 ), 
    .c0i0hs5tz64_ce5f0z                 (c0i0hs5tz64_ce5f0z                ), 
    .dmzdczrqcueolg3dzufj_by5rmf            (dmzdczrqcueolg3dzufj_by5rmf           ), 
    .a1sqko6fok9qzpbtyuw0                 (a1sqko6fok9qzpbtyuw0                ), 
    .bquohubxiv2rsayn62v                 (bquohubxiv2rsayn62v                ), 
    .kqyojh1maxy0x834htg                (kqyojh1maxy0x834htg               ), 

    .hpk3eafyque5ubt_c62flnny              (hpk3eafyque5ubt_c62flnny             ),       
    .sfezv1xz2ghvo8pkt                     (sfezv1xz2ghvo8pkt                    ),               
    .vagaza053272juvmo59v8w20s              (vagaza053272juvmo59v8w20s             ),       
    .rzf45534z36ejq96260                  (rzf45534z36ejq96260                 ),       
    .frzfsbt7hp3n4aj3zvvumnh0s               (frzfsbt7hp3n4aj3zvvumnh0s              ),         
    .zkuxqezrmlhyyjjgx                    (zkuxqezrmlhyyjjgx                   ),              
    .u3h5tvu1g2q93141j9o                    (u3h5tvu1g2q93141j9o                   ),              
    .pjh0wad7t_5du3cync_0c              (pjh0wad7t_5du3cync_0c             ),                        
    .wmkgrgf631pbq                      (wmkgrgf631pbq                     ),
    .oyq1p3qa2iffjuqns0jkgg                  (oyq1p3qa2iffjuqns0jkgg                 ),
                                                                           
    .qjw2q0j88rjr42lautsqnca              (qjw2q0j88rjr42lautsqnca             ),       
    .imkm56ujne9v4m6n08w1yf5622           (imkm56ujne9v4m6n08w1yf5622          ),     
    .txk1r9aiq_7l2nkw101w_                (txk1r9aiq_7l2nkw101w_               ),          
    .ih4hmwugasiodbx5da9_40kx               (ih4hmwugasiodbx5da9_40kx              ),        
    .x5vjq7mshfwr0h3q514t7mhdt               (x5vjq7mshfwr0h3q514t7mhdt              ),        
    .qrxtk7e03100_uwkx73sg7               (qrxtk7e03100_uwkx73sg7              ),        
    .i7qiq2q9c6hbeful9qu9lb               (i7qiq2q9c6hbeful9qu9lb              ),         
    .yr0s3skqk7cdqflsrbsxg9znu               (yr0s3skqk7cdqflsrbsxg9znu              ),         
    .adqieke11qo0elfz93hlouwjc0         (adqieke11qo0elfz93hlouwjc0        ),   
    .w93gdpnnxuydy53eu0s9nxw7xdct7       (w93gdpnnxuydy53eu0s9nxw7xdct7      ), 

    .cn8o3075eju6dycby     (cuxedtph_mmf5zt      ), 
    .zi39s8s7rmgo_lyocr_(axp009bfo575n9sjnnf ), 
    .g1cek93tezrlyyt    (brl3pfi8fhhizf3u     ), 
    .i22z6k7eo0it77lz2     (zcfxekf7ptrviima      ), 
    .ldj4m511gvpu12mdu1_ (f29yand0_mv30jc6grvj6  ), 
    .sl5f3k5g9ln8_zvzr  (uys2_c7rmnm5gjf6t   ), 
    .w2h8uh3l463qbgqmv       (umnrzb6pv8dzc        ), 


    .af5qc04tmn51e4u2h1z    (af5qc04tmn51e4u2h1z),
    .ciw6wwc7i33adp5         (chezfp7x0va2ea9tdq),
    .elspwgn4qhqqwg31epb      (elspwgn4qhqqwg31epb),
    .phk590vi2           (phk590vi2       ),
    .rnx27onf2lbe          (rnx27onf2lbe), 
    .ya8t4ev_aidf0t0x4or    (ya8t4ev_aidf0t0x4or),
    .rb050tnl             (rb050tnl),
    .e1go3iu             (e1go3iu),
    .el7_p8jit09           (el7_p8jit09),
    .a94vd35etec4           (a94vd35etec4),
    .l9erxxpnphqd26vg9        (l9erxxpnphqd26vg9),
    .vf5xcr67bqhzlo43_        (vf5xcr67bqhzlo43_),

    .vmx1fh4kmh4c             (vmx1fh4kmh4c),


    .wtd_nuaeb_mpye           (wtd_nuaeb_mpye    ), 
    .x7eg618xaszd4f21cl_g       (x7eg618xaszd4f21cl_g),


    .elth4vimq_j               (cmt_epc        ),
    .jlud6jeuxe0espga           (jlud6jeuxe0espga    ),




    .xd66pm611ai1dg             (xd66pm611ai1dg      ),
    .r9uxubpl2h2alj1q         (r9uxubpl2h2alj1q  ),
    .ftp0juzjm2b587cyw5       (ftp0juzjm2b587cyw5  ),

    .sf0uuehfhfa              (sf0uuehfhfa       ),
    .hvy2cpsp75f3               (hvy2cpsp75f3        ),
    .k3z202os              (k3z202os       ),
    .z35xlcc6bt4               (z35xlcc6bt4        ),
    .ew08uu2kn2p9e11s           (ew08uu2kn2p9e11s    ),
    .xv08lot3vi9dag4vs0       (xv08lot3vi9dag4vs0),
    .mtc04rctrfyb          (mtc04rctrfyb    ),
    .if5jz8qk0aqefy3v35o      (if5jz8qk0aqefy3v35o),

    .jw4fsjecr0u919fr7  (cmt_dret_ena     ),
    .rrujrlc85mhm  (rrujrlc85mhm     ),



    .r4bs4k_53n5wp         (r4bs4k_53n5wp      ),
    .i7lgezdqu4bmka         (i7lgezdqu4bmka      ),

    .h_qwsgi7nk2           (h_qwsgi7nk2        ),
    .bde41te346q515l            (bde41te346q515l         ),
    .tvh1llq2i3_y            (tvh1llq2i3_y         ),
    .w632tcbtqncn6         (w632tcbtqncn6      ),

    .ai169tbqp4seb3            (ai169tbqp4seb3         ),
    .b0zz_ornhz010            (b0zz_ornhz010         ),
    .yw4o4kdms07_32            (yw4o4kdms07_32         ),
    .ezl3jzeqhltgj7h            (ezl3jzeqhltgj7h         ),
    .w529wbj853            (w529wbj853         ),
    .i9xvsmm45fp0f58            (i9xvsmm45fp0f58         ),

    .u25pqekq4df            (u25pqekq4df         ),
    .dhjwho76fa8hqc        (dhjwho76fa8hqc     ),
    .xel6gw173w5x0           (xel6gw173w5x0        ),
    .icauf4l_12_c2xkj53lf       (icauf4l_12_c2xkj53lf    ),
    .v8ydjtlz16x9tx          (v8ydjtlz16x9tx       ),
    .e_z6d7r9kxqg32te      (e_z6d7r9kxqg32te   ),
    .p5jpgn4rvarpo              (p5jpgn4rvarpo           ),
    .z2g63deibg1b1quqr          (z2g63deibg1b1quqr       ),
    .tlgcdv86voe9          (tlgcdv86voe9       ),
    .u_ufp_wg29ieoklxxz1      (u_ufp_wg29ieoklxxz1   ),
    .s_m3pbf5m2tr6v          (s_m3pbf5m2tr6v       ),

    .bj7h5jqg66r51jxki6emra     (bj7h5jqg66r51jxki6emra  ),
    .zmfo8cca_77pc         (zmfo8cca_77pc      ),

    .miax48k27o484e8a         (miax48k27o484e8a      ),

    .fzdb65fcrotwcaccus_cwo     (fzdb65fcrotwcaccus_cwo  ),
    .tcy_87vt9vet39knuw      (tcy_87vt9vet39knuw   ),
    .fc_4ns_w1nh4h02z_dgg    (fc_4ns_w1nh4h02z_dgg ),

    .d3hccrck1fl7jjf6          (d3hccrck1fl7jjf6       ),

    .vkyge0q4mfc5          (vkyge0q4mfc5       ),
    .cppkd01vpwwnlfy           (cppkd01vpwwnlfy        ),

    .psx330qmvh5so1to4iq     (psx330qmvh5so1to4iq  ),
    .sefocn4wjn2k2f_zvlvnz   (sefocn4wjn2k2f_zvlvnz),  
    .qknomh2kbth19r1osddvzly   (qknomh2kbth19r1osddvzly),  
    .bzz8x0np0dpmdjt1d0w7uf   (bzz8x0np0dpmdjt1d0w7uf),  
    .rl9a96pgy3troiao05jel   (rl9a96pgy3troiao05jel),  
    .hzsp_nydab9ghw59v      (hzsp_nydab9ghw59v   ),  

    .pldoasxyzlvx2    (pldoasxyzlvx2       ),


    .unbt3q05xijb   (unbt3q05xijb     ),
    .hawbmpz6j7pzibqr   (hawbmpz6j7pzibqr),

    .o7hoht1pqz01v7            (o7hoht1pqz01v7),
    .kbv2bs_lxmvu             (kbv2bs_lxmvu ),


    .j0qaxhuqtdi       (j0qaxhuqtdi     ),
    .pbzpk52jinfscit4mm     (pbzpk52jinfscit4mm   ),
    .gwj6ow6qvbhs0tc31     (gwj6ow6qvbhs0tc31   ),
    .iwdkm52x_w4hpak_a2_w  (iwdkm52x_w4hpak_a2_w),
    .mm0ssgy582fv_j       (mm0ssgy582fv_j     ),
    .ir2913p9xpmq_1bvfd1  (ir2913p9xpmq_1bvfd1),
    .bsjo0v5e0t556pph  (bsjo0v5e0t556pph),
    .mwegg_7inaca6povsw(mwegg_7inaca6povsw),
    .wnkp7091zrsevkbl  (wnkp7091zrsevkbl),

    .r21i4by0bu3ks             (r21i4by0bu3ks),

    .zmwq3e9oijvo7d7          (zmwq3e9oijvo7d7),

    .sxvvsxtbhyvt        (sxvvsxtbhyvt      ),


    .pydatzxqqi       (pydatzxqqi       ),


    .cwwkpmk260lrt      (nmi_mode),

    .aw82i964do        (aw82i964do),
    .rvr30vvllni    (rvr30vvllni),
    .z1cj655u31    (z1cj655u31),
    .y8_gkxsfle        (y8_gkxsfle),
    .lhu2z948o3n    (lhu2z948o3n),

    .v09gw6e6rfjf05qg  (v09gw6e6rfjf05qg),

    .s5f_36xvqrtq7  (status_mie_r),

    .x6eltyshbu5            (x6eltyshbu5        ),
    .lt3v_fm0ipu            (lt3v_fm0ipu        ),
    .v3ne7glf8d8            (v3ne7glf8d8        ),
    .v9dnbgjy6c0vf          (v9dnbgjy6c0vf      ),
    .hmzw4exmjn8k921c           (hmzw4exmjn8k921c       ),

    .siifnhwgancn8            (siifnhwgancn8        ),
    .mfzl2fqml69hx            (mfzl2fqml69hx        ),
    .aw0hbwfkx3f63s            (aw0hbwfkx3f63s        ),
    .u83p4flbuvkqt26z          (u83p4flbuvkqt26z      ),
    .tvglhc8o_izdq           (tvglhc8o_izdq       ),

    .ij_sgq3rtvw2               (ij_sgq3rtvw2           ),
    .k9jntnqwqp              (k9jntnqwqp          ),

    .b0ry73kp6sc2 (b0ry73kp6sc2),
    .hr64e6c3gy  (hr64e6c3gy ),
    .cz1hh6af7xp2 (cz1hh6af7xp2),
    .st2zalpx0uf (st2zalpx0uf),          
    .w30ye15yns15 (w30ye15yns15),
    .ni01kj42oob2x (ni01kj42oob2x),          
    .ah8kjlmvnaxzbi (ah8kjlmvnaxzbi),          
    .fkuqlh34r (fkuqlh34r), 
    .hnc10arn_rd (hnc10arn_rd),
    .b2ulqcjb  (b2ulqcjb ),

    .dk2xhkj77a       (dk2xhkj77a      ),
    .gf33atgy           (gf33atgy          ),
    .ru_wi         (ru_wi        ) 
  );

  assign emc_bywzarijbo = (~tw5xnp59d8x) & (
                      (~(vi03qlql8tkd5 & ~b0ylmw5xa8oytsw3j6n)) | jjzotrbn | qo5p9t6s74zxpo 

                    | enwn0u48p2_ls5az80
                    | miax48k27o484e8a
                    | (~refz65mt7g99f_cb9h)
                    | (kvpemhoim1tq5y8mzwvix5)   
                    | (~f29yand0_mv30jc6grvj6)
                    | p7ah58va5_2njbtv  
                      )
                    ;


  assign z1l_kkshyf_56cwmaq2dm = fkuqlh34r;
  assign w7u50np_chxy7wq5n9et_q = hnc10arn_rd;
  assign l2dse4sd3runnrb1rcbydauc  = b2ulqcjb;
  assign kr1rhzlb5gr_wty1pe392s5oqet  = rm1dxjejhq7dh3q5m;
  assign ox2ptuhum_e2aodz8wine6h  = st2zalpx0uf;
  assign g_qmxgznvfin609fmm97kuc2dm02  = ni01kj42oob2x;
  assign i9oln6xm1pi9dzsd61s1kg4dmo7j  = ah8kjlmvnaxzbi;
  assign hei_cs0rbwsv  = w30ye15yns15;
  assign yf_5vs18cke5xg660my  = sxvvsxtbhyvt;
  

  assign uzevp4zrbs9gi = rnx27onf2lbe;





  assign aykpj7s87z_wdrbcx0hx  = f1k1tltm39p_5uxhp5l80q4;


  assign se2buoxmq91dbic3y2m5hu =    f0jwv0n5olimpf4vnvqpb4hs
                                 || dw2ygdedledlm7ps830qgbwonu
                                 ;




























endmodule                                      
























module m5_5v7i1cz62p(



  input                          cxkzjh6fduft16beuemi, 
  output                         uej0jzoacitho9mnzs, 
  input  [64-1:0]        hw1xobm2iv3kaij,
  input  [5-1:0] uwtwaa7c9764reokvm5,
  input                          f12hi8g2fiznovp,
  input                          k7wz0kgj7f94f7hml,
  input                          fkcyj1aq49159mfj,
  input                          i68lo1vqlv0o48k7,   
  input [4-1:0]   pupdpprs2srhv_sg,




  input                           j26xb89a8xae2cmtqfby, 
  output                          mpl24r05br_tctrlxtx8d6p, 
  input  [64-1:0]         k9ahcr_bj7e3lceyvmetj8,
  input  [5-1:0]                  axktcwwx1l7erym3mvldq,
  input  [5-1:0]  qil8zvwqkkfkcj8129d,
  input                           x5ug4xxlpdw8ph_oo7x_m,
  input                           fctsirgaydqowic465q,
  input                           mcnqahf70rz3wm2ilvhef,
  input [4-1:0]       u6gfx2g2h7t88vvhusrs5j,




  input                           owijmnymkyht7li_w68, 
  output                          a3ns4toutens4xm0pf6a, 
  input [4-1:0]       i_2sypygf_zqo5p_t7fy ,

  output                          seccdclbkfl        ,
  output [4-1:0]      g6hr2opjly0       ,
  output                          l9193amyxxm9g        ,
  output [4-1:0]      gehkicmawq02an4       ,
  output                          fcl5ybv5a2t4y        ,
  output [4-1:0]      ukjsioluzl5t       ,



  output                          v1kvt26zg5d2p1i3,
  output  [64-1:0]        z6cksoto8caeb0w8461f,
  output  [5-1:0] v5l563s9x82qkxwsx,

  output                          r7sap4hhn2lpgz_5t1t,
  output  [64-1:0]        safx984k5yjm7fd8b3i,
  output  [5-1:0] pvrou_4d1woq_z6q,

  output                          hvxtf10aywneycg3,
  output  [64-1:0]        qs405gb8afw52z6eyxi,
  output  [5-1:0] e_277pojqob91detq806,

  output                          f71k3zhdtjavw19c52g45,  
  output  vpzy7702dz4cc20ajy,
  output  [64-1:0] nwd_h3lrfk59xijt4s7qh1,
  output  [5-1:0] s0n0jneoy6ez4dfj5y_9eq,
  output  [5-1:0] sta4f_rkbcr520sb707nff,
  output ptyuk4efbbdu9asp0b8cmreeh,  


  output  mt0fxo7jph1jww9bml7,
  output  katolbldvqgqsog94,
  output  z22u8178eey1vl3,  




  input  gf33atgy,
  input  ru_wi
  );







    
    
    assign mpl24r05br_tctrlxtx8d6p = 1'b1;
    assign uej0jzoacitho9mnzs   = f12hi8g2fiznovp ? (i68lo1vqlv0o48k7 & cxkzjh6fduft16beuemi) : 1'b1;
    
    wire   j7ncmxtfohotzfc9  = cxkzjh6fduft16beuemi & uej0jzoacitho9mnzs & f12hi8g2fiznovp & i68lo1vqlv0o48k7;
    assign v1kvt26zg5d2p1i3   =  j7ncmxtfohotzfc9 & (~k7wz0kgj7f94f7hml);
    assign z6cksoto8caeb0w8461f  = hw1xobm2iv3kaij[64-1:0];
    assign v5l563s9x82qkxwsx = uwtwaa7c9764reokvm5;




    assign r7sap4hhn2lpgz_5t1t   = 1'b0;
    assign safx984k5yjm7fd8b3i  = 64'b0;
    assign pvrou_4d1woq_z6q = 5'b0;

    assign hvxtf10aywneycg3    = j26xb89a8xae2cmtqfby & mpl24r05br_tctrlxtx8d6p & (~x5ug4xxlpdw8ph_oo7x_m) & fctsirgaydqowic465q;
    assign qs405gb8afw52z6eyxi   = k9ahcr_bj7e3lceyvmetj8[64-1:0];
    assign e_277pojqob91detq806  = qil8zvwqkkfkcj8129d;

    assign mt0fxo7jph1jww9bml7   = cxkzjh6fduft16beuemi & uej0jzoacitho9mnzs & f12hi8g2fiznovp & fkcyj1aq49159mfj;


    assign katolbldvqgqsog94   = 1'b0;

    assign z22u8178eey1vl3   = j26xb89a8xae2cmtqfby & mpl24r05br_tctrlxtx8d6p & fctsirgaydqowic465q & mcnqahf70rz3wm2ilvhef;

      wire l7jdt7plpa0cj8eyq = cxkzjh6fduft16beuemi & uej0jzoacitho9mnzs & k7wz0kgj7f94f7hml & f12hi8g2fiznovp;
      wire kbf7vccq5wdokidaop1 = j26xb89a8xae2cmtqfby & mpl24r05br_tctrlxtx8d6p & x5ug4xxlpdw8ph_oo7x_m & fctsirgaydqowic465q;


      wire [4:0] vs4ta1kq798ck = l7jdt7plpa0cj8eyq ? 5'b0  : axktcwwx1l7erym3mvldq;
      wire [5-1:0] afgjc4gl7iktp1cf = l7jdt7plpa0cj8eyq ? uwtwaa7c9764reokvm5 : qil8zvwqkkfkcj8129d;
      wire yydetudxf41g = l7jdt7plpa0cj8eyq ? k7wz0kgj7f94f7hml : x5ug4xxlpdw8ph_oo7x_m;
      wire mqbwvne2qsvl1xp   = l7jdt7plpa0cj8eyq ? f12hi8g2fiznovp   : fctsirgaydqowic465q;
      wire [64-1:0] um__n7hbw6b   = l7jdt7plpa0cj8eyq ? hw1xobm2iv3kaij[64-1:0] : k9ahcr_bj7e3lceyvmetj8[64-1:0];

      wire ffn89_zo5701ravt5qz = l7jdt7plpa0cj8eyq | kbf7vccq5wdokidaop1;

      assign vpzy7702dz4cc20ajy    = ffn89_zo5701ravt5qz;
      assign nwd_h3lrfk59xijt4s7qh1   = um__n7hbw6b;
      assign s0n0jneoy6ez4dfj5y_9eq  = vs4ta1kq798ck;
      assign sta4f_rkbcr520sb707nff  = afgjc4gl7iktp1cf;
      assign ptyuk4efbbdu9asp0b8cmreeh =  ffn89_zo5701ravt5qz;

    assign f71k3zhdtjavw19c52g45  = v1kvt26zg5d2p1i3 | r7sap4hhn2lpgz_5t1t | hvxtf10aywneycg3;



  assign seccdclbkfl  = (cxkzjh6fduft16beuemi & uej0jzoacitho9mnzs);
  assign g6hr2opjly0 = pupdpprs2srhv_sg ;


  assign l9193amyxxm9g  = j26xb89a8xae2cmtqfby & mpl24r05br_tctrlxtx8d6p & (~x5ug4xxlpdw8ph_oo7x_m) ;
  assign gehkicmawq02an4 = u6gfx2g2h7t88vvhusrs5j;




  wire fhv19ylanj51_yq;
  wire [4-1:0] p_59ub3fg0fho9hq0pax8;
  ux607_gnrl_dfflr #(1) wixkpmz0j8doaxe6  (1'b1  , owijmnymkyht7li_w68      , fhv19ylanj51_yq      , gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(4) fy8qtapdyp3hhcwxih  (owijmnymkyht7li_w68  , i_2sypygf_zqo5p_t7fy      , p_59ub3fg0fho9hq0pax8      , gf33atgy, ru_wi);
  assign fcl5ybv5a2t4y        = fhv19ylanj51_yq      ;
  assign ukjsioluzl5t       = p_59ub3fg0fho9hq0pax8 ;


  assign a3ns4toutens4xm0pf6a = 1'b1;

endmodule                                      





















module fqo7x_ckpw9266xb2d57x8(



  input                          cxkzjh6fduft16beuemi, 
  output                         uej0jzoacitho9mnzs, 
  input  [5-1:0] uwtwaa7c9764reokvm5,
  input  [64-1:0]        hw1xobm2iv3kaij,
  input                          f12hi8g2fiznovp,
  input                          k7wz0kgj7f94f7hml,
  input                          fkcyj1aq49159mfj,
  input                          i68lo1vqlv0o48k7,   
  input [4-1:0]   pupdpprs2srhv_sg,




  input                           j26xb89a8xae2cmtqfby, 
  output                          mpl24r05br_tctrlxtx8d6p, 
  input  [64-1:0]         k9ahcr_bj7e3lceyvmetj8,
  input  [5-1:0]                  axktcwwx1l7erym3mvldq,
  input  [5-1:0]  qil8zvwqkkfkcj8129d,
  input                           x5ug4xxlpdw8ph_oo7x_m,
  input                           fctsirgaydqowic465q,
  input                           mcnqahf70rz3wm2ilvhef,
  input [4-1:0]       u6gfx2g2h7t88vvhusrs5j,



  input                           owijmnymkyht7li_w68, 
  output                          a3ns4toutens4xm0pf6a, 
  input [4-1:0]       i_2sypygf_zqo5p_t7fy ,

  output                          seccdclbkfl        ,
  output [4-1:0]      g6hr2opjly0       ,
  output                          l9193amyxxm9g        ,
  output [4-1:0]      gehkicmawq02an4       ,
  output                          fcl5ybv5a2t4y        ,
  output [4-1:0]      ukjsioluzl5t       ,



  output                          v1kvt26zg5d2p1i3,
  output  [64-1:0]        z6cksoto8caeb0w8461f,
  output  [5-1:0] v5l563s9x82qkxwsx,

  output                          r7sap4hhn2lpgz_5t1t,
  output  [64-1:0]        safx984k5yjm7fd8b3i,
  output  [5-1:0] pvrou_4d1woq_z6q,

  output                          hvxtf10aywneycg3,
  output  [64-1:0]        qs405gb8afw52z6eyxi,
  output  [5-1:0] e_277pojqob91detq806,

  output                          f71k3zhdtjavw19c52g45,  
  output  vpzy7702dz4cc20ajy,
  output  [64-1:0] nwd_h3lrfk59xijt4s7qh1,
  output  [5-1:0] s0n0jneoy6ez4dfj5y_9eq,
  output  [5-1:0] sta4f_rkbcr520sb707nff,
  output ptyuk4efbbdu9asp0b8cmreeh,  


  output  mt0fxo7jph1jww9bml7,
  output  katolbldvqgqsog94,
  output  z22u8178eey1vl3,  

  output                          uy7dkgcktef73e762sbkgdq2teb, 
  output  [4 -1:0] wsnaf53u3elqrc9oym2gh69u5 ,
  output  [64 -1:0]       e49tm9dpy3o9o2w9ac5yowmx ,

  input  gf33atgy,
  input  ru_wi
  );
  wire                         h1qsftcbdojcb1s5en;
  wire                         o68w5q05bpjtka;
  wire                         tnqagwcmpxu0c  ;
  wire [64 -1:0]       grqmvi5e4v7fp ;
  wire [4 -1:0] mcs6931j0dy0tx ;

  assign uy7dkgcktef73e762sbkgdq2teb   = h1qsftcbdojcb1s5en;
  assign wsnaf53u3elqrc9oym2gh69u5    = mcs6931j0dy0tx ;
  assign e49tm9dpy3o9o2w9ac5yowmx    = grqmvi5e4v7fp ;



  localparam aafrtcd422sh = 1+64+4;



  wire [aafrtcd422sh-1:0] uhh5eeau4yulwu7 = {
                                          f12hi8g2fiznovp,
                                          hw1xobm2iv3kaij,
                                          pupdpprs2srhv_sg   
                                        };   
  wire [aafrtcd422sh-1:0] tvaqurc_gjqpnyqr; 
  ux607_gnrl_bypbuf # (
    .DP(1),
    .DW(aafrtcd422sh) 
  ) kmbgh2n3oqe7wck0d8hj(
      .i_vld   (cxkzjh6fduft16beuemi),
      .i_rdy   (uej0jzoacitho9mnzs),

      .o_vld   (h1qsftcbdojcb1s5en),
      .o_rdy   (o68w5q05bpjtka),

      .i_dat   (uhh5eeau4yulwu7),
      .o_dat   (tvaqurc_gjqpnyqr),

      .clk     (gf33atgy  ),
      .rst_n   (ru_wi)
  );
  assign { 
           tnqagwcmpxu0c,
           grqmvi5e4v7fp,
           mcs6931j0dy0tx   
         } = tvaqurc_gjqpnyqr;




  m5_5v7i1cz62p bx3md36rhpuhyflzadfh(
    .mt0fxo7jph1jww9bml7   (mt0fxo7jph1jww9bml7),
    .katolbldvqgqsog94   (katolbldvqgqsog94),
    .z22u8178eey1vl3   (z22u8178eey1vl3),

    .cxkzjh6fduft16beuemi   (h1qsftcbdojcb1s5en   ), 
    .uej0jzoacitho9mnzs   (o68w5q05bpjtka   ),
    .hw1xobm2iv3kaij    (grqmvi5e4v7fp    ),
    .pupdpprs2srhv_sg    (mcs6931j0dy0tx    ),  
    .f12hi8g2fiznovp     (tnqagwcmpxu0c     ), 
    .i68lo1vqlv0o48k7     (i68lo1vqlv0o48k7   ), 
    .uwtwaa7c9764reokvm5   (uwtwaa7c9764reokvm5 ),
    .k7wz0kgj7f94f7hml   (k7wz0kgj7f94f7hml ), 
    .fkcyj1aq49159mfj    (1'b0   ), 

    .j26xb89a8xae2cmtqfby (j26xb89a8xae2cmtqfby),  
    .mpl24r05br_tctrlxtx8d6p (mpl24r05br_tctrlxtx8d6p),  
    .k9ahcr_bj7e3lceyvmetj8  (k9ahcr_bj7e3lceyvmetj8 ),  
    .qil8zvwqkkfkcj8129d (qil8zvwqkkfkcj8129d),  
    .x5ug4xxlpdw8ph_oo7x_m (x5ug4xxlpdw8ph_oo7x_m),  
    .axktcwwx1l7erym3mvldq (axktcwwx1l7erym3mvldq),  
    .fctsirgaydqowic465q   (fctsirgaydqowic465q  ),  
    .u6gfx2g2h7t88vvhusrs5j  (u6gfx2g2h7t88vvhusrs5j ),  

    .mcnqahf70rz3wm2ilvhef  (1'b0   ), 



    .v1kvt26zg5d2p1i3      (v1kvt26zg5d2p1i3   ),
    .z6cksoto8caeb0w8461f     (z6cksoto8caeb0w8461f  ),
    .v5l563s9x82qkxwsx    (v5l563s9x82qkxwsx ),

    .r7sap4hhn2lpgz_5t1t      (r7sap4hhn2lpgz_5t1t    ),
    .safx984k5yjm7fd8b3i     (safx984k5yjm7fd8b3i    ),
    .pvrou_4d1woq_z6q    (pvrou_4d1woq_z6q   ),

    .hvxtf10aywneycg3      (hvxtf10aywneycg3    ),
    .qs405gb8afw52z6eyxi     (qs405gb8afw52z6eyxi    ),
    .e_277pojqob91detq806    (e_277pojqob91detq806   ),

    .owijmnymkyht7li_w68  (owijmnymkyht7li_w68), 
    .a3ns4toutens4xm0pf6a  (a3ns4toutens4xm0pf6a), 
    .i_2sypygf_zqo5p_t7fy   (i_2sypygf_zqo5p_t7fy ),

    .seccdclbkfl          (seccdclbkfl      ),
    .g6hr2opjly0         (g6hr2opjly0     ),
    .l9193amyxxm9g          (l9193amyxxm9g      ),
    .gehkicmawq02an4         (gehkicmawq02an4     ),
    .fcl5ybv5a2t4y          (fcl5ybv5a2t4y      ),
    .ukjsioluzl5t         (ukjsioluzl5t     ),



    .vpzy7702dz4cc20ajy      (vpzy7702dz4cc20ajy    ),
    .nwd_h3lrfk59xijt4s7qh1     (nwd_h3lrfk59xijt4s7qh1   ),
    .s0n0jneoy6ez4dfj5y_9eq    (s0n0jneoy6ez4dfj5y_9eq  ),
    .sta4f_rkbcr520sb707nff    (sta4f_rkbcr520sb707nff  ),
    .ptyuk4efbbdu9asp0b8cmreeh   (ptyuk4efbbdu9asp0b8cmreeh ),
    .f71k3zhdtjavw19c52g45       (f71k3zhdtjavw19c52g45),


    .gf33atgy                 (gf33atgy          ),
    .ru_wi               (ru_wi        ) 
  );


endmodule




















module hprqrck8t9y3rksec (
  input lodtxdqjnwvx, 
  input cbbcxlflqkqoklckuekt, 
  input n37wgp2u95gc5b_, 
  input ewe_b1wv9zhrc8rc6hhr, 
  input z28w9as50xav1c2ms, 

  
  
  
  

  
  input                   s6ypv533tdywrez9dra,
  input                   wtxn5hz27d1ke0cp5p,
  input                   z_g_9tmwi_9phwpm,
  input [12-1:0]          zy04ur_r6ibez7,
  input  [64-1:0] tpenqez_048wjs0mji00,
  output [64-1:0] wg_nk5anc77k66ap,

  output                  m9i5nb3fpl7i1c2f7aqnda5a,
  output                  o9n8q26y9zbsj6n3w7zzdgn_d7n90v,
  output                  fc8jy9eix4zbo26a2l3mebjykj99y,
  
  output                  zds0n3s_2vya92r6p0iu18ede83st,
  output                  j_oxbujpaq4zahlaf42l9paa_kjbrj,
  

  
  
  output                             x8rpm78rvvycis, 
  input                              bwbmafs1inesgjyn, 
  input                              bkkiffh6ob85nh79doya_, 
  input  [5:0]                       qhqqh0lyehgtfop1tc, 
  output [74-1:0] canacnkc7zibtkn418i, 

  output                             sxhicsqvufwfbnk0, 
  input                              ydydp69z03wvr97, 
  input                              pjic5x84bqxpvdduy4r2s, 
  input                              w5az87bw32r0tjbo0tdrv2ouvx, 
  output [74-1:0] x03ux1utw4qem5kk3c, 

  
  
  output                             vs6ryzcr0bwqs5so, 
  output [32-1:0]            j25ub196dc_agl8oovaex4, 
  output                             pi2nokcm8qf7och7l4g, 
  output                             c0i0hs5tz64_ce5f0z, 
  output                             dmzdczrqcueolg3dzufj_by5rmf, 
  output                             a1sqko6fok9qzpbtyuw0, 
  output                             bquohubxiv2rsayn62v, 
  input                              kqyojh1maxy0x834htg, 


  
  

  input                                    fkuqlh34r,                  
  input                                    ni01kj42oob2x,                  
  input                                    ah8kjlmvnaxzbi,                  
  input  [1:0]                             st2zalpx0uf,                  
  input                                    rm1dxjejhq7dh3q5m,                  
  input                                    sxvvsxtbhyvt,                  

  
  output                                   hpk3eafyque5ubt_c62flnny,        
  output [27-1:0]      sfezv1xz2ghvo8pkt,               
  output [1:0]                             vagaza053272juvmo59v8w20s,        
  output                                   rzf45534z36ejq96260,                        
  output [26-1:0]    frzfsbt7hp3n4aj3zvvumnh0s,         
  output [64-1:0]                  zkuxqezrmlhyyjjgx,              
  output [64-1:0]                  u3h5tvu1g2q93141j9o,              
  output                                   pjh0wad7t_5du3cync_0c,                        
  
  output                                   wmkgrgf631pbq,
  input                                    oyq1p3qa2iffjuqns0jkgg,

  
  input                                    qjw2q0j88rjr42lautsqnca,        
  input [26-1:0]     imkm56ujne9v4m6n08w1yf5622,     
  input [20-1:0]          txk1r9aiq_7l2nkw101w_,          
  input                                    ih4hmwugasiodbx5da9_40kx,         
  input                                    x5vjq7mshfwr0h3q514t7mhdt,         
  input                                    qrxtk7e03100_uwkx73sg7,         
  input                                    i7qiq2q9c6hbeful9qu9lb,         
  input                                    yr0s3skqk7cdqflsrbsxg9znu,         
  input                                    adqieke11qo0elfz93hlouwjc0,   
  input                                    w93gdpnnxuydy53eu0s9nxw7xdct7, 

  
  
  
  output                             cn8o3075eju6dycby,  
  output                             zi39s8s7rmgo_lyocr_, 
  output [5-1:0]  g1cek93tezrlyyt, 
  output [64-1:0]            i22z6k7eo0it77lz2, 
  
  output                             ldj4m511gvpu12mdu1_,           
  output                             sl5f3k5g9ln8_zvzr,            
  input                              w2h8uh3l463qbgqmv,



  input  gf33atgy,
  input  ru_wi

  );

  wire aw82i964do = lodtxdqjnwvx;
  wire pydatzxqqi = z28w9as50xav1c2ms;
  wire y8_gkxsfle = n37wgp2u95gc5b_ & ~pydatzxqqi;
  wire s36z1abpqp = ~aw82i964do & ~pydatzxqqi & ~y8_gkxsfle;

  wire nyj60jhovrm8ck221y      = (zy04ur_r6ibez7 == 12'h7cb);
  wire wbpgavgnkjjioa8e3u9jm        = (zy04ur_r6ibez7 == 12'h7cc);
  wire xwz38wal3a2otarp2q2vo1pc;
  wire r97lptnbuajdq           = (zy04ur_r6ibez7 == 12'h7cd);
  wire ykmql1hqw3n46ozed            = (zy04ur_r6ibez7 == 12'h7ce);
  wire xsr2q02ms3e_kgdajc      = (zy04ur_r6ibez7 == 12'h5cb);
  wire idj84m6wh4hfma_4ko        = (zy04ur_r6ibez7 == 12'h5cc);
  wire zckng96c3vahiptf5xbt;
  wire zx9t7k1djh2xjrdy1i           = (zy04ur_r6ibez7 == 12'h5cd);
  wire vms1aagsjxnv;            
  wire p2s3rf_4d5qsvgov3eid_zq      = (zy04ur_r6ibez7 == 12'h4cb);
  wire vbla5rqpxkbflrtm        = (zy04ur_r6ibez7 == 12'h4cc);
  wire y2wqtcjri2rtyk60djlh;
  wire wbr64ehh7_1bx           = (zy04ur_r6ibez7 == 12'h4cd);
    
  wire hz3z0shjzrq3zuflmge      = nyj60jhovrm8ck221y      & z_g_9tmwi_9phwpm;
  wire hwwmcp9n_lron4dyadi        = wbpgavgnkjjioa8e3u9jm        & z_g_9tmwi_9phwpm;
  wire jm3juv14fels           = r97lptnbuajdq           & z_g_9tmwi_9phwpm;
  wire j5eu9hpjatwy6347            = ykmql1hqw3n46ozed            & z_g_9tmwi_9phwpm;
  wire n00xak5ss49lfu8hojy      = xsr2q02ms3e_kgdajc      & z_g_9tmwi_9phwpm;
  wire m6wvsbta6h7uz9w        = idj84m6wh4hfma_4ko        & z_g_9tmwi_9phwpm;
  wire iiqf_1ral3nh9o           = zx9t7k1djh2xjrdy1i           & z_g_9tmwi_9phwpm;
  wire lal8o4x20d5059pi0k7z      = p2s3rf_4d5qsvgov3eid_zq      & z_g_9tmwi_9phwpm;
  wire ubtmpc65a9oq6qvwghu1        = vbla5rqpxkbflrtm        & z_g_9tmwi_9phwpm;
  wire snfhp659sfq2           = wbr64ehh7_1bx           & z_g_9tmwi_9phwpm;
    
  wire vtuhwpwy1u_h059d2f      = nyj60jhovrm8ck221y      & wtxn5hz27d1ke0cp5p & s6ypv533tdywrez9dra;
  
  
  
  
  
  
  wire abniijg5zst5pbmx4q        = wbpgavgnkjjioa8e3u9jm        & wtxn5hz27d1ke0cp5p & s6ypv533tdywrez9dra;
  wire qi7ljmpbj6_hp_           = r97lptnbuajdq           & wtxn5hz27d1ke0cp5p & s6ypv533tdywrez9dra;
  wire yyxw_dgmuxg34z            = ykmql1hqw3n46ozed            & wtxn5hz27d1ke0cp5p & s6ypv533tdywrez9dra;
  wire ganxldhqmi26thelvrc5      = xsr2q02ms3e_kgdajc      & wtxn5hz27d1ke0cp5p & s6ypv533tdywrez9dra;
  
  
  
  
  
  
  wire szntcqan754qrdh        = idj84m6wh4hfma_4ko        & wtxn5hz27d1ke0cp5p & s6ypv533tdywrez9dra;
  wire evd4lbrrfrlt           = zx9t7k1djh2xjrdy1i           & wtxn5hz27d1ke0cp5p & s6ypv533tdywrez9dra;
  wire pqghoaaf_0uy5o7vmmvd6d      = p2s3rf_4d5qsvgov3eid_zq      & wtxn5hz27d1ke0cp5p & s6ypv533tdywrez9dra;
  
  
  
  
  
  
  wire cll6ubptbwvtxo0lc        = vbla5rqpxkbflrtm        & wtxn5hz27d1ke0cp5p & s6ypv533tdywrez9dra;
  wire kqn3xki834s2uls           = wbr64ehh7_1bx           & wtxn5hz27d1ke0cp5p & s6ypv533tdywrez9dra;

  
  wire uv8iclz1yq8 = 1'b1;

  wire [64-1:0] k2zur8td8o4265j5k1;
  wire [64-1:0] i6yyrngwp25i53cqkim9;
  wire [64-1:0] tzxdf39sspr1_q0sfb;
  
  wire                 p2smibeuelrp8hsca6vc8w6q;
  wire                 kidn1h9_lj8wzplj4kd32;
  wire                 gr5iv52qlkdgsjcutlh5ae;
  wire [64-1:0] b7kat6xkt_rgc2hdogj3k =   ({64{p2smibeuelrp8hsca6vc8w6q}} & k2zur8td8o4265j5k1)
                                                 | ({64{gr5iv52qlkdgsjcutlh5ae}} & i6yyrngwp25i53cqkim9)
                                                 | ({64{kidn1h9_lj8wzplj4kd32}} & tzxdf39sspr1_q0sfb)
                                                 ;
  wire [64-1:0] tqv0jti68ruy0moh = b7kat6xkt_rgc2hdogj3k + (1<<5); 

  wire batr98hpda = x8rpm78rvvycis | sxhicsqvufwfbnk0;
  wire x5bkt27dkr_7 = bwbmafs1inesgjyn | ydydp69z03wvr97;
  wire xjrmfp3ofdru4pyfjw = bkkiffh6ob85nh79doya_ | pjic5x84bqxpvdduy4r2s;
  wire [3-1:0] td1nncrrbp273gpbj6cq;
  wire en1q7v03lnxlj7aw4dpakyg0;
  wire igimbt9i77_wg1s8b6;

  
  
   wire fdc8111sh6h232;

   wire xbia17vq5zswh4 = fdc8111sh6h232 & igimbt9i77_wg1s8b6 & p2smibeuelrp8hsca6vc8w6q;
   wire oswe4ru1tv0 = xbia17vq5zswh4 ;
   wire bomw_wos9tnq5p5oe4q7sh = uv8iclz1yq8  & (vtuhwpwy1u_h059d2f | oswe4ru1tv0);
   wire [64-1:0] wepgerwk8uekz56dukn = ({64{vtuhwpwy1u_h059d2f}} & tpenqez_048wjs0mji00[64-1:0])
                                                 | ({64{oswe4ru1tv0}} & tqv0jti68ruy0moh[64-1:0])
                                                 ;
  ux607_gnrl_dfflr #(64) lpdc8omkmdjv_p9mk9kedg9l (bomw_wos9tnq5p5oe4q7sh, wepgerwk8uekz56dukn, k2zur8td8o4265j5k1, gf33atgy, ru_wi);
  wire [64-1:0] acpehvvxyfly37b3c4 = k2zur8td8o4265j5k1;

  
  
  wire ef3mzj71z281qrhxkun = uv8iclz1yq8 & abniijg5zst5pbmx4q;
  wire [64-1:0] pxj0thyzt9xckb7jppl;
  wire [64-1:0] kgdfan3om9krz_2smrw = {{64-5{1'b0}},tpenqez_048wjs0mji00[4:0]};
  ux607_gnrl_dfflr #(64) xvoqjidn177hhk5dyxmqino (ef3mzj71z281qrhxkun, kgdfan3om9krz_2smrw, pxj0thyzt9xckb7jppl, gf33atgy, ru_wi);
  wire [64-1:0]  tpj5e_qxsx38fs13tz = pxj0thyzt9xckb7jppl;
  
  ux607_gnrl_dffr #(1) iga_m000cl0v1v2pc0w0b9ilrgk2 (wbpgavgnkjjioa8e3u9jm, xwz38wal3a2otarp2q2vo1pc, gf33atgy, ru_wi);

  
  
  wire owhsxmah_o1vvv; 
  wire v9e1mwv5cah8h3od8jj = (owhsxmah_o1vvv & en1q7v03lnxlj7aw4dpakyg0 & p2smibeuelrp8hsca6vc8w6q); 
  wire h339d11vb2g9mh8 = uv8iclz1yq8 & (qi7ljmpbj6_hp_ | v9e1mwv5cah8h3od8jj);
  wire [64-1:0] fo1ut1do_1s86qf5;
  wire [64-1:0] b_5z6kaetv_3t7 = ({64{qi7ljmpbj6_hp_}} & {{64-3{1'b0}},tpenqez_048wjs0mji00[3-1:0]})
                                      | ({{64-3{1'b0}},td1nncrrbp273gpbj6cq})  
                                      ;
  ux607_gnrl_dfflr #(64) dnzs3g5ycutfv1yhi_ (h339d11vb2g9mh8, b_5z6kaetv_3t7, fo1ut1do_1s86qf5, gf33atgy, ru_wi);
  wire [64-1:0]  ks5lhl6mm0f68vt6 = fo1ut1do_1s86qf5;

  
  
  wire otgnrw7onbihzy1 = uv8iclz1yq8 & yyxw_dgmuxg34z;
  wire [64-1:0] ydw7u0ctnbhr;
  wire [64-1:0] iednlto8u4l3 = ({64{yyxw_dgmuxg34z}} & {{64-1{1'b0}},tpenqez_048wjs0mji00[0]});

  ux607_gnrl_dfflr #(64) k95fo1ww14sumuji (otgnrw7onbihzy1, iednlto8u4l3, ydw7u0ctnbhr, gf33atgy, ru_wi);
  wire [64-1:0]  xvvnu00tutw2 = ydw7u0ctnbhr;
  assign vms1aagsjxnv = xvvnu00tutw2[0];

  
  

   wire vvwgviupu768t6 = fdc8111sh6h232 & igimbt9i77_wg1s8b6 & kidn1h9_lj8wzplj4kd32;
   wire qvttcf3sbu8fo0hj= vvwgviupu768t6 ;
   wire toaxnsm8_p7pf1z7x8 = uv8iclz1yq8  & (ganxldhqmi26thelvrc5 | qvttcf3sbu8fo0hj);
   wire [64-1:0] l2fmsgojt52_zbzwhtb = ({64{ganxldhqmi26thelvrc5}} & tpenqez_048wjs0mji00[64-1:0])
                                                 | ({64{qvttcf3sbu8fo0hj}} & tqv0jti68ruy0moh[64-1:0])
                                                 ;
  ux607_gnrl_dfflr #(64) a9wsf_0mj6r5lwiw94rpz2 (toaxnsm8_p7pf1z7x8, l2fmsgojt52_zbzwhtb, tzxdf39sspr1_q0sfb, gf33atgy, ru_wi);
  wire [64-1:0] gs404nvjckm3gkxt3k = tzxdf39sspr1_q0sfb;

  
  
  wire qvrzkfitjxh5vkq6 = uv8iclz1yq8 & szntcqan754qrdh;
  wire [64-1:0] h7he7il3sxskkvpyg;
  wire [64-1:0] sp8oq_omzj3qe7myv5m = {{64-5{1'b0}},tpenqez_048wjs0mji00[4:0]};
  ux607_gnrl_dfflr #(64) p9awqcjda4yn7pwjgm5g41 (qvrzkfitjxh5vkq6, sp8oq_omzj3qe7myv5m, h7he7il3sxskkvpyg, gf33atgy, ru_wi);
  wire [64-1:0]  b0asn01va6mrjxk0 = h7he7il3sxskkvpyg;
  
  ux607_gnrl_dffr #(1) y3xyw__ailvs23ndm9ime07ziqstnd (idj84m6wh4hfma_4ko, zckng96c3vahiptf5xbt, gf33atgy, ru_wi);

  
  
  wire f0_6sq9mpnatn6gr8 = (owhsxmah_o1vvv & en1q7v03lnxlj7aw4dpakyg0 & kidn1h9_lj8wzplj4kd32); 
  wire xsz5__8terkg65pdx = uv8iclz1yq8 & (evd4lbrrfrlt | f0_6sq9mpnatn6gr8);
  wire [64-1:0] qdusaaydan1;
  wire [64-1:0] c46rl_wkzo4bkfw = ({64{evd4lbrrfrlt}} & {{64-3{1'b0}},tpenqez_048wjs0mji00[3-1:0]})
                                      | ({{64-3{1'b0}},td1nncrrbp273gpbj6cq})  
                                      ;
  ux607_gnrl_dfflr #(64) ta8bn3qughrs5wg (xsz5__8terkg65pdx, c46rl_wkzo4bkfw, qdusaaydan1, gf33atgy, ru_wi);
  wire [64-1:0]  sfv_3s9pduczih0od_ = qdusaaydan1;

  
  

   wire jv18ebc_1qg = fdc8111sh6h232 & igimbt9i77_wg1s8b6 & gr5iv52qlkdgsjcutlh5ae;
   wire l4lfyk6dj6lr= jv18ebc_1qg ;
   wire ud3q24jy214q9xltxw = uv8iclz1yq8  & (pqghoaaf_0uy5o7vmmvd6d | l4lfyk6dj6lr);
   wire [64-1:0] bw2e4nehpwf1v68h6hx = ({64{pqghoaaf_0uy5o7vmmvd6d}} & tpenqez_048wjs0mji00[64-1:0])
                                                 | ({64{l4lfyk6dj6lr}} & tqv0jti68ruy0moh[64-1:0])
                                                 ;
  ux607_gnrl_dfflr #(64) jbtw2gspe3g22ydnkg2ymjj (ud3q24jy214q9xltxw, bw2e4nehpwf1v68h6hx, i6yyrngwp25i53cqkim9, gf33atgy, ru_wi);
  wire [64-1:0] p_kkuyzrt1jtpp3remf1p0 = i6yyrngwp25i53cqkim9;

  
  
  wire q3rqwxg4lpne86conydxb = uv8iclz1yq8 & cll6ubptbwvtxo0lc;
  wire [64-1:0] gy6l0tq0aapmht624q;
  wire [64-1:0] uposvqc0t2qfvyn7 = {{64-5{1'b0}},tpenqez_048wjs0mji00[4:0]};
  ux607_gnrl_dfflr #(64) hkf4thaqgtfukfswpmuz (q3rqwxg4lpne86conydxb, uposvqc0t2qfvyn7, gy6l0tq0aapmht624q, gf33atgy, ru_wi);
  wire [64-1:0]  b7jun2_699m09sjv2m = gy6l0tq0aapmht624q;
  
  ux607_gnrl_dffr #(1) t3dtoseco_6tapxxzybg90thct (vbla5rqpxkbflrtm, y2wqtcjri2rtyk60djlh, gf33atgy, ru_wi);

  
  
  wire q32kv7agk03dyx3t5qtv9 = (owhsxmah_o1vvv & en1q7v03lnxlj7aw4dpakyg0 & gr5iv52qlkdgsjcutlh5ae); 
  wire c5i0c9a2petotk2vo = uv8iclz1yq8 & (kqn3xki834s2uls | q32kv7agk03dyx3t5qtv9);
  wire [64-1:0] uge5i5dpo9wpp;
  wire [64-1:0] ipbv5fdjko9xcwi21 = ({64{kqn3xki834s2uls}} & {{64-3{1'b0}},tpenqez_048wjs0mji00[3-1:0]})
                                      | ({{64-3{1'b0}},td1nncrrbp273gpbj6cq})  
                                      ;
  ux607_gnrl_dfflr #(64) i0afb1d868m6rtn8 (c5i0c9a2petotk2vo, ipbv5fdjko9xcwi21, uge5i5dpo9wpp, gf33atgy, ru_wi);
  wire [64-1:0]  yxt_oznssyj11tc = uge5i5dpo9wpp;


  
  
  assign {m9i5nb3fpl7i1c2f7aqnda5a, wg_nk5anc77k66ap} = {1'b0,64'b0} 
                 | {nyj60jhovrm8ck221y, ({64{hz3z0shjzrq3zuflmge}} & acpehvvxyfly37b3c4)}
                 | {wbpgavgnkjjioa8e3u9jm  , ({64{hwwmcp9n_lron4dyadi  }} & tpj5e_qxsx38fs13tz  )}
                 | {r97lptnbuajdq     , ({64{jm3juv14fels     }} & ks5lhl6mm0f68vt6     )}
                 | {ykmql1hqw3n46ozed      , ({64{j5eu9hpjatwy6347      }} & xvvnu00tutw2      )}
                 | {p2s3rf_4d5qsvgov3eid_zq, ({64{lal8o4x20d5059pi0k7z}} & p_kkuyzrt1jtpp3remf1p0)}
                 | {vbla5rqpxkbflrtm  , ({64{ubtmpc65a9oq6qvwghu1  }} & b7jun2_699m09sjv2m  )}
                 | {wbr64ehh7_1bx     , ({64{snfhp659sfq2     }} & yxt_oznssyj11tc     )}
                 | {xsr2q02ms3e_kgdajc, ({64{n00xak5ss49lfu8hojy}} & gs404nvjckm3gkxt3k)}
                 | {idj84m6wh4hfma_4ko  , ({64{m6wvsbta6h7uz9w  }} & b0asn01va6mrjxk0  )}
                 | {zx9t7k1djh2xjrdy1i     , ({64{iiqf_1ral3nh9o     }} & sfv_3s9pduczih0od_     )}
              ;

  assign o9n8q26y9zbsj6n3w7zzdgn_d7n90v = 
                 | p2s3rf_4d5qsvgov3eid_zq
                 | vbla5rqpxkbflrtm  
                 | wbr64ehh7_1bx     
                 ;

  assign fc8jy9eix4zbo26a2l3mebjykj99y = s36z1abpqp &  
               (
                 | (~vms1aagsjxnv & p2s3rf_4d5qsvgov3eid_zq)
                 | (~vms1aagsjxnv & vbla5rqpxkbflrtm  ) 
                 | (~vms1aagsjxnv & wbr64ehh7_1bx     )   
               )
                 ;


  assign zds0n3s_2vya92r6p0iu18ede83st = 
                 | xsr2q02ms3e_kgdajc
                 | idj84m6wh4hfma_4ko  
                 | zx9t7k1djh2xjrdy1i     
                 | p2s3rf_4d5qsvgov3eid_zq
                 | vbla5rqpxkbflrtm  
                 | wbr64ehh7_1bx     
                 ;

  assign j_oxbujpaq4zahlaf42l9paa_kjbrj = y8_gkxsfle &  
               (
                 | (~vms1aagsjxnv & xsr2q02ms3e_kgdajc)
                 | (~vms1aagsjxnv & idj84m6wh4hfma_4ko  ) 
                 | (~vms1aagsjxnv & zx9t7k1djh2xjrdy1i     )   
                 | (~vms1aagsjxnv & p2s3rf_4d5qsvgov3eid_zq)
                 | (~vms1aagsjxnv & vbla5rqpxkbflrtm  ) 
                 | (~vms1aagsjxnv & wbr64ehh7_1bx     )   
               )
                 ;


  
  
  wire [64-1:0]mj62ywr =   ({64{p2smibeuelrp8hsca6vc8w6q}} & tpj5e_qxsx38fs13tz)
                                 | ({64{kidn1h9_lj8wzplj4kd32}} & b0asn01va6mrjxk0)
                                 | ({64{gr5iv52qlkdgsjcutlh5ae}} & b7jun2_699m09sjv2m)
                                 ;
  
  wire [64-1:0]xgg3cweyrd0uj_9ekh = b7kat6xkt_rgc2hdogj3k; 

  wire pu7da028_tz7r = (mj62ywr[2:0] == 3'b000);
  wire xnsc6qdckok83v0y = (mj62ywr[2:0] == 3'b001);
  wire em88l_e2n0l = (mj62ywr[2:0] == 3'b010);
  wire oogo4cx3q8tv9mbo = (mj62ywr[2:0] == 3'b011);
  wire fpop_x33d6ai = (mj62ywr[2:0] == 3'b100);
  wire h9ohvklruyeg = (mj62ywr[2:0] == 3'b101);
  wire abh4vum0nod88rk7 = (mj62ywr[2:0] == 3'b110);
  wire ibnxpm9kzoqm5y = (mj62ywr[2:0] == 3'b111);

  wire n6hzwnw9zs  = (mj62ywr[4:3] == 2'b00);
  wire mftzpw3hqrbum  = (mj62ywr[4:3] == 2'b01);
  wire h_zklq46k29uk3  = (mj62ywr[4:3] == 2'b10);
  wire d5yz35iuocu  = (mj62ywr[4:3] == 2'b11);
  
  
  wire rrki1m97jmtyk2r;
  wire i1g4vxhyij_qk9u;
  wire zij1fmhqno571ee5 = ~rrki1m97jmtyk2r
                        & ~i1g4vxhyij_qk9u
                        ;
  wire x3pdmlbidudtcfe    = n6hzwnw9zs & pu7da028_tz7r;
  wire y_lhuhvde       = n6hzwnw9zs & xnsc6qdckok83v0y;
  wire knep835je_uzqghqf  = n6hzwnw9zs & em88l_e2n0l; 
  wire md9w_qvcupymt5     = n6hzwnw9zs & oogo4cx3q8tv9mbo;
  wire pdje7bg4uudiwmaizj   = n6hzwnw9zs & fpop_x33d6ai;
  wire t__jcg4w9op      = n6hzwnw9zs & ibnxpm9kzoqm5y;
  wire ufj54jrgxdnsw4v_   = h_zklq46k29uk3 & ibnxpm9kzoqm5y & (rrki1m97jmtyk2r | i1g4vxhyij_qk9u);
  wire v64tquaebtsdj1cgmtr = (n6hzwnw9zs & abh4vum0nod88rk7)
                       | (h_zklq46k29uk3 & ibnxpm9kzoqm5y & zij1fmhqno571ee5) 
                       ; 
                                                    
  
  wire a601v24iimk0q23vf;
  wire hmtyprargqxng = a601v24iimk0q23vf;
  wire v8lyodmb_xbnrq1r5f5vib_1;
  wire tvr8zxsmimyd3j7y4;
  wire wkpz9dk71bcfhgjwdb1b;

  wire [74-1:0] wfa5o72ctktgt55fgv2eo;
  assign wfa5o72ctktgt55fgv2eo[5  ] = tvr8zxsmimyd3j7y4;  
  assign wfa5o72ctktgt55fgv2eo[6  ] = rrki1m97jmtyk2r;  
  assign wfa5o72ctktgt55fgv2eo[8  ] = v8lyodmb_xbnrq1r5f5vib_1;  
  assign wfa5o72ctktgt55fgv2eo[7  ] = i1g4vxhyij_qk9u;  
  assign wfa5o72ctktgt55fgv2eo[9  ] = wkpz9dk71bcfhgjwdb1b;  
  assign wfa5o72ctktgt55fgv2eo[0     ] = y_lhuhvde | knep835je_uzqghqf | t__jcg4w9op | v64tquaebtsdj1cgmtr;  
  assign wfa5o72ctktgt55fgv2eo[1    ] = x3pdmlbidudtcfe | knep835je_uzqghqf | ufj54jrgxdnsw4v_ | v64tquaebtsdj1cgmtr  ;  
  assign wfa5o72ctktgt55fgv2eo[2   ] = md9w_qvcupymt5 ;  
  assign wfa5o72ctktgt55fgv2eo[3 ] = pdje7bg4uudiwmaizj;  
  assign wfa5o72ctktgt55fgv2eo[4     ] = x3pdmlbidudtcfe | y_lhuhvde | knep835je_uzqghqf | md9w_qvcupymt5 | pdje7bg4uudiwmaizj;  
  wire hn06o8bac7m4y72hse;
  assign wfa5o72ctktgt55fgv2eo[74-1:10   ] = hn06o8bac7m4y72hse ? xgg3cweyrd0uj_9ekh[64-1:0] : {{64-20-12{1'b0}}, txk1r9aiq_7l2nkw101w_, xgg3cweyrd0uj_9ekh[11:0]};  
  wire [64-1:0] xqt00lwbx__r_z4f6tfsp7 = wfa5o72ctktgt55fgv2eo[74-1:10];

  
  wire tfa79b6o6viuffzd    = mftzpw3hqrbum & pu7da028_tz7r;
  wire feaio68lvlpv0pv     = mftzpw3hqrbum & oogo4cx3q8tv9mbo;
  wire zalvrup6tbluro_t   = mftzpw3hqrbum & fpop_x33d6ai;
  wire plauwcknx568sxh4z   = mftzpw3hqrbum & h9ohvklruyeg;

  wire [74-1:0] f71s92bjwuhpisqhx13nk;
  assign f71s92bjwuhpisqhx13nk[5  ] = tvr8zxsmimyd3j7y4;  
  assign f71s92bjwuhpisqhx13nk[6  ] = rrki1m97jmtyk2r;  
  assign f71s92bjwuhpisqhx13nk[8  ] = v8lyodmb_xbnrq1r5f5vib_1;  
  assign f71s92bjwuhpisqhx13nk[9  ] = wkpz9dk71bcfhgjwdb1b;  
  assign f71s92bjwuhpisqhx13nk[7  ] = i1g4vxhyij_qk9u;  
  assign f71s92bjwuhpisqhx13nk[0     ] = plauwcknx568sxh4z;  
  assign f71s92bjwuhpisqhx13nk[1    ] = tfa79b6o6viuffzd | plauwcknx568sxh4z;  
  assign f71s92bjwuhpisqhx13nk[2   ] = feaio68lvlpv0pv    ;  
  assign f71s92bjwuhpisqhx13nk[3 ] = zalvrup6tbluro_t  ;  
  assign f71s92bjwuhpisqhx13nk[4     ] = tfa79b6o6viuffzd | feaio68lvlpv0pv | zalvrup6tbluro_t;  
  assign f71s92bjwuhpisqhx13nk[74-1:10   ] = xgg3cweyrd0uj_9ekh[64-1:0];  
 

  assign fdc8111sh6h232 = 1'b0 
                    | x3pdmlbidudtcfe   
                    | y_lhuhvde      
                    | knep835je_uzqghqf 
                    | md9w_qvcupymt5    
                    | pdje7bg4uudiwmaizj  
                    | tfa79b6o6viuffzd   
                    | feaio68lvlpv0pv    
                    | zalvrup6tbluro_t  
                    ;

  assign owhsxmah_o1vvv = 1'b0
                      | md9w_qvcupymt5
                      | pdje7bg4uudiwmaizj  
                      | feaio68lvlpv0pv    
                      | zalvrup6tbluro_t  
                      ; 

  wire lqmar0e = fdc8111sh6h232   
                 
               | plauwcknx568sxh4z  
               | v64tquaebtsdj1cgmtr
               | t__jcg4w9op     
               | ufj54jrgxdnsw4v_  
               ;


  assign canacnkc7zibtkn418i = f71s92bjwuhpisqhx13nk;
  assign x03ux1utw4qem5kk3c = wfa5o72ctktgt55fgv2eo;

  wire t8pnaxivsp11y;
  wire o1cudx277m8xr;
  wire stxr8fa544k8i6tqe;
  wire a5mvas76kenria5gi34;
  wire xszf10lmqmdfvdacx82;
  
  
  
  
  
  assign cn8o3075eju6dycby = 1'b0;
  
  
  
  
  
  
  
  
  
  
  

  assign zi39s8s7rmgo_lyocr_ = 1'b0;
  
  
  
  
  
  
  
  
  
  
  
  
  
  

  assign g1cek93tezrlyyt = 5'd0;
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  assign i22z6k7eo0it77lz2 = 64'b0;
  

  
  
  
  wire csvyewfoj_2dyhz       =   (
                               tfa79b6o6viuffzd  
                             | feaio68lvlpv0pv   
                             | zalvrup6tbluro_t 
                             | plauwcknx568sxh4z 
                            )
                           ;
  
  wire tujozwjl_1      = csvyewfoj_2dyhz;
  
  wire wsso1l3roo     =     (
                               x3pdmlbidudtcfe    
                             | y_lhuhvde       
                             | knep835je_uzqghqf  
                             | md9w_qvcupymt5     
                             | pdje7bg4uudiwmaizj   
                             | t__jcg4w9op      
                             | ufj54jrgxdnsw4v_   
                             | v64tquaebtsdj1cgmtr 
                            )
                           ;
  wire x6iacisl6_ir1ub      = wsso1l3roo;
 
  assign a601v24iimk0q23vf =  abniijg5zst5pbmx4q  
                       | szntcqan754qrdh 
                       | cll6ubptbwvtxo0lc
                       ;

  wire ktto7e9umj7dov;

  
  
  localparam rqzr_eaa  = 4'b0000; 
  localparam ioaaz4ufczj  = 4'b0001; 
  localparam fb7psuwcbwuti  = 4'b0010; 
  localparam fdma9st8q43nuns   = 4'b0011; 
  localparam qcpy4fycbt   = 4'b0100; 
  localparam r1t9p6mx_ra    = 4'b0101; 
  localparam c686_234if9z23e   = 4'b0110; 
  localparam ygm_h85q0x9n   = 4'b0111; 
  localparam fb3blm21_xwu   = 4'b1000; 

  wire [3:0] f8m0yygpetis;
  wire [3:0] tztm2dxlxm;
  wire gmvq6zbjfg;

  wire xntpwh2cyhb = (tztm2dxlxm == rqzr_eaa);
  wire vfxezjwbi8a = (tztm2dxlxm == ioaaz4ufczj);
  assign ktto7e9umj7dov = (tztm2dxlxm == fb7psuwcbwuti);
  wire tt7bgy6ulfeivcyf = (tztm2dxlxm == fdma9st8q43nuns);
  wire dalyz6cgj0a5uolc = (tztm2dxlxm == qcpy4fycbt);
  wire pxk8z0f1z4cgkbk = (tztm2dxlxm == fb3blm21_xwu);
  assign t8pnaxivsp11y = (tztm2dxlxm == ygm_h85q0x9n);
  wire jk0c_m61_wt35 = (tztm2dxlxm == r1t9p6mx_ra);
  wire nqzeiapkstv_5 = (tztm2dxlxm == c686_234if9z23e);

  assign ldj4m511gvpu12mdu1_ = xntpwh2cyhb;
  
  wire fn22ct7oo31a51601y;
  wire [3:0] wgrd6wm9974g7ezyq;
  wire n1jimlhvuntydx703f25ft;
  wire [3:0] c50tv7mimwy79;
  wire ms00q96_l_6ybkbpkdyd6h;
  wire [3:0] xmr18pucnal9xg;
  wire nbxih33qqt2yi461gczx;
  wire [3:0] icx1msle9uf5ow;
  wire twa5abff7v9zkqfjzf6yxle5;
  wire [3:0] fzq2ed9hkh092uvxvuz;
  wire x8aa4ng6e22soilavroar;
  wire [3:0] a82yw5un6rt36e4;
  wire q4kn7leuy6psrwb6eky3i9s;
  wire [3:0] qx31lq1cfib5uox;
  wire iwuvkevvdgv8nypv7v3;
  wire [3:0] i72_codnw9hftldm;
  wire i49b10h6halpyqw7129ml;
  wire [3:0] wr1x_jb8cte_n_3f6;

  
  assign fn22ct7oo31a51601y = xntpwh2cyhb & a601v24iimk0q23vf;
  assign wgrd6wm9974g7ezyq = ioaaz4ufczj;

  
  assign n1jimlhvuntydx703f25ft = vfxezjwbi8a & (tujozwjl_1 ? 1'b1 : x6iacisl6_ir1ub ? ~w2h8uh3l463qbgqmv : 1'b1); 
  assign c50tv7mimwy79 = tujozwjl_1 ? fdma9st8q43nuns : 
                        x6iacisl6_ir1ub ? (~fdc8111sh6h232 ? qcpy4fycbt : hn06o8bac7m4y72hse ? fb3blm21_xwu :  r1t9p6mx_ra) : 
                        fb7psuwcbwuti;

  
  assign ms00q96_l_6ybkbpkdyd6h = ktto7e9umj7dov;
  assign xmr18pucnal9xg = rqzr_eaa;

  
  assign nbxih33qqt2yi461gczx = tt7bgy6ulfeivcyf & bwbmafs1inesgjyn;
  assign icx1msle9uf5ow = rqzr_eaa;

  
  assign hn06o8bac7m4y72hse = ~fkuqlh34r | rrki1m97jmtyk2r | tvr8zxsmimyd3j7y4;
  assign twa5abff7v9zkqfjzf6yxle5 = dalyz6cgj0a5uolc & ydydp69z03wvr97;
  assign fzq2ed9hkh092uvxvuz = rqzr_eaa;

  
  wire fqxauxh4hyx_b;
  wire oge7q1uaup7yuy9t;
  assign iwuvkevvdgv8nypv7v3 = pxk8z0f1z4cgkbk;
  assign i72_codnw9hftldm = 
                          kqyojh1maxy0x834htg  ? ygm_h85q0x9n : 
                          fqxauxh4hyx_b           ? ygm_h85q0x9n :
                          oge7q1uaup7yuy9t          ? ygm_h85q0x9n :
                          qcpy4fycbt;

  
  assign i49b10h6halpyqw7129ml = t8pnaxivsp11y;
  assign wr1x_jb8cte_n_3f6 = rqzr_eaa;


  
  wire plgrerx7_ny1kdg16ie831 = hpk3eafyque5ubt_c62flnny & oyq1p3qa2iffjuqns0jkgg;
  assign x8aa4ng6e22soilavroar = jk0c_m61_wt35 & plgrerx7_ny1kdg16ie831;
  assign a82yw5un6rt36e4 = c686_234if9z23e;

  
  wire covhkab5l4p5vyb4_k5; 
  assign q4kn7leuy6psrwb6eky3i9s = nqzeiapkstv_5 & qjw2q0j88rjr42lautsqnca;
  assign qx31lq1cfib5uox = covhkab5l4p5vyb4_k5 ? ygm_h85q0x9n : fb3blm21_xwu;

 
  assign gmvq6zbjfg =   fn22ct7oo31a51601y
                   | n1jimlhvuntydx703f25ft
                   | ms00q96_l_6ybkbpkdyd6h
                   | nbxih33qqt2yi461gczx
                   | twa5abff7v9zkqfjzf6yxle5
                   | iwuvkevvdgv8nypv7v3
                   | i49b10h6halpyqw7129ml
                   | x8aa4ng6e22soilavroar
                   | q4kn7leuy6psrwb6eky3i9s
                   ; 

  assign f8m0yygpetis =   ({4{fn22ct7oo31a51601y}}   & wgrd6wm9974g7ezyq)
                   | ({4{n1jimlhvuntydx703f25ft}}   & c50tv7mimwy79)
                   | ({4{ms00q96_l_6ybkbpkdyd6h}}   & xmr18pucnal9xg)
                   | ({4{nbxih33qqt2yi461gczx}} & icx1msle9uf5ow)
                   | ({4{twa5abff7v9zkqfjzf6yxle5}} & fzq2ed9hkh092uvxvuz)
                   | ({4{iwuvkevvdgv8nypv7v3}} & i72_codnw9hftldm)
                   | ({4{i49b10h6halpyqw7129ml}} & wr1x_jb8cte_n_3f6)
                   | ({4{x8aa4ng6e22soilavroar}}  & a82yw5un6rt36e4)
                   | ({4{q4kn7leuy6psrwb6eky3i9s}} & qx31lq1cfib5uox)
                   ;

  ux607_gnrl_dfflr #(4) zy9agrte859 (gmvq6zbjfg, f8m0yygpetis, tztm2dxlxm, gf33atgy, ru_wi); 

  
  wire hd_fpok_kvptm7d9zjsjwhe = abniijg5zst5pbmx4q;
  wire sgkr3sgtoqp3j1_x6g8akcy82we = gmvq6zbjfg & (f8m0yygpetis == rqzr_eaa);
  wire xav3_b1w49lodyw3ky41uhgl = hd_fpok_kvptm7d9zjsjwhe | sgkr3sgtoqp3j1_x6g8akcy82we;
  wire p02zov_3lxukr7rlvks2yey = hd_fpok_kvptm7d9zjsjwhe | (~sgkr3sgtoqp3j1_x6g8akcy82we);

  ux607_gnrl_dfflr #(1) oskhizapxqhv0l8ntoatnxwwp7kkj7 (xav3_b1w49lodyw3ky41uhgl, p02zov_3lxukr7rlvks2yey, p2smibeuelrp8hsca6vc8w6q, gf33atgy, ru_wi); 

  
  wire on_xwis2hg9o98dsgj7cwwcgawhl = szntcqan754qrdh;
  wire pi3umaqf0w6ou0u47478zhk = gmvq6zbjfg & (f8m0yygpetis == rqzr_eaa);
  wire vzpk8ye3g8exn176vk94ipiu1 = on_xwis2hg9o98dsgj7cwwcgawhl | pi3umaqf0w6ou0u47478zhk;
  wire lg7idlpn50hhmmtxxoh2qrah = on_xwis2hg9o98dsgj7cwwcgawhl | (~pi3umaqf0w6ou0u47478zhk);

  ux607_gnrl_dfflr #(1) aibwxirks94c9cx41l2p9woghqhp (vzpk8ye3g8exn176vk94ipiu1, lg7idlpn50hhmmtxxoh2qrah, kidn1h9_lj8wzplj4kd32, gf33atgy, ru_wi); 

  
  wire kt2wlmxeega8v3xmxf04ais6hh6j = cll6ubptbwvtxo0lc;
  wire n4n65ty4ni_hr35_ymczpc2muc3 = gmvq6zbjfg & (f8m0yygpetis == rqzr_eaa);
  wire xnxki0uvry7vj4sadtlzrgfiu = kt2wlmxeega8v3xmxf04ais6hh6j | n4n65ty4ni_hr35_ymczpc2muc3;
  wire o4ib5rt87k4t4tdyb7zwvvjoe0 = kt2wlmxeega8v3xmxf04ais6hh6j | (~n4n65ty4ni_hr35_ymczpc2muc3);

  ux607_gnrl_dfflr #(1) dtk65gx3npsy9b2itpjt32vk59y0 (xnxki0uvry7vj4sadtlzrgfiu, o4ib5rt87k4t4tdyb7zwvvjoe0, gr5iv52qlkdgsjcutlh5ae, gf33atgy, ru_wi); 

  
  
  wire uys2_c7rmnm5gjf6t;
  wire yhte_l42subrkndmdewly6ed = a601v24iimk0q23vf;
  wire jgy2u9imfeirozi9eglwglq = gmvq6zbjfg & (f8m0yygpetis == rqzr_eaa);
  wire a8qosapxeb5vai1uy9s = yhte_l42subrkndmdewly6ed | jgy2u9imfeirozi9eglwglq;
  wire fvd4_fyn059jua6pp041uu5 = yhte_l42subrkndmdewly6ed | (~jgy2u9imfeirozi9eglwglq);

  ux607_gnrl_dfflr #(1) q5v2_zkz0s81_48ydhmm6gkl1d (a8qosapxeb5vai1uy9s, fvd4_fyn059jua6pp041uu5, uys2_c7rmnm5gjf6t, gf33atgy, ru_wi); 

  assign sl5f3k5g9ln8_zvzr = uys2_c7rmnm5gjf6t;

  
  
  
  
  
  
  
  assign x8rpm78rvvycis     = tt7bgy6ulfeivcyf;

  
  
  
  
  
  
  
  assign sxhicsqvufwfbnk0     = dalyz6cgj0a5uolc;

  

  assign vs6ryzcr0bwqs5so = pxk8z0f1z4cgkbk;
  assign j25ub196dc_agl8oovaex4 = xqt00lwbx__r_z4f6tfsp7[32-1:0];
  assign pi2nokcm8qf7och7l4g = md9w_qvcupymt5;   
  assign c0i0hs5tz64_ce5f0z = 1'b0; 
  assign dmzdczrqcueolg3dzufj_by5rmf = v8lyodmb_xbnrq1r5f5vib_1; 
  assign a1sqko6fok9qzpbtyuw0 = rrki1m97jmtyk2r;
  assign bquohubxiv2rsayn62v = tvr8zxsmimyd3j7y4;

  wire t7_wd7s1ayipd6fch8xgh3n = pxk8z0f1z4cgkbk | t8pnaxivsp11y; 
  wire rffe_iwy5__m2ffjdoobl = pxk8z0f1z4cgkbk ? kqyojh1maxy0x834htg : 1'b0; 

  ux607_gnrl_dfflr #(1) oj9q5dmh_sl7oq7rtr_bw5 (t7_wd7s1ayipd6fch8xgh3n, rffe_iwy5__m2ffjdoobl, stxr8fa544k8i6tqe, gf33atgy, ru_wi);



  
  

  
  wire       vgsz5pn_3kjggra6ueuqr_;
  wire [1:0] w01sf2h97q68k5msmjfsgb;
  wire       sho0i24sqotphrb09e3c0yy;
  wire       b9qdzfuqngpv3oj8qn60ex;
  wire       pvfop2o8otpcjkgqm3v6eswr;

  ux607_gnrl_dfflr #(1) mv4wlq4ofhg017onppr9klih6dij (hmtyprargqxng, rm1dxjejhq7dh3q5m, vgsz5pn_3kjggra6ueuqr_, gf33atgy, ru_wi); 
  ux607_gnrl_dfflr #(2) rijb7rgg2svtjlvt01ru45n0qpl_m23  (hmtyprargqxng, st2zalpx0uf,  w01sf2h97q68k5msmjfsgb,  gf33atgy, ru_wi); 
  ux607_gnrl_dfflr #(1) h9v2r6d_4zj8mhd3d2eyxuz3xzce8  (hmtyprargqxng, ni01kj42oob2x,  sho0i24sqotphrb09e3c0yy,  gf33atgy, ru_wi); 
  ux607_gnrl_dfflr #(1) wkaacv0eoxtx3ng18e8ebfd8ao2xnq  (hmtyprargqxng, ah8kjlmvnaxzbi,  b9qdzfuqngpv3oj8qn60ex,  gf33atgy, ru_wi); 
  ux607_gnrl_dfflr #(1) z85rcd1mtc57uoogknsh9mmrl6a   (hmtyprargqxng, sxvvsxtbhyvt,   pvfop2o8otpcjkgqm3v6eswr,   gf33atgy, ru_wi); 


  wire x0j1djmcr7nvs77eqi_6;
  wire ba_mmm9llu4g4hxtzc3jfsiqk9f;
  assign covhkab5l4p5vyb4_k5 =  x0j1djmcr7nvs77eqi_6
                          | ba_mmm9llu4g4hxtzc3jfsiqk9f
                          ;

  assign hpk3eafyque5ubt_c62flnny = jk0c_m61_wt35; 
  assign sfezv1xz2ghvo8pkt = b7kat6xkt_rgc2hdogj3k[27-1+12:12]; 
  assign frzfsbt7hp3n4aj3zvvumnh0s = b7kat6xkt_rgc2hdogj3k[64-1 : 27+12-1]; 
  assign vagaza053272juvmo59v8w20s = {1'b0, i1g4vxhyij_qk9u}; 
  assign rzf45534z36ejq96260 = tvr8zxsmimyd3j7y4; 
  assign zkuxqezrmlhyyjjgx = b7kat6xkt_rgc2hdogj3k; 
  assign u3h5tvu1g2q93141j9o = 64'b0; 
  assign pjh0wad7t_5du3cync_0c = 1'b0; 
  assign wmkgrgf631pbq = 1'b0; 


  wire [1:0] e5suv95h3yjoa = {1'b0, i1g4vxhyij_qk9u};

  cqpjxz2qb247thego6htwvkw_aiu lpcbtkgnuc86ae4xr8g1d9jqhojv_j(
  .f_8ecse5wf0jrndlozy2070bja                       (qjw2q0j88rjr42lautsqnca              ),        
  .e4sprh35cvfb6sw6lnskyaga91                    (imkm56ujne9v4m6n08w1yf5622           ),
  .qrvtg_49_dmoggu94orq0                        (ih4hmwugasiodbx5da9_40kx               ),         
  .iocew24g1qos_gvi3_r3uoqfdf                        (x5vjq7mshfwr0h3q514t7mhdt               ),         
  .qh_y92pv7dp1us9t5wxdmm57                        (qrxtk7e03100_uwkx73sg7               ),         
  .cznjry8adajzgi6gkmyr830m_u                        (i7qiq2q9c6hbeful9qu9lb               ),         
  .ugixcggahb26m1glzpuqvpq                        (yr0s3skqk7cdqflsrbsxg9znu               ),         
  .vbpz6tidsg3o93kih6nmamlyg9wmr1zz                  (adqieke11qo0elfz93hlouwjc0         ),   
  .j2dtuvq0m4iir947lery9tpxqwhjj2g3                (w93gdpnnxuydy53eu0s9nxw7xdct7       ), 
  .wzqcq7ug3_gv3tuf0o                           (1'b0                               ),
  .ng5gq72xr47fw8fztwfo8hw                         (vgsz5pn_3kjggra6ueuqr_              ), 
  .cmyy3ooatm0bn2s6fv8_r                          (w01sf2h97q68k5msmjfsgb               ), 
  .ckgybqpbvuzwgxv1ixd_6rpf                          (sho0i24sqotphrb09e3c0yy               ),
  .nguthky_k_yqsf8fa9btry1                          (b9qdzfuqngpv3oj8qn60ex               ),
  .w30ye15yns15                                     (e5suv95h3yjoa                       ),
  .jyl_xsaj6z1u9wndwpi                               (pvfop2o8otpcjkgqm3v6eswr                ),
  .idg19n7mm21jtb                                  (tvr8zxsmimyd3j7y4                     ),
  .o_4mw1alrjmdzl                                 (x0j1djmcr7nvs77eqi_6               ),
  .nkjxsm02z2_q5_0_                               (ba_mmm9llu4g4hxtzc3jfsiqk9f             ),
  .gf33atgy                                          (gf33atgy                                ),
  .ru_wi                                        (ru_wi                              )
);



  wire z2_i1jboefgvd3i6evnwsj5 = nqzeiapkstv_5 | t8pnaxivsp11y;
  wire xbgwtlk5_9oiewa9xdpqf5bfa = nqzeiapkstv_5 ? x0j1djmcr7nvs77eqi_6 : 1'b0;
  ux607_gnrl_dfflr #(1) r8khybyteg83hxbcovhw06hpe (z2_i1jboefgvd3i6evnwsj5, xbgwtlk5_9oiewa9xdpqf5bfa, a5mvas76kenria5gi34, gf33atgy, ru_wi);

  wire m0lr0ty_ia3x1g5cpqna424 = nqzeiapkstv_5 | t8pnaxivsp11y;
  wire gz3vuyxkdvci4hhp9u1kt3n1dgk = nqzeiapkstv_5 ? ba_mmm9llu4g4hxtzc3jfsiqk9f : 1'b0;
  ux607_gnrl_dfflr #(1) f2yexm49yp76lguh0qta0yk1maf (m0lr0ty_ia3x1g5cpqna424, gz3vuyxkdvci4hhp9u1kt3n1dgk, xszf10lmqmdfvdacx82, gf33atgy, ru_wi);




  assign o1cudx277m8xr = 1'b0 
                     | a5mvas76kenria5gi34  
                     | xszf10lmqmdfvdacx82 
                     | stxr8fa544k8i6tqe
                     ;


  
  
wc2lipjaiimwuy7fx9zp32mr  lbpbwc1x5lhcs71rg3inpdi1d2xu(
     .e98zc_xde8d   (xqt00lwbx__r_z4f6tfsp7[32-1:0]),
     .lms849k     (fqxauxh4hyx_b ),
     .dhzk00cwbk (oge7q1uaup7yuy9t)
  );





  assign td1nncrrbp273gpbj6cq = bwbmafs1inesgjyn & bkkiffh6ob85nh79doya_ ? 
                                 (
                                    qhqqh0lyehgtfop1tc[0]   ? 3'd1 :   
                                    qhqqh0lyehgtfop1tc[1]   ? 3'd2 :   
                                    qhqqh0lyehgtfop1tc[2]   ? 3'd3 :   
                                    qhqqh0lyehgtfop1tc[3]   ? 3'd4 :   
                                                              3'd0 
                                 ) :
                              ydydp69z03wvr97 & pjic5x84bqxpvdduy4r2s ?
                                 (
                                    w5az87bw32r0tjbo0tdrv2ouvx ? 3'd3 :   
                                                              3'd1     
                                 ) :
                              t8pnaxivsp11y ?                 3'd2 :
                                                              3'd0 ;   
  
  assign en1q7v03lnxlj7aw4dpakyg0 = bwbmafs1inesgjyn | ydydp69z03wvr97 | t8pnaxivsp11y;
  assign igimbt9i77_wg1s8b6 = en1q7v03lnxlj7aw4dpakyg0;

  

  ux607_gnrl_dfflr #(1) o972gi91r4j36ftxumx4lvxdnwa8 (hmtyprargqxng, cbbcxlflqkqoklckuekt, v8lyodmb_xbnrq1r5f5vib_1, gf33atgy, ru_wi); 
  ux607_gnrl_dfflr #(1) w48e7wdkr9y2kf0u_x10p (hmtyprargqxng, lodtxdqjnwvx, rrki1m97jmtyk2r, gf33atgy, ru_wi); 
  ux607_gnrl_dfflr #(1) b3c3qdin2ugiu0wv08z6 (hmtyprargqxng, z28w9as50xav1c2ms, tvr8zxsmimyd3j7y4, gf33atgy, ru_wi); 


  ux607_gnrl_dfflr #(1) nbf3cjdgpo9x7njxtdu0lu1v4 (hmtyprargqxng, ewe_b1wv9zhrc8rc6hhr, wkpz9dk71bcfhgjwdb1b, gf33atgy, ru_wi); 
  ux607_gnrl_dfflr #(1) ozt5t1pvs5eulpi7bs08 (hmtyprargqxng, n37wgp2u95gc5b_, i1g4vxhyij_qk9u, gf33atgy, ru_wi); 




endmodule




















module r5e39tculmqtcj5 (
  input [31:0] ticq8ng,
  input [31:0] y4a7pqq0kkz,
  input nn8hi7fy9,

  output uwkhmy2e_yju,
  output k1fnd9t0fsu,
  output la186rvvv7gcy,
  output kd65qo8qkm0kgmw,
  output a7atgbs19h1,
  output kzl0hy0qswsidji5,
  output boll1pzurodbj,
  output kt7mps652so,
  output em08qdw,
  output fij5gpv,

  output [9:0] tcfrqq029
);

wire wtomt4uy4ek = nn8hi7fy9 ? ticq8ng[31] : y4a7pqq0kkz[31];

wire eecpw_svltkog5 = nn8hi7fy9 ? (ticq8ng[30:20] == 11'h7FF) : (y4a7pqq0kkz[30:23] == 8'hFF);

wire y4n9i2ze4fjy04 = nn8hi7fy9 ? (ticq8ng[30:20] == 11'h000) : (y4a7pqq0kkz[30:23] == 8'h00);

wire nl14snhbt2qj = nn8hi7fy9 ? ({ticq8ng[19:0],y4a7pqq0kkz} == 52'b0) : (y4a7pqq0kkz[22:0] == 23'b0);

wire c5969aj90uti = y4n9i2ze4fjy04 & (~nl14snhbt2qj);

wire q8cfxdt_ = nn8hi7fy9 ? ticq8ng[19] : y4a7pqq0kkz[22];

wire wnbogvv = (~eecpw_svltkog5) & (~y4n9i2ze4fjy04);

assign em08qdw = eecpw_svltkog5 & (~nl14snhbt2qj) & (~q8cfxdt_);

assign fij5gpv = eecpw_svltkog5 & (~nl14snhbt2qj) & q8cfxdt_;

wire zwtvtr2 = fij5gpv | em08qdw;

wire ijny0n8caa = eecpw_svltkog5 & nl14snhbt2qj;

wire mwdn3z1 = (y4n9i2ze4fjy04 & nl14snhbt2qj);

assign kd65qo8qkm0kgmw = mwdn3z1 & wtomt4uy4ek;
assign a7atgbs19h1 = mwdn3z1 & (~wtomt4uy4ek);

assign la186rvvv7gcy = c5969aj90uti & wtomt4uy4ek;
assign kzl0hy0qswsidji5 = c5969aj90uti & (~wtomt4uy4ek);

assign k1fnd9t0fsu = wnbogvv & wtomt4uy4ek;
assign boll1pzurodbj = wnbogvv & (~wtomt4uy4ek);

assign uwkhmy2e_yju = ijny0n8caa & wtomt4uy4ek;
assign kt7mps652so = ijny0n8caa & (~wtomt4uy4ek);



assign tcfrqq029 [0] = uwkhmy2e_yju;

assign tcfrqq029 [1] = k1fnd9t0fsu;

assign tcfrqq029 [2] = la186rvvv7gcy;

assign tcfrqq029 [3] = kd65qo8qkm0kgmw;

assign tcfrqq029 [4] = a7atgbs19h1;

assign tcfrqq029 [5] = kzl0hy0qswsidji5;

assign tcfrqq029 [6] = boll1pzurodbj;

assign tcfrqq029 [7] = kt7mps652so;

assign tcfrqq029 [8] = em08qdw;

assign tcfrqq029 [9] = fij5gpv;

endmodule




















module swhs3pkf0sfg9ix (
    input  gf33atgy,
    input  ru_wi,
    input  cr7bv45kj7l,
    input  [31:0] ticq8ng,
    input  [31:0] y4a7pqq0kkz,
    input  v659v2hvrtej,
    input  p940nw4duiie64,
    input  ersv4d_m80ir1,
    input  lc9pop79cuks,
    input  af8gggx2rbk5w,
    input  z9ydb68fp_la3j,
    input  im1jxeoei8g,
    input  c2o9xduz06,
    input  azpnhv65b4,
    input  ji57bityrdt,
    input  ex14gbip3a,
    input  f_xw6g_ldgz,
    input  cix9qipqelc7k,
    input  wpio23m13to3o0,
    input  u9bwc77pa3,
    input  k937n2wbqgq,
    input  ayc3vpo7,
    input  goy441jl,
    input  [2:0] vc529nuu,
    output [63:0] uiwlxd,
    output [4:0] adnx9wgdt2

);

  
  wire nn8hi7fy9 = ersv4d_m80ir1 
                | lc9pop79cuks 
                | ex14gbip3a 
                | f_xw6g_ldgz 
                | ayc3vpo7;

   wire v0da13u6ykrw = nn8hi7fy9 ? (ticq8ng[30:20] == 11'h7FF) : (y4a7pqq0kkz[30:23] == 8'hFF);
   wire rg17tsy6wwx = nn8hi7fy9 ? (ticq8ng[30:20] == 11'h000) : (y4a7pqq0kkz[30:23] == 8'h00);
   wire wb75liyzd6vmew7 = nn8hi7fy9 ? ({ticq8ng[19:0],y4a7pqq0kkz} == 52'b0) : (y4a7pqq0kkz[22:0] == 23'b0);
   wire bml43dgqbvm = rg17tsy6wwx & (~wb75liyzd6vmew7);
   wire ib3hkx1k0t = nn8hi7fy9 ? ticq8ng[19] : y4a7pqq0kkz[22];
   wire mgvwdehh1 = (~v0da13u6ykrw) & (~rg17tsy6wwx);
   wire aswm0l3tr55 = v0da13u6ykrw & (~wb75liyzd6vmew7) & (~ib3hkx1k0t);
   wire r41nzg = v0da13u6ykrw & (~wb75liyzd6vmew7) & ib3hkx1k0t;
   wire jqgto = r41nzg | aswm0l3tr55;
   wire ak6syfq = v0da13u6ykrw & wb75liyzd6vmew7;
   wire sy1qjmixh5e = (rg17tsy6wwx & wb75liyzd6vmew7);

   wire [51:0]  jd1t0763x = {ticq8ng[19:0],y4a7pqq0kkz};
   wire [22:0]  lkish79hpt = y4a7pqq0kkz[22:0];
   wire [10:0]  vropxwawb = ticq8ng[30:20];
   wire [ 7:0]  dbw_bap_jqyl = y4a7pqq0kkz[30:23];
   wire         rhaf675bn = ticq8ng[31];
   wire         a8rijdb567ulj = y4a7pqq0kkz[31];


   wire [51:0]  d86mct = nn8hi7fy9 ? jd1t0763x : {lkish79hpt,29'b0};
   wire         mp3k_c3d = nn8hi7fy9 ? rhaf675bn : a8rijdb567ulj;
   wire [10:0]  eff76eu5r  = nn8hi7fy9 ? vropxwawb  : {3'b0,dbw_bap_jqyl};

   wire zpwosdnwv0 = ak6syfq & (~mp3k_c3d);
   wire h2pw9rtks0i = ak6syfq & mp3k_c3d;

   wire eqi5fiol = sy1qjmixh5e & (~mp3k_c3d);
   wire kc2obnf0fo = sy1qjmixh5e & mp3k_c3d;

  wire [3-1:0] hr6uuvr3izh;
  wire  hr_5q_o87l78el0;
  wire  rau7b3otce5zq;
  wire  pz73hz7q5h3oazsw;
  wire  ieq_x45icc_ygmzwu;
  wire  dmqidngg044lka0;
  wire  f4vcs6htny8xk9;
  wire  fj4nn1kh724bow;
  wire  chfklna44pacjcho;
  wire  s4mabzvk_lget7;
  wire  ade81kyp0620xstvq;
  wire  sn7ynh0j2u8h61;
  wire  uq85gpt70wdca;
  wire  dah1__e5zjv47wr;
  wire  zvw_q5tgix3s69c7o;
  wire  xurhhleqgmg8sy2;
  wire  rpn9v9ketinrb4o7oj;
  wire  hbc9h8mi5tp   ;
  wire  v41vgtsgcvch   ;
  wire  axgk4peda4gp   ;
  wire  bwqs5m4om61   ;
  wire  z1iavptcuyb   ;
  wire  sjt2wedeei_gmt0 ;
  wire  pdw2zx8bnrucv    ;
  wire  vnyuwuzda74sk9_  ;
  wire  se2fv2m60n1xym  ;
  wire  l4tu2pzv06wzg  ;
  wire  u75k9olcw2ovrh  ;
  wire  scjp5ckdygufd  ;
  wire  kcx64rdtzypzm  ;

  ux607_gnrl_dfflr #(3)    w5g6z591t60kamo(cr7bv45kj7l, vc529nuu  , hr6uuvr3izh  , gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1) dxm2rxi700ckuyplrd9 (cr7bv45kj7l, af8gggx2rbk5w, hr_5q_o87l78el0, gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1) v0knvpxc99h7mlx (cr7bv45kj7l, z9ydb68fp_la3j, rau7b3otce5zq, gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1) o5vbo36d6bi14deust (cr7bv45kj7l, im1jxeoei8g, pz73hz7q5h3oazsw, gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1) xj2i7kq2ilqr_tfz (cr7bv45kj7l, c2o9xduz06, ieq_x45icc_ygmzwu, gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1) cobhlfgdb0z_d6e (cr7bv45kj7l, v659v2hvrtej, dmqidngg044lka0, gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1) w_z54b32w1zg97gzisf0 (cr7bv45kj7l, p940nw4duiie64, f4vcs6htny8xk9, gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1) oik2q5uhh3r9a0a (cr7bv45kj7l, ersv4d_m80ir1, fj4nn1kh724bow, gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1) mkzgmnso8mgy5fu4 (cr7bv45kj7l, lc9pop79cuks, chfklna44pacjcho, gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1) mi37kjxy4xy0pf38tfo(cr7bv45kj7l, cix9qipqelc7k,s4mabzvk_lget7,gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1) u4tn2l1jthbizby6djz2(cr7bv45kj7l, wpio23m13to3o0,ade81kyp0620xstvq,gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1) s0hbuk2m76gddf53pym0u(cr7bv45kj7l, u9bwc77pa3,sn7ynh0j2u8h61,gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1) qfu28sbumblvg5ay76w(cr7bv45kj7l, k937n2wbqgq,uq85gpt70wdca,gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1) k5n30u66sp8d3z2p9p1h(cr7bv45kj7l, azpnhv65b4,dah1__e5zjv47wr,gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1) k3ikqtussshkh0go2(cr7bv45kj7l, ji57bityrdt,zvw_q5tgix3s69c7o,gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1) uh18x9e2uac079645(cr7bv45kj7l, ex14gbip3a,xurhhleqgmg8sy2,gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1) xxn6f86bw0utb4cti(cr7bv45kj7l, f_xw6g_ldgz,rpn9v9ketinrb4o7oj,gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1)    yq0y4mugwn2ud_m (cr7bv45kj7l, mp3k_c3d   , hbc9h8mi5tp   , gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1)    lfai2_hbgs7svna (cr7bv45kj7l, r41nzg   , v41vgtsgcvch   , gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1)    ha22lz3ge_tccsx (cr7bv45kj7l, aswm0l3tr55   , axgk4peda4gp   , gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1)    drxv7bef_c07bkk2s (cr7bv45kj7l, ak6syfq   , bwqs5m4om61   , gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1)    a8zt_cg79_f45y_e (cr7bv45kj7l, mgvwdehh1   , z1iavptcuyb   , gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1)  z6_5wmkudbfxd64 (cr7bv45kj7l, bml43dgqbvm , sjt2wedeei_gmt0 , gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1)     fqczcw2y69vxl (cr7bv45kj7l, jqgto    , pdw2zx8bnrucv    , gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1)   lx5lwcr9rqcfcn7m2p (cr7bv45kj7l, zpwosdnwv0  , vnyuwuzda74sk9_  , gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1)   gypcrav_osuorfday (cr7bv45kj7l, h2pw9rtks0i  , se2fv2m60n1xym  , gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1)   lvk7jedln7pqpdq (cr7bv45kj7l, eqi5fiol  , l4tu2pzv06wzg  , gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1)   kmp7vp7wu5v3lbt (cr7bv45kj7l, kc2obnf0fo  , u75k9olcw2ovrh  , gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1)   k4cjm8u5ws78u (cr7bv45kj7l, ayc3vpo7  , scjp5ckdygufd  , gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1)   p0k5c0vf3uy7ty (cr7bv45kj7l, goy441jl  , kcx64rdtzypzm  , gf33atgy, ru_wi);

   wire [64-1:0] spdu2kgfxi4hwqf5 = 64'h7FF80000_00000000;
   wire [32-1:0] yalqc1omcjhx6 = 32'h7FC00000;
   wire [64-1:0] l1gpd_rq1zeu6   = 64'h7FF00000_00000000;
   wire [64-1:0] tm080y4ksbj0jwufg   = 64'hFFF00000_00000000;
   wire [32-1:0] t56x59ztjm5zwnj56   = 32'h7F800000;
   wire [32-1:0] vembz3jnjwpwx   = 32'hFF800000;
   wire [64-1:0] uk4q4m8jvw0d8zp   = 64'h00000000_00000000;
   wire [64-1:0] wzqga1virp_encj   = 64'h80000000_00000000;
   wire [32-1:0] d40417qihw6rqg   = 32'h00000000;
   wire [32-1:0] ywnvnrprlg65x3uq   = 32'h80000000;







   
   
   
   
   
   
   
        
   wire wp_xp_nm2j7az = v659v2hvrtej | p940nw4duiie64 | ersv4d_m80ir1 | lc9pop79cuks;
   wire jzx0y049lp5cy0v= azpnhv65b4 | ji57bityrdt | ex14gbip3a | f_xw6g_ldgz;

   wire [52:0]  xf92vp2m3d = {mgvwdehh1, d86mct};

   wire [10:0] wvvpiph = nn8hi7fy9 ? 11'd1023 : 11'd127;



   wire [11:0] mvpt9rw8vb52stdz38p;
   wire [11:0] l1l1j1q86l7rjr2j;
   wire b7al416lol277;
   
   wire [11:0] xzraqync_3fsxk9k_3teii55y2 = {1'b0,eff76eu5r}   ;
   wire [11:0] eb0ctt_nl3e3d7d1w_4p9n7x93 = (~{1'b0,wvvpiph });
   wire        vc000h9sulun8dpbf0bz5fzxls = 1'b1;
   
   wire        i83vn2g75rui4ede6j9ioa70ugp = (wp_xp_nm2j7az | jzx0y049lp5cy0v);       
   wire [11:0] szdt_u65giz7 = mvpt9rw8vb52stdz38p[11:0];
   
   wire [11:0] jdn4wx2w8tno0b61k_srrv = {1'b0,wvvpiph }   ;
   wire [11:0] dslntpb2kksdjgkt0powur_ = (~{1'b0,eff76eu5r});
   wire        biyo66wdgpupq01jhemo3lq0 = 1'b1;
   
   wire        amxnkuchi7l1_0kudwvt84gbi = (wp_xp_nm2j7az | jzx0y049lp5cy0v);       
   wire [11:0] vyj0dzwxv00l94e = l1l1j1q86l7rjr2j[11:0];

   wire hw84i0_d96enyp517ctg = (vyj0dzwxv00l94e == 12'd1);
   wire s0xxswrrovk5qfz7tiaa = (vyj0dzwxv00l94e == 12'd2);

   wire [10:0] rd7fl26_y5h = szdt_u65giz7[11] ? vyj0dzwxv00l94e[10:0] : szdt_u65giz7[10:0];
   wire qjq45_mvimn5 = (~szdt_u65giz7[11]);
       
   wire h_qbebb = qjq45_mvimn5 & (|szdt_u65giz7[10:7]);
   wire [127:0] mejh707tq;
   wire [52:0]  fiyap2f_ig_f;

   wire [180:0] jkxd7ftbbh3xspajh = {128'b0,xf92vp2m3d};
   wire [  6:0] tzyyizq0dvvice8zgo5_n = szdt_u65giz7[6:0];
   
   wire         ejaudkhb58i42o3ci78 = (wp_xp_nm2j7az | jzx0y049lp5cy0v);       
   wire [180:0] joviasnyqgggsfacl;
   wire [180:0] iws06ubcqffir0mqtxhl7l = joviasnyqgggsfacl;

   assign {mejh707tq, fiyap2f_ig_f} = joviasnyqgggsfacl;


       
   wire [128:0] nxgosqul = (~qjq45_mvimn5) ? 129'b0 : {mejh707tq[127:0],fiyap2f_ig_f[52]};
   wire [63:0] d21dzbu556kk4rkuqye = jzx0y049lp5cy0v ? nxgosqul[63:0] : {32'b0,nxgosqul[31:0]};

   wire a5_ly4ex5a71hcq24a2jf = |fiyap2f_ig_f[49:0];

   wire f6dc_rhcaz;

   wire pazpiknp4h1    = qjq45_mvimn5 ? nxgosqul[0]          : 1'b0;
   wire g2sc17nqw10  = qjq45_mvimn5 ? fiyap2f_ig_f[51]     : hw84i0_d96enyp517ctg ? xf92vp2m3d[52]   : s0xxswrrovk5qfz7tiaa ? 1'b0             : 1'b0            ;
   wire etltckdy1zv  = qjq45_mvimn5 ? fiyap2f_ig_f[50]     : hw84i0_d96enyp517ctg ? xf92vp2m3d[51]   : s0xxswrrovk5qfz7tiaa ? xf92vp2m3d[52]   : 1'b0            ;
   wire a7e2y8e5thkno7f = qjq45_mvimn5 ? a5_ly4ex5a71hcq24a2jf : hw84i0_d96enyp517ctg ? (|xf92vp2m3d[50:0]) : s0xxswrrovk5qfz7tiaa ? (|xf92vp2m3d[51:0]) : (|xf92vp2m3d[52:0]);

   el7n_zz16sk_ntvue9v wjyg9zves44l3osv1y9 (
       .l      (pazpiknp4h1), 
       .g      (g2sc17nqw10 ),
       .r      (etltckdy1zv ),
       .s      (a7e2y8e5thkno7f),
       .ly53de   (mp3k_c3d),
       .nfj6b     (vc529nuu),
       .f6dc_rhcaz (f6dc_rhcaz) 
   );


  
  wire bip07ip5l5ft3aa2t3s4 = (|nxgosqul[128:64]) | (wp_xp_nm2j7az ? |nxgosqul[63:32] : 1'b0);
  wire e6axxabwbo852 = dmqidngg044lka0 | f4vcs6htny8xk9 | fj4nn1kh724bow | chfklna44pacjcho;
  wire gj1k4_k7peyb= dah1__e5zjv47wr | zvw_q5tgix3s69c7o | xurhhleqgmg8sy2 | rpn9v9ketinrb4o7oj;
  assign b7al416lol277 = cr7bv45kj7l & (wp_xp_nm2j7az | jzx0y049lp5cy0v);

  
  wire dzbfnnjnu5c2vi;
  wire w4ntspj0bg6ql8opwen7v55sa;
  wire [63:0] rwee3l_yahi8zjq8y_6six;
  wire v2yut51ojed2 ;
  wire enog_chi0waara08l    ;
  wire ia7awt7a85f2x8zfe  ;
  wire mjc2ko9ue08hnfniz8  ;
  wire v6p6tk4wn1g_mj7 ;

  ux607_gnrl_dfflr #(1)             q31xk608uoot9gf374t(b7al416lol277, f6dc_rhcaz               , dzbfnnjnu5c2vi            , gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1)  aykvry6minck1aikyhd9rgwgnkuah(b7al416lol277, bip07ip5l5ft3aa2t3s4 , w4ntspj0bg6ql8opwen7v55sa , gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(64)    rp7ls6ttig0_lmru708upgof6(b7al416lol277, d21dzbu556kk4rkuqye       , rwee3l_yahi8zjq8y_6six    , gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1)            cbhmwd7l2g2ayjv(b7al416lol277, h_qbebb              , v2yut51ojed2           , gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1)          bqtkvonczhgb7trgbqs(b7al416lol277, pazpiknp4h1            , enog_chi0waara08l         , gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1)        tk03rbxk1mwphqha_y7o(b7al416lol277, g2sc17nqw10          , ia7awt7a85f2x8zfe       , gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1)        cviqp1fply7uru_ulbl30b(b7al416lol277, etltckdy1zv          , mjc2ko9ue08hnfniz8       , gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1)       t2wk2yxwjc7g0vuadmzcz7(b7al416lol277, a7e2y8e5thkno7f         , v6p6tk4wn1g_mj7      , gf33atgy, ru_wi);



  wire [63:0] fbz5m81mktdw4uhv;
  wire        y2br9ri7kni_unin;











   wire [63:0] mk5gl3ippdiih78z_h8_ngwbgpt = rwee3l_yahi8zjq8y_6six[63:0];
   wire [63:0] qaufsfnnc9i8ce5deb847cksm = 64'b0;
   wire        mb8tn3wn2iqxl5a0jirs0h = dzbfnnjnu5c2vi;

   wire        z7zzynt4p6n91ltyfzw88yr = e6axxabwbo852 | gj1k4_k7peyb;

   wire [63:0] y4yutdej0620pote;
   wire        bb977ptd1fyw2vzt;
   wire [63:0] gflb0dmv454sowt17bx;
   wire        lgz5ovlgwou4qwx6k71sq;

   assign {y2br9ri7kni_unin,fbz5m81mktdw4uhv} = {bb977ptd1fyw2vzt,y4yutdej0620pote};

   wire c90da34p3x7kbsitpwjm = fbz5m81mktdw4uhv[32]; 
   

   wire s5v59vnb7umvyym6nbwlh0q4 = v2yut51ojed2 | w4ntspj0bg6ql8opwen7v55sa | (gj1k4_k7peyb ? y2br9ri7kni_unin : c90da34p3x7kbsitpwjm);

   wire a5ju5vvapnv = dmqidngg044lka0 | fj4nn1kh724bow;
   wire vrh7fcmgexv = dah1__e5zjv47wr | xurhhleqgmg8sy2;
   wire armn6_2e5hdgso = zvw_q5tgix3s69c7o | rpn9v9ketinrb4o7oj;

   wire llz0g84mdu21zmq = (~hbc9h8mi5tp) & s5v59vnb7umvyym6nbwlh0q4;
      
   wire fqmrukd2bhi20ngh6jl = (~(|fbz5m81mktdw4uhv)) & (~s5v59vnb7umvyym6nbwlh0q4);
   wire ulou78bd89d6sgy = hbc9h8mi5tp & (~fqmrukd2bhi20ngh6jl);
   wire x40te217wy90wsvbzda2r7n = fbz5m81mktdw4uhv[63];  
   wire ouw65j55ve26l_xayvvr8lvlb = fbz5m81mktdw4uhv[31];   
   wire cbmn5rtjbb68qbo = (~hbc9h8mi5tp) & (s5v59vnb7umvyym6nbwlh0q4 | (gj1k4_k7peyb ? x40te217wy90wsvbzda2r7n : ouw65j55ve26l_xayvvr8lvlb));
   wire mojy8yz4lgbnb2vi = hbc9h8mi5tp & (s5v59vnb7umvyym6nbwlh0q4 | (gj1k4_k7peyb ? (fbz5m81mktdw4uhv[63] & (|fbz5m81mktdw4uhv[62:0])) : (fbz5m81mktdw4uhv[31] & (|fbz5m81mktdw4uhv[30:0]))));

   wire [63:0] olk58do8mpdp18e6zbw2zzcwa = ~fbz5m81mktdw4uhv;
   wire [63:0] d4_gebt1q1dsvf_bvc3a0 = 64'b0;
   wire        c5381srmbn8numzwdtbkoy_9_4 = 1'b1; 
   
   
   
   
   
   

   wire        bkz3ex8j6dty_vo9us5iq9r = e6axxabwbo852 | gj1k4_k7peyb;

   
   
   
   wire [63:0] s25c523vk8wbn3kssl = gflb0dmv454sowt17bx;

   wire [63:0] hhqjnbrw2zq = cbmn5rtjbb68qbo ? (vrh7fcmgexv ? {32'h7FFF_FFFF,32'hFFFF_FFFF} : {32'h0000_0000,32'h7FFF_FFFF}): 
                          mojy8yz4lgbnb2vi ? (vrh7fcmgexv ? {32'h8000_0000,32'h0000_0000} : {32'hFFFF_FFFF,32'h8000_0000}):  
                          hbc9h8mi5tp  ? (vrh7fcmgexv ? s25c523vk8wbn3kssl : {{32{s25c523vk8wbn3kssl[31]}},s25c523vk8wbn3kssl[31:0]}):
                                         fbz5m81mktdw4uhv;
   wire [63:0] lii58p0oecj8xmc3 = llz0g84mdu21zmq ? {32'hFFFF_FFFF,32'hFFFF_FFFF} : 
                          ulou78bd89d6sgy ? {32'h0000_0000,32'h0000_0000} :  
                                         (armn6_2e5hdgso ? fbz5m81mktdw4uhv : {{32{fbz5m81mktdw4uhv[31]}},fbz5m81mktdw4uhv[31:0]});

   wire [63:0] ebd5a_t3vwkpflq = 
             
                 (pdw2zx8bnrucv | (bwqs5m4om61 & (~hbc9h8mi5tp))) ? (vrh7fcmgexv ? {32'h7FFF_FFFF,32'hFFFF_FFFF} : a5ju5vvapnv ? {32'h0000_0000,32'h7FFF_FFFF} : {32'hFFFF_FFFF,32'hFFFF_FFFF}) :
             
                 (bwqs5m4om61 & hbc9h8mi5tp) ? (vrh7fcmgexv ? {32'h8000_0000, 32'h0000_0000} : a5ju5vvapnv ? {32'hFFFF_FFFF,32'h8000_0000} : {32'h0000_0000,32'h0000_0000}) :
                 (a5ju5vvapnv | vrh7fcmgexv) ? hhqjnbrw2zq : lii58p0oecj8xmc3;

   
   
   
   wire t3xiz869kmsi_3wq = 
             
                 (pdw2zx8bnrucv | bwqs5m4om61) ? 1'b1 :  
                  (a5ju5vvapnv | vrh7fcmgexv) ? (cbmn5rtjbb68qbo | mojy8yz4lgbnb2vi) : (llz0g84mdu21zmq | ulou78bd89d6sgy);
   
   wire j6j8pa8aj_ipbu = 1'b0;
   
   
   wire wpx5ds4kagcnzl = 1'b0;
   
   
   wire x_gkjtpzcoygb_z = 1'b0;
   
   
   wire nhxsrct55nx7mr75b = (ia7awt7a85f2x8zfe | mjc2ko9ue08hnfniz8 | v6p6tk4wn1g_mj7) & (~t3xiz869kmsi_3wq);

   wire [4:0] y2wm4k1yrm37sbpjdf7u = {nhxsrct55nx7mr75b, wpx5ds4kagcnzl, x_gkjtpzcoygb_z, j6j8pa8aj_ipbu, t3xiz869kmsi_3wq};









  wire yr81i0s2 = af8gggx2rbk5w | im1jxeoei8g;
  wire rh_iqvuelzm = cix9qipqelc7k | u9bwc77pa3;
  wire bgx1o9epb0 = wpio23m13to3o0 | k937n2wbqgq;
  wire [63:0] mxm8oqd2lxz6 = (rh_iqvuelzm | bgx1o9epb0) ? {ticq8ng,y4a7pqq0kkz} : {32'b0,y4a7pqq0kkz};
  wire c3r259f43o3z7v = ~(|mxm8oqd2lxz6);
  
  
  
  

   wire [63:0] l71gng_e70xlmju6i04j = ~mxm8oqd2lxz6;
   wire [63:0] adolmfulsl08sg822k = 64'b0;
   wire        lvok_ngexfmtvo_hm407a = 1'b1; 

   wire        z45kmgu047lndnhmyt1 = af8gggx2rbk5w
                                   | z9ydb68fp_la3j
                                   | im1jxeoei8g
                                   | c2o9xduz06
                                   | cix9qipqelc7k
                                   | wpio23m13to3o0
                                   | u9bwc77pa3
                                   | k937n2wbqgq;

   wire [63:0] aglkl2uv0hawtn0uj = l71gng_e70xlmju6i04j + adolmfulsl08sg822k + lvok_ngexfmtvo_hm407a;

  wire w4dcqs0_8z8k = rh_iqvuelzm ? mxm8oqd2lxz6[63] : yr81i0s2 ? mxm8oqd2lxz6[31] : 1'b0;

  wire [63:0] mhfym4qmm = rh_iqvuelzm ? (w4dcqs0_8z8k ? aglkl2uv0hawtn0uj : mxm8oqd2lxz6) : yr81i0s2 ? (w4dcqs0_8z8k ? {32'b0,aglkl2uv0hawtn0uj[31:0]} : mxm8oqd2lxz6) : mxm8oqd2lxz6;


  wire [256-1:0] pf894p8faa = ({mhfym4qmm,{256-64{1'b0}}});
  wire [8-1:0] ht70;

  rwxldxdknfy97dlh i65hoqdmzb5rs8rl (
    .bjh (pf894p8faa),
    .ht70(ht70) 
  );

  wire [6-1:0] nwbg661y77_nqg = (rh_iqvuelzm | bgx1o9epb0) ? ht70[6-1:0] : {1'b0,ht70[5-1:0]};

  wire        e4_3ntz4xgj0u = af8gggx2rbk5w | z9ydb68fp_la3j | im1jxeoei8g | c2o9xduz06;
  wire        m70re9vay1 = cix9qipqelc7k | wpio23m13to3o0 | u9bwc77pa3 | k937n2wbqgq;
  wire        sb6nw06tetk = hr_5q_o87l78el0 | rau7b3otce5zq | pz73hz7q5h3oazsw | ieq_x45icc_ygmzwu;
  wire        g2r8zvzorupe187 = s4mabzvk_lget7 | ade81kyp0620xstvq | sn7ynh0j2u8h61 | uq85gpt70wdca;

  wire        xwxqw7_z001p = pz73hz7q5h3oazsw | ieq_x45icc_ygmzwu;
  wire        omvrz3vw7kq9t6 = sn7ynh0j2u8h61 | uq85gpt70wdca;
  wire        ugn5d14tezev = hr_5q_o87l78el0 | rau7b3otce5zq;
  wire        vc68wjfd30aavzk = s4mabzvk_lget7 | ade81kyp0620xstvq;

  wire jiv6seie_10do4 = cr7bv45kj7l & (e4_3ntz4xgj0u | m70re9vay1); 

  wire [6-1:0] ixcgnhvjijqxeuhp0;
  wire [64-1:0]bx1yhwlg4yqm;
  wire gx0lr2xgi7mj7;
  wire cm6nzdpeyik46rk;


  ux607_gnrl_dfflr #(6 )    rswmtt75dc4h41z0n9_xxz(jiv6seie_10do4, nwbg661y77_nqg, ixcgnhvjijqxeuhp0, gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(64)        ufj3iup33_yef0idg(jiv6seie_10do4, mhfym4qmm    , bx1yhwlg4yqm    , gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1 )      xjc06zu8ogj7e9ki8etu0771(jiv6seie_10do4, c3r259f43o3z7v  , gx0lr2xgi7mj7  , gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1 )      r2q7ugyr90rq1d507qklk(jiv6seie_10do4, w4dcqs0_8z8k  , cm6nzdpeyik46rk  , gf33atgy, ru_wi);

  wire [64-1:0] xm9fp5x8sdsgnnyv1vf = bx1yhwlg4yqm << ixcgnhvjijqxeuhp0;

  
  
  
  wire [10:0] xx70joqe2qlgyf6w = (omvrz3vw7kq9t6 ? 11'd1086 : 11'd1054)-{5'b0,ixcgnhvjijqxeuhp0};
  wire [ 7:0] y6sdjwxp0dt1h = (vc68wjfd30aavzk ? 8'd190 : 8'd158) -{2'b0,ixcgnhvjijqxeuhp0};

  wire [52:0] pe7gc9dqr37ph = omvrz3vw7kq9t6 ? xm9fp5x8sdsgnnyv1vf[63:11] : {xm9fp5x8sdsgnnyv1vf[31:0],21'b0};
  wire [23:0] usghctlpj2_46 = vc68wjfd30aavzk ? xm9fp5x8sdsgnnyv1vf[63:40] : xm9fp5x8sdsgnnyv1vf[31:8];

  wire sdqetqmk9q7fkv83ton;
  wire hho8ecwfuh3ja54mb    = omvrz3vw7kq9t6 ? pe7gc9dqr37ph[0] : usghctlpj2_46[0];
  wire hhtm0qxr0y3keri9in  = omvrz3vw7kq9t6 ? (xm9fp5x8sdsgnnyv1vf[10]) : vc68wjfd30aavzk ? (xm9fp5x8sdsgnnyv1vf[39]) : (xm9fp5x8sdsgnnyv1vf[7]);
  wire ed2aly5kzxxegumn  = omvrz3vw7kq9t6 ? (xm9fp5x8sdsgnnyv1vf[9]) : vc68wjfd30aavzk ? (xm9fp5x8sdsgnnyv1vf[38]) : (xm9fp5x8sdsgnnyv1vf[6]);
  wire gqyfq_havp408uqe = omvrz3vw7kq9t6 ? (|xm9fp5x8sdsgnnyv1vf[8:0]) : vc68wjfd30aavzk ? (|xm9fp5x8sdsgnnyv1vf[37:0]) : (|xm9fp5x8sdsgnnyv1vf[5:0]);

   el7n_zz16sk_ntvue9v a46sakzs911xk4 (
       .l      (hho8ecwfuh3ja54mb   ), 
       .g      (hhtm0qxr0y3keri9in ),
       .r      (ed2aly5kzxxegumn ),
       .s      (gqyfq_havp408uqe),
       .ly53de   (cm6nzdpeyik46rk),
       .nfj6b     (hr6uuvr3izh),
       .f6dc_rhcaz (sdqetqmk9q7fkv83ton) 
   );


  

  wire [63:0] owhmq9txebb2a9zyklrio9c_5 = omvrz3vw7kq9t6 ? {11'b0,pe7gc9dqr37ph} : {40'b0,usghctlpj2_46};
  wire [63:0] hfh_pcy6voxri913omng8m2a8ry0 = 64'b0;
  wire        j5tfly5h_wd6fmufafopdcm_ = sdqetqmk9q7fkv83ton;

  wire        spcrj9sis7u8esdkjajkdw6dcuv = sb6nw06tetk | g2r8zvzorupe187;

  wire [63:0] gsjuh3lhqf5dmqgse_tn8cemu = y4yutdej0620pote;
  wire [23:0] krh6hsdi49lxm = gsjuh3lhqf5dmqgse_tn8cemu[23:0];
  wire [52:0] g3sim70n20wxs1v = gsjuh3lhqf5dmqgse_tn8cemu[52:0];

  wire usou492tzhgqzjz9id = (&usghctlpj2_46[23:0]) & sdqetqmk9q7fkv83ton;
  wire ebqft_u7h83q6j_vz = (&pe7gc9dqr37ph[52:0]) & sdqetqmk9q7fkv83ton & omvrz3vw7kq9t6;

  wire [51:0] av94l5c_8l = ebqft_u7h83q6j_vz ? 52'b0 : omvrz3vw7kq9t6 ? g3sim70n20wxs1v[51:0] : pe7gc9dqr37ph[51:0];
  wire [22:0] lue2hslc3l4 = usou492tzhgqzjz9id ? 23'b0 : krh6hsdi49lxm[22:0];

  wire [10:0] idi7c9rdnli = ebqft_u7h83q6j_vz ? (xx70joqe2qlgyf6w + 1'b1) : xx70joqe2qlgyf6w;
  wire [ 7:0] st3z3s0rmosj4j = usou492tzhgqzjz9id ? (y6sdjwxp0dt1h + 1'b1) : y6sdjwxp0dt1h;

  wire [63:0] fhki71q1i = gx0lr2xgi7mj7 ? 64'b0 : {cm6nzdpeyik46rk,idi7c9rdnli,av94l5c_8l};
  wire [31:0] xrbruzney = gx0lr2xgi7mj7 ? 32'b0 : {cm6nzdpeyik46rk,st3z3s0rmosj4j,lue2hslc3l4};
   
   
   wire ykljt3ahha7e8mr2bsm0 = 1'b0;
   
   wire whcjgpc8x7reawnr1ak1o7 = 1'b0;
   
   wire b0m008ias_3_joo8ci = 1'b0;
   
   wire gtb7y9epksp_u7zqlj6u = 1'b0;
   
   wire ouakyql0g9e8sffn9ixyl = (xwxqw7_z001p ? 1'b0 : (hhtm0qxr0y3keri9in | ed2aly5kzxxegumn | gqyfq_havp408uqe)) | b0m008ias_3_joo8ci | gtb7y9epksp_u7zqlj6u;

   wire [4:0] f1flggli7x7mi5jwt9g10 = {ouakyql0g9e8sffn9ixyl, b0m008ias_3_joo8ci, gtb7y9epksp_u7zqlj6u, whcjgpc8x7reawnr1ak1o7, ykljt3ahha7e8mr2bsm0};









  wire vehdhv49gt6d2bj = cr7bv45kj7l & goy441jl;
  wire [ 7:0]  kvi4z7us5isov0a;
  wire [22:0]  dgudaduac_a7a;
  ux607_gnrl_dfflr #(8 ) q056qhvyf9x3hqvfu7e(vehdhv49gt6d2bj, dbw_bap_jqyl, kvi4z7us5isov0a, gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(23) xjwiwos4mhxqfn4qa(vehdhv49gt6d2bj, lkish79hpt, dgudaduac_a7a, gf33atgy, ru_wi);






  wire [10:0] ihvmf65uugl2ewbqg =  {3'b0,kvi4z7us5isov0a} + 11'd896; 
  wire [51:0] wqa5mpk3z64lvozs2q =  {dgudaduac_a7a,29'b0};
  wire [63:0] qhev__b7kylzel29z9w7f9 = {hbc9h8mi5tp,ihvmf65uugl2ewbqg,wqa5mpk3z64lvozs2q};



  wire [256-1:0] xyaajbvliil3bn2mr6 = ({1'b0,dgudaduac_a7a,{256-24{1'b0}}});
  wire [7:0] ftt0vhrwgob0c82_nc3ey;
  wire [5-1:0] ukt_g2cm_gifq9;

  rwxldxdknfy97dlh pnxhdxlxwdrqez3ci890d65nj (
    .bjh (xyaajbvliil3bn2mr6),
    .ht70(ftt0vhrwgob0c82_nc3ey) 
  );

  assign ukt_g2cm_gifq9 = ftt0vhrwgob0c82_nc3ey[5-1:0];

  wire [51:0] x57lprnbetqnwn4bkcv5;
  wire ui7e7chpi93voac2hm_dfzvyq;
  assign {ui7e7chpi93voac2hm_dfzvyq, x57lprnbetqnwn4bkcv5} =  {1'b0,dgudaduac_a7a,29'b0} << ukt_g2cm_gifq9;
  wire [10:0] y_u1ny5_14wq2rtwpqw83 = 11'd897 + (~{{6{1'b0}},ukt_g2cm_gifq9}) + 1'b1 ; 
  wire [63:0] f2yuodlbt822l1b6o2xm = {hbc9h8mi5tp,y_u1ny5_14wq2rtwpqw83,x57lprnbetqnwn4bkcv5};

  
  wire [63:0] pb1goy3hbcopmgu = 
                  ({64{z1iavptcuyb}} &   qhev__b7kylzel29z9w7f9) 
                | ({64{sjt2wedeei_gmt0}} & f2yuodlbt822l1b6o2xm) 
                | ({64{pdw2zx8bnrucv   }} & spdu2kgfxi4hwqf5 ) 
                | ({64{vnyuwuzda74sk9_   }} & l1gpd_rq1zeu6 ) 
                | ({64{se2fv2m60n1xym   }} & tm080y4ksbj0jwufg )  
                | ({64{l4tu2pzv06wzg   }} & uk4q4m8jvw0d8zp ) 
                | ({64{u75k9olcw2ovrh   }} & wzqga1virp_encj ); 

   
   wire a9fa29i9oppqitmjj = axgk4peda4gp;
   
   wire hq45kvlb4hjs381c663y3 = 1'b0;
   
   wire lvlpytojso100cxvhre_6 = 1'b0;
   
   wire zydjeq8gfzk97vrwqbmx = 1'b0;
   
   wire o4dov3p85cv36iopc6o = 1'b0;
   wire [4:0] eguplxhc_687urq5l0 = {o4dov3p85cv36iopc6o, lvlpytojso100cxvhre_6, zydjeq8gfzk97vrwqbmx, hq45kvlb4hjs381c663y3, a9fa29i9oppqitmjj};




















   wire [10:0]  hp9rd1eihd_z9;
   wire [10:0]  dd5hyb7iet0k8l;
   wire  dtzmrgu84s1mdscek9qo;
   wire  b5bbj3wjjezh0949e88y1;


   wire kqnn94hqa4r9;

   
   wire [11:0] sqpiekccxd2x4_ctvc2w0wi8 = {1'b0,vropxwawb};
   wire [11:0] i3slsg00pgw5vcpyqfv_3rxcw = (~(12'd896));
   wire        ha9di4e4z6dadblsh60250 = 1'b1;
   
   wire        ura_fvk48_k6iqthxf870q = ayc3vpo7;        
   assign      {dtzmrgu84s1mdscek9qo,hp9rd1eihd_z9} = mvpt9rw8vb52stdz38p[11:0];
   
   wire [11:0] y3cokke8yg3105dm4w_bbyy = 12'd896;
   wire [11:0] ueb1_pbdifwvfu3da_yito0e = (~{1'b0,vropxwawb});
   wire        dmuyykrx42nqxgusj55or = 1'b1;
   
   wire        lic9r65a3ssfzs_0n3gjmqu = ayc3vpo7;        
   assign      {b5bbj3wjjezh0949e88y1,dd5hyb7iet0k8l} = l1l1j1q86l7rjr2j[11:0];

 
   
   wire rgmk2oj9zacg0dcy4v_90k_= (&hp9rd1eihd_z9[7:0]);
   wire mnjeuoafst8sfo0jux3x= ~(|hp9rd1eihd_z9[7:0]);
   wire q4bt4op2nbaqlqxd2 = (~dtzmrgu84s1mdscek9qo) & ((|hp9rd1eihd_z9[10:8]) | rgmk2oj9zacg0dcy4v_90k_); 
   wire w7fmrmf7ghl938_mglbq_0 = dtzmrgu84s1mdscek9qo & (|dd5hyb7iet0k8l[10:5]);
 
   wire e1p_8oqyfr7t2qhap6 = (~dtzmrgu84s1mdscek9qo) & (~(|hp9rd1eihd_z9[10:8])) & (~rgmk2oj9zacg0dcy4v_90k_) & (~mnjeuoafst8sfo0jux3x);
 
   wire jga79_44n42d9bcjqf = (~(q4bt4op2nbaqlqxd2 | w7fmrmf7ghl938_mglbq_0 | e1p_8oqyfr7t2qhap6));
   wire rsp108bewnfhaswj_   = (~dtzmrgu84s1mdscek9qo) & (hp9rd1eihd_z9 == 11'd0);

   wire sxabvouyn80pvh;
   wire [23:0] q_o8yll2v1j49fdlm;
   wire m0wx272a4q0_zc2ww4w;
   wire xb2fgcgo_uwgc6jkf;
   wire [59:0] wns4jt3e4wkv0476ykwrf5k5b;
   wire f0de9y_8g8qmyn1k = |wns4jt3e4wkv0476ykwrf5k5b;

   
   
   
   wire omaxte58qmuedb = 
               ((vc529nuu == 3'b000) & 1'b1) 
              |((vc529nuu == 3'b011) & (~rhaf675bn)) 
              |((vc529nuu == 3'b010) & rhaf675bn)
              |((vc529nuu == 3'b001) & 1'b0)
              |((vc529nuu == 3'b100) & 1'b1);

   wire v7qlfzyd_lpbgae2ufm = (|xf92vp2m3d[26:0]);
   wire xvhmfh1tsn5foi6xea = (|xf92vp2m3d[52:27]);
   wire txiyqjrxqklqzoc = xvhmfh1tsn5foi6xea | v7qlfzyd_lpbgae2ufm;


   
   wire [180:0] n83bqbngxrxqxxo05_civdqb = {95'b0,xf92vp2m3d[52:0],33'b0};
   wire [  6:0] oup9k43j8btkzxiaite9 = {2'b0, dd5hyb7iet0k8l[4:0]};

   wire [180:0] gw0aqw1v_7ra026jbw3g9; 
   i6_4g5fspqlv1svn #(181) w7yt52pnla6jmoo93rklilolt(n83bqbngxrxqxxo05_civdqb, gw0aqw1v_7ra026jbw3g9);
   wire [  6:0] lj_r0gxh2jlgddmvmpdysrp = oup9k43j8btkzxiaite9;
   
   wire         p_ny_rf6klsay6sv = ayc3vpo7;           
   wire [180:0] pcgmvojsdhl5j7wtqek6 = joviasnyqgggsfacl;

   wire [180:0] b8zszqnll41ofx9dlmhg6mle;
   i6_4g5fspqlv1svn #(181) gyzuwmltjzi3fdsc8wwtidfwww(pcgmvojsdhl5j7wtqek6, b8zszqnll41ofx9dlmhg6mle);

   wire [ 85:0] oei3rxym1k6h = b8zszqnll41ofx9dlmhg6mle[85:0];

   assign {q_o8yll2v1j49fdlm, m0wx272a4q0_zc2ww4w, xb2fgcgo_uwgc6jkf, wns4jt3e4wkv0476ykwrf5k5b} =
                       
                 w7fmrmf7ghl938_mglbq_0 ? {26'b0,31'b0,txiyqjrxqklqzoc,28'b0} :
                       
                 (q4bt4op2nbaqlqxd2 & omaxte58qmuedb )? {  24'b0 ,1'b0,1'b0,32'b0,28'b0} :
                 (q4bt4op2nbaqlqxd2 & (~omaxte58qmuedb)) ? {(~24'b0),1'b0,1'b0,32'b0,28'b0} :
                       
                 e1p_8oqyfr7t2qhap6 ? {xf92vp2m3d[52:0], 5'b0,28'b0} :
                       
                       
                     
                     (oei3rxym1k6h >> 1'b1);


   el7n_zz16sk_ntvue9v nq0krmy09h3gmx (
       .l      (q_o8yll2v1j49fdlm[0]), 
       .g      (m0wx272a4q0_zc2ww4w),
       .r      (xb2fgcgo_uwgc6jkf),
       .s      (f0de9y_8g8qmyn1k),
       .ly53de   (mp3k_c3d),
       .nfj6b     (vc529nuu),
       .f6dc_rhcaz (sxabvouyn80pvh) 
   );

   wire [10:0] xki9rpxv59kysmzf2t;
   wire [23:0] mbpgpyw965o93zxcbedd ;
   wire qo4wnjwrpewhnsy      ;
   wire oldc8zjch_ivo2t4ivakjuj0w ;
   wire cq4p8wrizkn2w0muh9lz ;
   wire pkg9uh70m9r5qfr2br1krw    ;
   wire fnaj0ofqigt39ipd5_j    ;
   wire szk496rpt5gnjjwxw2    ;
   wire esm2i7auc4_ytlyxx96   ;
   wire mo_cnfk2_1t9m27pp6c2gft   ;
   wire d0l22goz68mi5gu0   ;
   wire h4vq176c1olpkhftm       ;

   assign kqnn94hqa4r9 = cr7bv45kj7l & ayc3vpo7;

  ux607_gnrl_dfflr #(11)     ymgr6lwk5ckagga3efs12ns4df(kqnn94hqa4r9, hp9rd1eihd_z9    , xki9rpxv59kysmzf2t    , gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(24)      gbo94lza8h27z7in98uprkcwv(kqnn94hqa4r9, q_o8yll2v1j49fdlm     , mbpgpyw965o93zxcbedd     , gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1 )      bvmylxvfxsv0uooqyp6xb(kqnn94hqa4r9, sxabvouyn80pvh     , qo4wnjwrpewhnsy     , gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1 ) xhjyismw0lz3mhnhsptppskw57d50x(kqnn94hqa4r9, w7fmrmf7ghl938_mglbq_0, oldc8zjch_ivo2t4ivakjuj0w, gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1 ) vfi5g2wjjw6mbnpv4tyu1npcdwp(kqnn94hqa4r9, q4bt4op2nbaqlqxd2, cq4p8wrizkn2w0muh9lz, gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1 )    b1pyt6sx2ifroxb211bkxxuyq(kqnn94hqa4r9, e1p_8oqyfr7t2qhap6   , pkg9uh70m9r5qfr2br1krw   , gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1 )    cq2j6j59d7m7vkzw95ie2bn(kqnn94hqa4r9, m0wx272a4q0_zc2ww4w   , fnaj0ofqigt39ipd5_j   , gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1 )    z1zsb4j7k7hbzai53vtjvkzeht1(kqnn94hqa4r9, xb2fgcgo_uwgc6jkf   , szk496rpt5gnjjwxw2   , gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1 )   h8pe7eu07c6hvzxvusnctuiutox(kqnn94hqa4r9, f0de9y_8g8qmyn1k  , esm2i7auc4_ytlyxx96  , gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1 )   z9iiakki7rqds970vle4hi01xk0(kqnn94hqa4r9, jga79_44n42d9bcjqf  , mo_cnfk2_1t9m27pp6c2gft  , gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1 )   fq7_u8nv88nbgqph5y5fsq5uqoz  (kqnn94hqa4r9, rsp108bewnfhaswj_    , d0l22goz68mi5gu0    , gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1 )   u3j0gbobv0_ihak2rqq91g0qu    (kqnn94hqa4r9, omaxte58qmuedb      , h4vq176c1olpkhftm      , gf33atgy, ru_wi);

  
  wire [63:0] lg0e3c0xtzym7r6qr3ldke = {40'b0,mbpgpyw965o93zxcbedd};
  wire [63:0] ibvdejo2hw6gfd5a53dhher4hoj = 64'b0;
  wire        igjyy7e1djo175nfpyefk6 = qo4wnjwrpewhnsy;

  wire        eg_gr5p9tp7d54mftb3ox2x = scjp5ckdygufd;

  wire [31:0] of0xk7mvylfujwckdmv1lfy3n = gflb0dmv454sowt17bx[31:0];
  wire [23:0] haga0vabnncrpfw3rkqn = of0xk7mvylfujwckdmv1lfy3n[23:0];

  wire ezi3qkvcv6hwxfrcflzte5oiob_unl;

  wire wgpbal5l2d098lnqyvz4ewn = (&mbpgpyw965o93zxcbedd[23:0]) & qo4wnjwrpewhnsy;

  wire [22:0] y27j95huqy27 = wgpbal5l2d098lnqyvz4ewn ? 23'b0 : haga0vabnncrpfw3rkqn[22:0];

  wire [ 7:0] zfff1e3chku1 = 
                       
                 oldc8zjch_ivo2t4ivakjuj0w ? 8'b0 :
                       
                 (cq4p8wrizkn2w0muh9lz & h4vq176c1olpkhftm )? 8'hFF : 
                 (cq4p8wrizkn2w0muh9lz & (~h4vq176c1olpkhftm)) ? 8'hFE : 
                       
                       
                 pkg9uh70m9r5qfr2br1krw ? (wgpbal5l2d098lnqyvz4ewn ? (xki9rpxv59kysmzf2t[7:0] + 1'b1) : xki9rpxv59kysmzf2t[7:0]) :
                       
                       ezi3qkvcv6hwxfrcflzte5oiob_unl ? 8'h1 : 8'h0;

  wire n74yqv89osk9_ljy9o8nywir = (~oldc8zjch_ivo2t4ivakjuj0w) & (~cq4p8wrizkn2w0muh9lz) 
                                & (pkg9uh70m9r5qfr2br1krw) 
                                & wgpbal5l2d098lnqyvz4ewn 
                                & (xki9rpxv59kysmzf2t == 11'hFE);

  assign ezi3qkvcv6hwxfrcflzte5oiob_unl = (~oldc8zjch_ivo2t4ivakjuj0w) & (~cq4p8wrizkn2w0muh9lz) & (~pkg9uh70m9r5qfr2br1krw) 
                                & (mo_cnfk2_1t9m27pp6c2gft) 
                                & qo4wnjwrpewhnsy  
                                & (mbpgpyw965o93zxcbedd == 24'h7F_FFFF) & d0l22goz68mi5gu0;

  wire [31:0] bf33foa4ntw0los =
  
                     
                 pdw2zx8bnrucv ? yalqc1omcjhx6 :
                     
                 vnyuwuzda74sk9_ ? t56x59ztjm5zwnj56 :
                 se2fv2m60n1xym ? vembz3jnjwpwx :
                     
                 l4tu2pzv06wzg ? d40417qihw6rqg :
                 u75k9olcw2ovrh ? ywnvnrprlg65x3uq : {hbc9h8mi5tp,zfff1e3chku1[7:0],y27j95huqy27};

   wire hq2a91udhq_o7gw56od9 = (pdw2zx8bnrucv | vnyuwuzda74sk9_ | se2fv2m60n1xym | l4tu2pzv06wzg | u75k9olcw2ovrh);
   
   wire ln95nxt09o6fqnio778 = axgk4peda4gp;
   
   wire zx3lu1stxlso4lsw3y_bc = 1'b0;
   
   
   wire kbqea1y9t9qqezy5fp = (~hq2a91udhq_o7gw56od9) & (oldc8zjch_ivo2t4ivakjuj0w | mo_cnfk2_1t9m27pp6c2gft) 
                          & (fnaj0ofqigt39ipd5_j | szk496rpt5gnjjwxw2 | esm2i7auc4_ytlyxx96);
   
        
   wire pm59oieq4ouggzsvl = (~hq2a91udhq_o7gw56od9) & (cq4p8wrizkn2w0muh9lz | n74yqv89osk9_ljy9o8nywir);
   
   wire h5owxrkl7pvby5psgobi7 = (~hq2a91udhq_o7gw56od9) & (fnaj0ofqigt39ipd5_j | szk496rpt5gnjjwxw2 | esm2i7auc4_ytlyxx96 | kbqea1y9t9qqezy5fp | pm59oieq4ouggzsvl);

   wire [4:0] mjge6k3zbamrbeai3d9 = {h5owxrkl7pvby5psgobi7, kbqea1y9t9qqezy5fp, pm59oieq4ouggzsvl, zx3lu1stxlso4lsw3y_bc, ln95nxt09o6fqnio778};







  assign uiwlxd =
        ({64{dmqidngg044lka0}} & ebd5a_t3vwkpflq) 
      | ({64{f4vcs6htny8xk9}} & ebd5a_t3vwkpflq)
      | ({64{hr_5q_o87l78el0}} & {32'hFFFF_FFFF,xrbruzney})
      | ({64{rau7b3otce5zq}} & {32'hFFFF_FFFF,xrbruzney})
      | ({64{dah1__e5zjv47wr}}& ebd5a_t3vwkpflq) 
      | ({64{zvw_q5tgix3s69c7o}}& ebd5a_t3vwkpflq)
      | ({64{s4mabzvk_lget7}}& {32'hFFFF_FFFF,xrbruzney})
      | ({64{ade81kyp0620xstvq}}& {32'hFFFF_FFFF,xrbruzney})
      | ({64{fj4nn1kh724bow}} & ebd5a_t3vwkpflq)
      | ({64{chfklna44pacjcho}} & ebd5a_t3vwkpflq)
      | ({64{pz73hz7q5h3oazsw}} & fhki71q1i)
      | ({64{ieq_x45icc_ygmzwu}} & fhki71q1i)
      | ({64{xurhhleqgmg8sy2}}& ebd5a_t3vwkpflq)
      | ({64{rpn9v9ketinrb4o7oj}}& ebd5a_t3vwkpflq)
      | ({64{sn7ynh0j2u8h61}}& fhki71q1i)
      | ({64{uq85gpt70wdca}}& fhki71q1i)
      | ({64{scjp5ckdygufd  }} & {32'hFFFF_FFFF,bf33foa4ntw0los})
      | ({64{kcx64rdtzypzm  }} & pb1goy3hbcopmgu) 
      ;

  wire [4:0] k6mvi11sj =
        ({5{dmqidngg044lka0}} & y2wm4k1yrm37sbpjdf7u)
      | ({5{f4vcs6htny8xk9}} & y2wm4k1yrm37sbpjdf7u)
      | ({5{hr_5q_o87l78el0}} & f1flggli7x7mi5jwt9g10)
      | ({5{rau7b3otce5zq}} & f1flggli7x7mi5jwt9g10)
      | ({5{dah1__e5zjv47wr}}& y2wm4k1yrm37sbpjdf7u)
      | ({5{zvw_q5tgix3s69c7o}}& y2wm4k1yrm37sbpjdf7u)
      | ({5{s4mabzvk_lget7}}& f1flggli7x7mi5jwt9g10)
      | ({5{ade81kyp0620xstvq}}& f1flggli7x7mi5jwt9g10)
      | ({5{fj4nn1kh724bow}} & y2wm4k1yrm37sbpjdf7u)
      | ({5{chfklna44pacjcho}} & y2wm4k1yrm37sbpjdf7u)
      | ({5{pz73hz7q5h3oazsw}} & f1flggli7x7mi5jwt9g10)
      | ({5{ieq_x45icc_ygmzwu}} & f1flggli7x7mi5jwt9g10)
      | ({5{xurhhleqgmg8sy2}}& y2wm4k1yrm37sbpjdf7u)
      | ({5{rpn9v9ketinrb4o7oj}}& y2wm4k1yrm37sbpjdf7u)
      | ({5{sn7ynh0j2u8h61}}& f1flggli7x7mi5jwt9g10)
      | ({5{uq85gpt70wdca}}& f1flggli7x7mi5jwt9g10)
      | ({5{scjp5ckdygufd  }} & mjge6k3zbamrbeai3d9)
      | ({5{kcx64rdtzypzm  }} & eguplxhc_687urq5l0)
      ;

  assign adnx9wgdt2 = {k6mvi11sj[0],k6mvi11sj[1],k6mvi11sj[2],k6mvi11sj[3],k6mvi11sj[4]}; 







   wire [180:0] p9c35mkpvg26ai1w062k; 
   wire [6:0]   oaeo91pwh63pd616dvkra; 
   
   assign { p9c35mkpvg26ai1w062k
          , oaeo91pwh63pd616dvkra} = 
              ({188{ejaudkhb58i42o3ci78 }} & 
                      {jkxd7ftbbh3xspajh
                      ,tzyyizq0dvvice8zgo5_n}
              ) |   
              ({188{p_ny_rf6klsay6sv }} & 
                      {gw0aqw1v_7ra026jbw3g9
                      ,lj_r0gxh2jlgddmvmpdysrp}
              ) ;   

   assign joviasnyqgggsfacl = p9c35mkpvg26ai1w062k << oaeo91pwh63pd616dvkra;


   wire [11:0] d9f8vcehnlpmw_oj7q; 
   wire [11:0] f8uvzururdrgxefwye; 
   wire        pco31x2lqnnejhzghke; 
   wire        osa_5u8ky1l89q9a; 

   wire [11:0] wm9pbpaf3izvyuh; 
   wire [11:0] p4m1e78vqg1kf0wx; 
   wire        dtdye51qcfpfm6spusw; 
   wire        k_ohwd25n61e250r7esc6; 

   assign {osa_5u8ky1l89q9a, mvpt9rw8vb52stdz38p} = d9f8vcehnlpmw_oj7q + f8uvzururdrgxefwye + pco31x2lqnnejhzghke;
   assign {k_ohwd25n61e250r7esc6, l1l1j1q86l7rjr2j} = wm9pbpaf3izvyuh + p4m1e78vqg1kf0wx + dtdye51qcfpfm6spusw;

   assign { d9f8vcehnlpmw_oj7q  
          , f8uvzururdrgxefwye  
          , pco31x2lqnnejhzghke} =
              ({25{i83vn2g75rui4ede6j9ioa70ugp }} & 
                      {xzraqync_3fsxk9k_3teii55y2
                      ,eb0ctt_nl3e3d7d1w_4p9n7x93
                      ,vc000h9sulun8dpbf0bz5fzxls}
              ) |   
              ({25{ura_fvk48_k6iqthxf870q}} & 
                      {sqpiekccxd2x4_ctvc2w0wi8
                      ,i3slsg00pgw5vcpyqfv_3rxcw
                      ,ha9di4e4z6dadblsh60250}
              ) ;   

   assign { wm9pbpaf3izvyuh  
          , p4m1e78vqg1kf0wx  
          , dtdye51qcfpfm6spusw} =
              ({25{amxnkuchi7l1_0kudwvt84gbi }} & 
                      {jdn4wx2w8tno0b61k_srrv
                      ,dslntpb2kksdjgkt0powur_
                      ,biyo66wdgpupq01jhemo3lq0}
              ) 
              |   ({25{lic9r65a3ssfzs_0n3gjmqu}} & 
                      {y3cokke8yg3105dm4w_bbyy
                      ,ueb1_pbdifwvfu3da_yito0e
                      ,dmuyykrx42nqxgusj55or}
              ) 
              ;   


   wire [63:0] r5pno8wfxkm303iiv; 
   wire [63:0] dwobwamcr_yq0u_v6p; 
   wire        sojgdhmnusto0fbz; 

   wire [63:0] o398vdz_cc_f542uvt; 
   wire [63:0] tykqrm68tpdpycge; 
   wire        iqftzud8t42tevt_l_8h; 

   assign {bb977ptd1fyw2vzt, y4yutdej0620pote} = r5pno8wfxkm303iiv + dwobwamcr_yq0u_v6p + sojgdhmnusto0fbz;
   assign {lgz5ovlgwou4qwx6k71sq, gflb0dmv454sowt17bx} = o398vdz_cc_f542uvt + tykqrm68tpdpycge + iqftzud8t42tevt_l_8h;

   assign { r5pno8wfxkm303iiv  
          , dwobwamcr_yq0u_v6p  
          , sojgdhmnusto0fbz} =
              ({129{z7zzynt4p6n91ltyfzw88yr }} & 
                      {mk5gl3ippdiih78z_h8_ngwbgpt
                      ,qaufsfnnc9i8ce5deb847cksm
                      ,mb8tn3wn2iqxl5a0jirs0h}
              ) |   
              ({129{spcrj9sis7u8esdkjajkdw6dcuv}} & 
                      {owhmq9txebb2a9zyklrio9c_5
                      ,hfh_pcy6voxri913omng8m2a8ry0
                      ,j5tfly5h_wd6fmufafopdcm_}
              ) ;   

   assign { o398vdz_cc_f542uvt  
          , tykqrm68tpdpycge  
          , iqftzud8t42tevt_l_8h} =
              ({129{bkz3ex8j6dty_vo9us5iq9r }} & 
                      {olk58do8mpdp18e6zbw2zzcwa
                      ,d4_gebt1q1dsvf_bvc3a0
                      ,c5381srmbn8numzwdtbkoy_9_4}
              ) 
              |   ({129{eg_gr5p9tp7d54mftb3ox2x}} & 
                      {lg0e3c0xtzym7r6qr3ldke
                      ,ibvdejo2hw6gfd5a53dhher4hoj
                      ,igjyy7e1djo175nfpyefk6}
              ) 
              ;   


endmodule























module avxgym1nr_i6e(
  
  
  input  yq7_jyt__u, 
  input  p1oz3zlyx9z099ko, 
  output i7xpott8rcin,
  input  [64-1:0] xfxtnu32e4,
  input  [64-1:0] bzyabkjyg5aufwj,
  input  [64-1:0] w_vtk6165e,
  input  [48-1:0]  nog5k2tkaj_,  
  input  [64-1:0] a1nhqrkfzavps,
  input  [4-1:0] p3g2fj0yq04eh,
  input  [3-1:0] k1hmos4y13oq40h,
  output hh9xkcr7e1fpzxae1ybn,

  
  input                             eg8yja9aryvtp8s,
  input  [64-1:0]           ti187a_zcpeoww6gv,
  input  [64-1:0]           zpr8r800wvts9w_mx,
  input  [64-1:0]           gv1t0hwgea_5zw0eibk,
  input  [64-1:0]           ccwkp0gpz76bmkrz,
  input  [48-1:0]  k8zoj8eu8lhoa3e82,  


  output q5h0basu9fqsocd,

  
  
  output bum_0_4oz7eoli40, 
  output i53j9zqmffz8y6oqz7t, 
  input  zt7k3255akax0ouek346m,
  output [64-1:0] vw3plvpp665o9dv9,
  output [64-1:0] bzyry2czkd6xk6zjhye,
  output [64-1:0] cp61fga88rjw8r82n3v,
  output [48-1:0]  je_9freaj3uhcgylh63_,  
  output [64-1:0] fqbjly2wnzhx63l,
  output [4-1:0] bzjarqiyu0mfd0z3p,
  output [3-1:0] v79ay3621ggo4h0d5aaj,
 
  
  
  
  output kf2dpoq324swtgxgs6p, 
  output l8kc7o3jpu34qr5q7, 
  input  zgtqckuiafu2aw2bjsy,
  output [64-1:0] sw6wc3aq6kk892q79y32,
  output [64-1:0] bgldh5yqcsal9_d,
  output [64-1:0] pflh54d0tzca0r8_,
  output [48-1:0]  rbuzk7rvhcg5f8qo25j,  
  output [64-1:0] k1d77g2k6dmwycm9z8,
  output [4-1:0] tkda6753pw4u9iq3ht,
  output [3-1:0] win4d4amp0pkd57fchc,

  
  
  output ywvgb6n56j5hgb2jrff, 
  output cbk5zw3f620wbbj1dvrxi, 
  input  kisnmwl5fk22ydrmv4,
  output [64-1:0] jf1prsiac8pb9waq4q,
  output [64-1:0] utnh02m2bfr89kp,
  output [64-1:0] nc5jui2ngra88qjivem,
  output [48-1:0]  pr309tdfjv528m400czp,  
  output [64-1:0] vchmkej8wq81b86w2qhu,
  output [4-1:0] i0d65n3vieh6ywu9yts,
  output [3-1:0] bucityy4pde4rrsrgrrqj,

  
  
  output ddc4jxtzijwcnfg, 
  output h_ur90x_3ax0srnyj, 
  input  dytkvkta2hudyfw07,
  input  mdk0j4bk2l0pmkz25px_h,
  output [64-1:0] xuixtwz82z81xfu02cgu,
  output [64-1:0] r1okty2iji67yzm9,
  output [64-1:0] keu9vxu53w1s5zr,
  output [48-1:0]  a0qgx1mu_gmlc7c6t5,  
  output [64-1:0] x0083y1q_m2c9h6,
  output [4-1:0] z94qawv75fwplf5ze90 

  );


  
  wire [2-1:0] o13hosud54289421  = nog5k2tkaj_ [6:5];

  wire oci0aoa9px8px = eg8yja9aryvtp8s; 
  wire cjj78pjxcu = (o13hosud54289421 == 2'd2); 
  wire ddr4_obijt7hd = (o13hosud54289421 == 2'd0); 
  wire bnjnczs_68_5tp = (o13hosud54289421 == 2'd3); 

  assign bum_0_4oz7eoli40 = yq7_jyt__u & oci0aoa9px8px & (~q5h0basu9fqsocd); 
  assign kf2dpoq324swtgxgs6p = yq7_jyt__u & cjj78pjxcu & (~q5h0basu9fqsocd); 
  assign ywvgb6n56j5hgb2jrff = yq7_jyt__u & bnjnczs_68_5tp & (~q5h0basu9fqsocd); 
  assign ddc4jxtzijwcnfg = yq7_jyt__u & ddr4_obijt7hd & (~mdk0j4bk2l0pmkz25px_h); 

  assign i53j9zqmffz8y6oqz7t = p1oz3zlyx9z099ko & oci0aoa9px8px;
  assign l8kc7o3jpu34qr5q7 = p1oz3zlyx9z099ko & cjj78pjxcu;
  assign cbk5zw3f620wbbj1dvrxi = p1oz3zlyx9z099ko & bnjnczs_68_5tp;
  assign h_ur90x_3ax0srnyj = p1oz3zlyx9z099ko & ddr4_obijt7hd;

  assign hh9xkcr7e1fpzxae1ybn = ~(
                            (q5h0basu9fqsocd & oci0aoa9px8px) 
                          | (q5h0basu9fqsocd & cjj78pjxcu) 
                          | (q5h0basu9fqsocd & bnjnczs_68_5tp) 
                          | (mdk0j4bk2l0pmkz25px_h & ddr4_obijt7hd)
                          ); 
  
  assign i7xpott8rcin     = (zt7k3255akax0ouek346m & oci0aoa9px8px) 
                          | (zgtqckuiafu2aw2bjsy & cjj78pjxcu) 
                          | (kisnmwl5fk22ydrmv4 & bnjnczs_68_5tp) 
                          | (dytkvkta2hudyfw07 & ddr4_obijt7hd); 
  
  wire [3-1:0] c6mh24qx7gmbl8cxpw  = eg8yja9aryvtp8s ? k8zoj8eu8lhoa3e82[9:7] : nog5k2tkaj_ [9:7];
  wire m7clc8vb7t9hcht7x         = (c6mh24qx7gmbl8cxpw == 3'b111);   
  wire [3-1:0] f3xyh1exzhxz394v   = m7clc8vb7t9hcht7x ? k1hmos4y13oq40h : c6mh24qx7gmbl8cxpw;
  
  
  
  assign q5h0basu9fqsocd    = 
                              (f3xyh1exzhxz394v == 3'b101)
                            | (f3xyh1exzhxz394v == 3'b110)
                            | (f3xyh1exzhxz394v == 3'b111);

  
  
  
  
  
  
  
  
  
  
  
  
  
             
             
             
  
             
  
             
  wire i1f2d0e21mc0d6jd209 = nog5k2tkaj_[19:19 ];
  wire t07ozrftfq49v1xpf = nog5k2tkaj_[20:20];
  wire p404nfi6aa16ixku3k1= nog5k2tkaj_[30:30 ];
  wire usxh0_qchzh4nshwu= nog5k2tkaj_[31:31];

  wire cuod7gqjnrbx7n_0p = nog5k2tkaj_[29:29];
  wire c7ttmuql_vy82  = nog5k2tkaj_[11:11 ];
  wire gig6pyl3lvde2tj = nog5k2tkaj_[12:12];
  wire ckylhcympzjnlf3 = nog5k2tkaj_[13:13];
  wire t59ya121g5qoi = nog5k2tkaj_[16:16];
  wire xuwi8b5_ahi4_o = nog5k2tkaj_[24:24 ];
  wire aiwxtk8ws0p11f = k8zoj8eu8lhoa3e82[23:23];
  wire x5e7sr5xdixajvq7ko = nog5k2tkaj_[13:13];

  wire gqw26qq65l0p9dw7ug     =  (oci0aoa9px8px & (~aiwxtk8ws0p11f))
                          | (cjj78pjxcu & (~x5e7sr5xdixajvq7ko)); 

  wire jujoq3mt3ztufhq7q2a  = bnjnczs_68_5tp & (~cuod7gqjnrbx7n_0p) & (c7ttmuql_vy82 | gig6pyl3lvde2tj | ckylhcympzjnlf3);

  wire hhxnr8xtx5u1ih9ph   = (bnjnczs_68_5tp & (i1f2d0e21mc0d6jd209 | t07ozrftfq49v1xpf)); 

  wire qvrj8r1frp_uaofspi7   = (bnjnczs_68_5tp & (p404nfi6aa16ixku3k1 | usxh0_qchzh4nshwu)); 

  wire mhm0lrcg4yd7ny = bnjnczs_68_5tp & t59ya121g5qoi &(~cuod7gqjnrbx7n_0p);

  wire b78fi3xv8fp_a = bnjnczs_68_5tp & xuwi8b5_ahi4_o &(~cuod7gqjnrbx7n_0p); 
 
  wire hrkl3eazhqtpgvtwlwdwf = gqw26qq65l0p9dw7ug | jujoq3mt3ztufhq7q2a | hhxnr8xtx5u1ih9ph | qvrj8r1frp_uaofspi7 | mhm0lrcg4yd7ny | b78fi3xv8fp_a;   

  wire vvci_dacs5h8pwa = hrkl3eazhqtpgvtwlwdwf & (~(&xfxtnu32e4[63:32]));
  wire hjlzvltivyqcgn = hrkl3eazhqtpgvtwlwdwf & (~(&bzyabkjyg5aufwj[63:32]));
  wire bqg0qzvhjlk = hrkl3eazhqtpgvtwlwdwf & (~(&w_vtk6165e[63:32]));
  wire [64-1:0] gxb7vkuoyr5ez5ytsp85xg = {32'hFFFF_FFFF,32'h7FC0_0000};
  wire [64-1:0] yvj78iqi3vkr191cwe3 = {32'hFFFF_FFFF,32'h7FC0_0000};
  wire [64-1:0] ai4k83ar37uryuo45kqiq = {32'hFFFF_FFFF,32'h7FC0_0000};
  wire [64-1:0] artnbioj = vvci_dacs5h8pwa ? gxb7vkuoyr5ez5ytsp85xg : xfxtnu32e4;
  wire [64-1:0] emfjxicm = hjlzvltivyqcgn ? yvj78iqi3vkr191cwe3 : bzyabkjyg5aufwj;
  wire [64-1:0] jtcy9rup = bqg0qzvhjlk ? ai4k83ar37uryuo45kqiq : w_vtk6165e;

  wire z09slkkjbcqyy93z = hrkl3eazhqtpgvtwlwdwf & (~(&ti187a_zcpeoww6gv[63:32]));
  wire eg3jrsaxae27l0e = hrkl3eazhqtpgvtwlwdwf & (~(&zpr8r800wvts9w_mx[63:32]));
  wire s1wv8zzbqf70q58_ = hrkl3eazhqtpgvtwlwdwf & (~(&gv1t0hwgea_5zw0eibk[63:32]));
  wire [64-1:0] evsynalol06cn5who0wrhtwj = {32'hFFFF_FFFF,32'h7FC0_0000};
  wire [64-1:0] h6sa95y1y8t676dg79_num = {32'hFFFF_FFFF,32'h7FC0_0000};
  wire [64-1:0] wtsymynctnf4dsnbb5ubfj2ix_v = {32'hFFFF_FFFF,32'h7FC0_0000};
  wire [64-1:0] wqcl9su8_9 = z09slkkjbcqyy93z ? evsynalol06cn5who0wrhtwj : ti187a_zcpeoww6gv;
  wire [64-1:0] h7r6ma08wi40 = eg3jrsaxae27l0e ? h6sa95y1y8t676dg79_num : zpr8r800wvts9w_mx;
  wire [64-1:0] bpwytpqr2n = s1wv8zzbqf70q58_ ? wtsymynctnf4dsnbb5ubfj2ix_v : gv1t0hwgea_5zw0eibk;


  
  assign vw3plvpp665o9dv9   = {64{oci0aoa9px8px}} & wqcl9su8_9[64-1:0];
  assign bzyry2czkd6xk6zjhye   = {64{oci0aoa9px8px}} & h7r6ma08wi40[64-1:0];
  assign cp61fga88rjw8r82n3v   = {64{oci0aoa9px8px}} & bpwytpqr2n[64-1:0];
  assign je_9freaj3uhcgylh63_  = {48{oci0aoa9px8px}} & k8zoj8eu8lhoa3e82;  
  assign fqbjly2wnzhx63l   = {64{oci0aoa9px8px}} & ccwkp0gpz76bmkrz;  
  assign bzjarqiyu0mfd0z3p  = {4{oci0aoa9px8px}} & p3g2fj0yq04eh;  
  assign v79ay3621ggo4h0d5aaj = {3{oci0aoa9px8px}} & f3xyh1exzhxz394v;  
  
  assign jf1prsiac8pb9waq4q   = {64{bnjnczs_68_5tp}} & artnbioj;
  assign utnh02m2bfr89kp   = {64{bnjnczs_68_5tp}} & emfjxicm;
  assign nc5jui2ngra88qjivem   = {64{bnjnczs_68_5tp}} & jtcy9rup;
  assign pr309tdfjv528m400czp  = {48{bnjnczs_68_5tp}} & nog5k2tkaj_;  
  assign vchmkej8wq81b86w2qhu   = {64{bnjnczs_68_5tp}} & a1nhqrkfzavps;  
  assign i0d65n3vieh6ywu9yts  = {4{bnjnczs_68_5tp}} & p3g2fj0yq04eh;  
  assign bucityy4pde4rrsrgrrqj = {3{bnjnczs_68_5tp}} & f3xyh1exzhxz394v;  
  
  assign sw6wc3aq6kk892q79y32   = {64{cjj78pjxcu}} & artnbioj[64-1:0];
  assign bgldh5yqcsal9_d   = {64{cjj78pjxcu}} & emfjxicm[64-1:0];
  assign pflh54d0tzca0r8_   = {64{cjj78pjxcu}} & jtcy9rup[64-1:0];
  assign rbuzk7rvhcg5f8qo25j  = {48{cjj78pjxcu}} & nog5k2tkaj_;  
  assign k1d77g2k6dmwycm9z8   = {64{cjj78pjxcu}} & a1nhqrkfzavps;  
  assign tkda6753pw4u9iq3ht  = {4{cjj78pjxcu}} & p3g2fj0yq04eh;  
  assign win4d4amp0pkd57fchc = {3{cjj78pjxcu}} & f3xyh1exzhxz394v;  
  
  assign xuixtwz82z81xfu02cgu   = {64{ddr4_obijt7hd}} & artnbioj[64-1:0];
  assign r1okty2iji67yzm9   = {64{ddr4_obijt7hd}} & emfjxicm[64-1:0];
  assign keu9vxu53w1s5zr   = {64{ddr4_obijt7hd}} & jtcy9rup[64-1:0];
  assign a0qgx1mu_gmlc7c6t5  = {48{ddr4_obijt7hd}} & nog5k2tkaj_;  
  assign x0083y1q_m2c9h6   = {64{ddr4_obijt7hd}} & a1nhqrkfzavps;  
  assign z94qawv75fwplf5ze90  = {4{ddr4_obijt7hd}} & p3g2fj0yq04eh;  

endmodule                                      






















module s4uzmkluo__rou46olor5a (
    input  [15:0] v2aj2jo,
    input  m10yxa5jl,

    output [64-1:0] uiwlxd,
    output [4:0] adnx9wgdt2

);

  
   wire [3-1:0] vc529nuu = 3'b001; 
  
   wire v0da13u6ykrw = (v2aj2jo[14:10] == 5'h1F);
   wire rg17tsy6wwx = (v2aj2jo[14:10] == 5'h00);
   wire wb75liyzd6vmew7 = (v2aj2jo[9:0] == 10'b0);
   wire bml43dgqbvm = rg17tsy6wwx & (~wb75liyzd6vmew7);
   wire ib3hkx1k0t = v2aj2jo[9];
   wire mgvwdehh1 = (~v0da13u6ykrw) & (~rg17tsy6wwx);
   wire aswm0l3tr55 = v0da13u6ykrw & (~wb75liyzd6vmew7) & (~ib3hkx1k0t);
   wire r41nzg = v0da13u6ykrw & (~wb75liyzd6vmew7) & ib3hkx1k0t;
   wire jqgto = r41nzg | aswm0l3tr55;
   wire ak6syfq = v0da13u6ykrw & wb75liyzd6vmew7;
   wire sy1qjmixh5e = (rg17tsy6wwx & wb75liyzd6vmew7);

   wire [ 9:0]  sfe6a4twd3cd = v2aj2jo[9:0];
   wire [ 4:0]  sq69mif63dg99 = v2aj2jo[14:10];
   wire         u1rd7n0pab = v2aj2jo[15];



   wire         mp3k_c3d = u1rd7n0pab;


   wire zpwosdnwv0 = ak6syfq & (~mp3k_c3d);
   wire h2pw9rtks0i = ak6syfq & mp3k_c3d;

   wire eqi5fiol = sy1qjmixh5e & (~mp3k_c3d);
   wire kc2obnf0fo = sy1qjmixh5e & mp3k_c3d;


   wire [32-1:0] e5otgqgjkm78gyd   = 32'h7FC00000;
   wire [16-1:0] rphhy7og5shc   = 16'h7E00;
   wire [32-1:0] lkpuz8x2a1y5   = 32'h7F800000;
   wire [16-1:0] wztskukp1m94m   = 16'h7C00;
   wire [32-1:0] w4m58zc6vxjqm   = 32'hFF800000;
   wire [16-1:0] os3en__39s   = 16'hFC00;
   wire [32-1:0] ppp30tohtvbsq   = 32'h00000000;
   wire [32-1:0] l2mifwazi5t_   = 32'h80000000;
   wire [16-1:0] c89mpiadrlqqb   = 16'h0000;
   wire [16-1:0] ged2mj90blbvit   = 16'h8000;
   wire [16-1:0] gz6qduuihnykm = 16'h7BFF;
   wire [16-1:0] s1th5gccdkngj = 16'hFBFF;













  wire [ 7:0] l05thqln33vhhqzuis =  {3'b0,sq69mif63dg99} + 8'd112; 
  wire [22:0] yhlqdyor8nfuccdf =  {sfe6a4twd3cd,13'b0};
  wire [31:0] r3udjcwxoemur9evh1j = {mp3k_c3d,l05thqln33vhhqzuis,yhlqdyor8nfuccdf};



  wire [256-1:0] nxmh4n8ce2t97t = ({1'b0,sfe6a4twd3cd,{256-11{1'b0}}});
  wire [7:0] t1c6_ahypwh7r;
  wire [4-1:0] um5umfozmuf0pe;

  rwxldxdknfy97dlh eya9fmk_n7n3e8f00xgpbpl (
    .bjh (nxmh4n8ce2t97t),
    .ht70(t1c6_ahypwh7r) 
  );

  assign um5umfozmuf0pe = t1c6_ahypwh7r[4-1:0];

  wire [22:0] p_govy3cw_xlgp8rv;
  wire kkepb15l85cjoik70gn;
  assign {kkepb15l85cjoik70gn, p_govy3cw_xlgp8rv} =  {1'b0,sfe6a4twd3cd,13'b0} << um5umfozmuf0pe;
  wire [ 7:0] qjwjqpc5mh_50mbncafo = 8'd113 + (~{{4{1'b0}},um5umfozmuf0pe}) + 1'b1 ; 
  wire [31:0] won_q7rfal4pajgg_r = {mp3k_c3d,qjwjqpc5mh_50mbncafo,p_govy3cw_xlgp8rv};

  
  wire [64-1:0] eif8v0b04 = 
                  ({64{mgvwdehh1    }} & {{32{r3udjcwxoemur9evh1j[31]}}  ,r3udjcwxoemur9evh1j}) 
                | ({64{bml43dgqbvm  }} & {{32{won_q7rfal4pajgg_r[31]}},won_q7rfal4pajgg_r}) 
                | ({64{jqgto     }} & {{32{e5otgqgjkm78gyd[31]}}      ,e5otgqgjkm78gyd} ) 
                | ({64{zpwosdnwv0   }} & {{32{lkpuz8x2a1y5[31]}}      ,lkpuz8x2a1y5} ) 
                | ({64{h2pw9rtks0i   }} & {{32{w4m58zc6vxjqm[31]}}      ,w4m58zc6vxjqm} )  
                | ({64{eqi5fiol   }} & {{32{ppp30tohtvbsq[31]}}      ,ppp30tohtvbsq} ) 
                | ({64{kc2obnf0fo   }} & {{32{l2mifwazi5t_[31]}}      ,l2mifwazi5t_} ); 
   
   
   
   
   wire ah_qis35wkxsqu = aswm0l3tr55;
   
   wire x42gpr4k4m8ef = 1'b0;
   
   wire rfzeewvlhzgm14k = 1'b0;
   
   wire ix_48__mqlfcey = 1'b0;
   
   wire yk2f_mtl5j5ydp = 1'b0;
   wire [4:0] rukged0k_aoegt_ro1f = {yk2f_mtl5j5ydp, rfzeewvlhzgm14k, ix_48__mqlfcey, x42gpr4k4m8ef, ah_qis35wkxsqu};








  assign uiwlxd = eif8v0b04;

  wire [4:0] k6mvi11sj = ({5{m10yxa5jl}} & rukged0k_aoegt_ro1f);

  assign adnx9wgdt2 = {k6mvi11sj[0],k6mvi11sj[1],k6mvi11sj[2],k6mvi11sj[3],k6mvi11sj[4]}; 

endmodule























module xpl5poo_wcl1vxzty7q #(
  parameter onr7l = 8 
)(
  input  [onr7l-1:0] ii,
  input  [onr7l-1:0] fij51v,
  input  [onr7l-1:0] cuzhl9,
  input           c,
  output [onr7l-1:0] s 
);

wire [onr7l-1:0] qk5ekvko5;
wire [onr7l-1:0] m01g6zl;

j3aa8h4yagvjsr416mg #(onr7l) r2oayxmv31tprr(
    .frgfco(ii  ),
    .ii(fij51v  ),
    .fij51v(cuzhl9  ),
    .c(qk5ekvko5), 
    .s(m01g6zl));

assign s = ({qk5ekvko5[onr7l-1:1],c} + m01g6zl);

endmodule


module m4df8f44pc8gto0crv(
  input  rj9pxiv3u3_pir,
  output b972jgf18d478vs1,
  input  [4-1:0] lw3kfp2bybej9,

  output ct0b7_gmchg9rz, 
  input  xvcpof07ihp69zc, 
  output [4 -1:0] bqcca4rpw2hdc6m1,

  output nyxl3jayn42b,
     output i0twiyq2wbmlvd6,
     output ql50zn__j2hmc8re,
     output ba0penccyqijkya4,

  output frfkcvpr3s1e,

  input gf33atgy,
  input ru_wi
);

  

  
  
  wire cns7w0cqkrz9uox; 
  wire jz8ky7a75l; 
  wire g1kx9xyy4gu1; 
  wire hkd5epsmvlz; 
  wire aubyyhgkel71; 
  wire ycwba7ldw34; 
  
  

  
  wire [4-1:0] x__lgcfoyn8;
  wire [4-1:0] taxi8w9ug_3ckl;
  wire [4-1:0] d2hhe5i9jn8;
  

  ux607_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(4)
  ) ay67o7ygpe34ch (
   .i_vld(rj9pxiv3u3_pir), 
   .i_rdy(b972jgf18d478vs1), 
   .i_dat(lw3kfp2bybej9),
   .o_vld(cns7w0cqkrz9uox), 
   .o_rdy(jz8ky7a75l), 
   .o_dat(x__lgcfoyn8),
 
   .clk  (gf33atgy  ),
   .rst_n(ru_wi)  
  );

  ux607_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(4)
  ) q4tuajzt5dbqj01qk6h (
   .i_vld(cns7w0cqkrz9uox), 
   .i_rdy(jz8ky7a75l), 
   .i_dat(x__lgcfoyn8),
   .o_vld(g1kx9xyy4gu1), 
   .o_rdy(hkd5epsmvlz), 
   .o_dat(taxi8w9ug_3ckl),
 
   .clk  (gf33atgy  ),
   .rst_n(ru_wi)  
  );

  ux607_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(4)
  ) ts657vjj488dibmw3 (
   .i_vld(g1kx9xyy4gu1), 
   .i_rdy(hkd5epsmvlz), 
   .i_dat(taxi8w9ug_3ckl),
   .o_vld(aubyyhgkel71), 
   .o_rdy(ycwba7ldw34), 
   .o_dat(d2hhe5i9jn8),
 
   .clk  (gf33atgy  ),
   .rst_n(ru_wi)  
  );


  
  
  
  

  
  
  
  
  assign nyxl3jayn42b = 1'b1;
  assign ycwba7ldw34 = xvcpof07ihp69zc;
  assign ct0b7_gmchg9rz = aubyyhgkel71;
  assign bqcca4rpw2hdc6m1 = d2hhe5i9jn8;
  assign i0twiyq2wbmlvd6 = rj9pxiv3u3_pir;
  assign ql50zn__j2hmc8re = cns7w0cqkrz9uox & jz8ky7a75l;
  assign ba0penccyqijkya4 = g1kx9xyy4gu1 & hkd5epsmvlz;
  assign frfkcvpr3s1e = cns7w0cqkrz9uox | g1kx9xyy4gu1 | aubyyhgkel71;

endmodule





module ggzvoy2zvu8ryca4ylw0(
  input [2:0] jq6ebmv,
  input [2:0] f7rj,
  output uriczc 
);

wire kqxmwtnmf = jq6ebmv[2] ^ f7rj[2];

wire x9ut0 =   jq6ebmv[1]  &   f7rj[1];
wire qzhlz = (~jq6ebmv[1]) & (~f7rj[1]);

wire z9k7hkt =   jq6ebmv[0]  &   f7rj[0];
wire bqaor4kps7 = (~jq6ebmv[0]) & (~f7rj[0]);

assign uriczc = (kqxmwtnmf & (
                        (x9ut0 & (~bqaor4kps7)) | 
                        (qzhlz & (~z9k7hkt))
                      )
            ) | 
           ((~kqxmwtnmf) & (
                          (qzhlz & (~bqaor4kps7)) | 
                          (x9ut0 & (~z9k7hkt))
                        )
           );

endmodule


module u6rhkw924ptxmc8p5wde #(
  parameter onr7l = 256 
)(
  input          a856yvdz,
  input [onr7l-1:0] bjh,
  input [7:0]    w40py,
  output[onr7l-1:0] adqhji 
);


wire[onr7l-1:0] x3vrpy = a856yvdz ? (~bjh) : bjh;

wire[onr7l-1:0] s4ir7c8hg=
		 {onr7l{w40py[1:0] == 2'b00}} & x3vrpy 
		|{onr7l{w40py[1:0] == 2'b01}} & {x3vrpy[onr7l-1-1:00],{1{a856yvdz}}}  
		|{onr7l{w40py[1:0] == 2'b10}} & {x3vrpy[onr7l-1-2:00],{2{a856yvdz}}}  
		|{onr7l{w40py[1:0] == 2'b11}} & {x3vrpy[onr7l-1-3:00],{3{a856yvdz}}} ;

wire[onr7l-1:0] lfpprd5dtfy=
		 {onr7l{w40py[3:2] == 2'b00}} & s4ir7c8hg 
		|{onr7l{w40py[3:2] == 2'b01}} & {s4ir7c8hg[onr7l-1-4:00] ,{4{a856yvdz}}}  
		|{onr7l{w40py[3:2] == 2'b10}} & {s4ir7c8hg[onr7l-1-8:00] ,{8{a856yvdz}}}  
		|{onr7l{w40py[3:2] == 2'b11}} & {s4ir7c8hg[onr7l-1-12:00],{12{a856yvdz}}} ;

wire[onr7l-1:0] cs8evrvizs=
		 {onr7l{w40py[5:4] == 2'b00}} & lfpprd5dtfy 
		|{onr7l{w40py[5:4] == 2'b01}} & {lfpprd5dtfy[onr7l-1-16:00],{16{a856yvdz}}}  
		|{onr7l{w40py[5:4] == 2'b10}} & {lfpprd5dtfy[onr7l-1-32:00],{32{a856yvdz}}}  
		|{onr7l{w40py[5:4] == 2'b11}} & {lfpprd5dtfy[onr7l-1-48:00],{48{a856yvdz}}} ;

wire[256-1:0] anl5941suw0xhcu;
generate
    if(onr7l > 192) begin: ukhn_zj0m74u_xu20f
      assign anl5941suw0xhcu =
		 {256{w40py[7:6] == 2'b00}} & {{256-onr7l{1'b0}},cs8evrvizs[onr7l-1:0]} 
		|{256{w40py[7:6] == 2'b01}} & {{256-onr7l{1'b0}},cs8evrvizs[onr7l-1-64:00],{64{a856yvdz}}}  
		|{256{w40py[7:6] == 2'b10}} & {{256-onr7l{1'b0}},cs8evrvizs[onr7l-1-128:00],{128{a856yvdz}}}  
		|{256{w40py[7:6] == 2'b11}} & {{256-onr7l{1'b0}},cs8evrvizs[onr7l-1-192:00],{192{a856yvdz}}} ;
    end
    else begin: l3rr903chra5y7
      assign anl5941suw0xhcu =
		 {256{w40py[7:6] == 2'b00}} & {{256-onr7l{1'b0}} ,cs8evrvizs[onr7l-1:0]} 
		|{256{w40py[7:6] == 2'b01}} & {{256-onr7l{1'b0}} ,cs8evrvizs[onr7l-1-64:00],{64{a856yvdz}}}  
		|{256{w40py[7:6] == 2'b10}} & {{256-onr7l{1'b0}} ,cs8evrvizs[onr7l-1-128:00],{128{a856yvdz}}}  
		|{256{w40py[7:6] == 2'b11}} & {{256-192{1'b0}},{192{a856yvdz}}} ;
    end
endgenerate

wire[onr7l-1:0] o6r0pl8eou = anl5941suw0xhcu[onr7l-1:0];

assign adqhji = o6r0pl8eou;

endmodule


module uwtp9d4cv1y3gqfa7u3jo #(
  parameter onr7l     = 256,
  parameter hw3qvr = 8
)(
  input [onr7l-1:0] bjh,
  output [hw3qvr-1:0] ht70
);

wire [onr7l-1:0] cvf2uttd2wy;

assign cvf2uttd2wy[onr7l-1] = bjh[onr7l-1];

genvar j;
generate 
 for (j=onr7l-2; j>=0; j=j-1) begin: m_j0ywdyf2
    assign cvf2uttd2wy[j] = (|bjh[onr7l-1:j]);
 end
endgenerate

wire [onr7l-1:0] i = cvf2uttd2wy & {1'b1,~cvf2uttd2wy[onr7l-1:1]};

assign ht70[0] = |{i[000], i[002], i[004], i[006], i[008], i[010], i[012], i[014], i[016], i[018],
                  i[020], i[022], i[024], i[026], i[028], i[030], i[032], i[034], i[036], i[038],
                  i[040], i[042], i[044], i[046], i[048], i[050], i[052], i[054], i[056], i[058],
                  i[060], i[062], i[064], i[066], i[068], i[070], i[072], i[074], i[076], i[078],
                  i[080], i[082], i[084], i[086], i[088], i[090], i[092], i[094], i[096], i[098],
                  i[100], i[102], i[104], i[106], i[108], i[110], i[112], i[114], i[116], i[118],
                  i[120], i[122], i[124], i[126], i[128], i[130], i[132], i[134], i[136], i[138],
                  i[140], i[142], i[144], i[146], i[148], i[150], i[152], i[154], i[156], i[158],
                  i[160], i[162], i[164], i[166], i[168], i[170], i[172], i[174], i[176], i[178],
                  i[180], i[182], i[184], i[186], i[188], i[190], i[192], i[194], i[196], i[198],
                  i[200], i[202], i[204], i[206], i[208], i[210], i[212], i[214], i[216], i[218],
                  i[220], i[222], i[224], i[226], i[228], i[230], i[232], i[234], i[236], i[238],
                  i[240], i[242], i[244], i[246], i[248], i[250], i[252], i[254]};

assign ht70[1] = |{i[000], i[001], i[004], i[005], i[008], i[009], i[012], i[013], 
                  i[016], i[017], i[020], i[021], i[024], i[025], i[028], i[029], 
                  i[032], i[033], i[036], i[037], i[040], i[041], i[044], i[045], 
                  i[048], i[049], i[052], i[053], i[056], i[057], i[060], i[061],
                  i[064], i[065], i[068], i[069], i[072], i[073], i[076], i[077],
                  i[080], i[081], i[084], i[085], i[088], i[089], i[092], i[093], 
                  i[096], i[097], i[100], i[101], i[104], i[105], i[108], i[109], 
                  i[112], i[113], i[116], i[117], i[120], i[121], i[124], i[125],
                  i[128], i[129], i[132], i[133], i[136], i[137], i[140], i[141],
                  i[144], i[145], i[148], i[149], i[152], i[153], i[156], i[157],
                  i[160], i[161], i[164], i[165], i[168], i[169], i[172], i[173],
                  i[176], i[177], i[180], i[181], i[184], i[185], i[188], i[189],
                  i[192], i[193], i[196], i[197], i[200], i[201], i[204], i[205],
                  i[208], i[209], i[212], i[213], i[216], i[217], i[220], i[221],
                  i[224], i[225], i[228], i[229], i[232], i[233], i[236], i[237],
                  i[240], i[241], i[244], i[245], i[248], i[249], i[252], i[253]};

assign ht70[2] = |{i[000], i[001], i[002], i[003], i[008], i[009], i[010], i[011], 
                  i[016], i[017], i[018], i[019], i[024], i[025], i[026], i[027], 
                  i[032], i[033], i[034], i[035], i[040], i[041], i[042], i[043], 
                  i[048], i[049], i[050], i[051], i[056], i[057], i[058], i[059],
                  i[064], i[065], i[066], i[067], i[072], i[073], i[074], i[075],
                  i[080], i[081], i[082], i[083], i[088], i[089], i[090], i[091], 
                  i[096], i[097], i[098], i[099], i[104], i[105], i[106], i[107], 
                  i[112], i[113], i[114], i[115], i[120], i[121], i[122], i[123],
                  i[128], i[129], i[130], i[131], i[136], i[137], i[138], i[139],
                  i[144], i[145], i[146], i[147], i[152], i[153], i[154], i[155],
                  i[160], i[161], i[162], i[163], i[168], i[169], i[170], i[171],
                  i[176], i[177], i[178], i[179], i[184], i[185], i[186], i[187],
                  i[192], i[193], i[194], i[195], i[200], i[201], i[202], i[203],
                  i[208], i[209], i[210], i[211], i[216], i[217], i[218], i[219],
                  i[224], i[225], i[226], i[227], i[232], i[233], i[234], i[235],
                  i[240], i[241], i[242], i[243], i[248], i[249], i[250], i[251]};

assign ht70[3] = |{i[000], i[001], i[002], i[003], i[004], i[005], i[006], i[007], 
                  i[016], i[017], i[018], i[019], i[020], i[021], i[022], i[023], 
                  i[032], i[033], i[034], i[035], i[036], i[037], i[038], i[039], 
                  i[048], i[049], i[050], i[051], i[052], i[053], i[054], i[055],
                  i[064], i[065], i[066], i[067], i[068], i[069], i[070], i[071],
                  i[080], i[081], i[082], i[083], i[084], i[085], i[086], i[087], 
                  i[096], i[097], i[098], i[099], i[100], i[101], i[102], i[103], 
                  i[112], i[113], i[114], i[115], i[116], i[117], i[118], i[119],
                  i[128], i[129], i[130], i[131], i[132], i[133], i[134], i[135],
                  i[144], i[145], i[146], i[147], i[148], i[149], i[150], i[151],
                  i[160], i[161], i[162], i[163], i[164], i[165], i[166], i[167],
                  i[176], i[177], i[178], i[179], i[180], i[181], i[182], i[183],
                  i[192], i[193], i[194], i[195], i[196], i[197], i[198], i[199],
                  i[208], i[209], i[210], i[211], i[212], i[213], i[214], i[215],
                  i[224], i[225], i[226], i[227], i[228], i[229], i[230], i[231],
                  i[240], i[241], i[242], i[243], i[244], i[245], i[246], i[247]};

assign ht70[4] = |{i[000], i[001], i[002], i[003], i[004], i[005], i[006], i[007], i[008], i[009], i[010], i[011], i[012], i[013], i[014], i[015], 
                  i[032], i[033], i[034], i[035], i[036], i[037], i[038], i[039], i[040], i[041], i[042], i[043], i[044], i[045], i[046], i[047], 
                  i[064], i[065], i[066], i[067], i[068], i[069], i[070], i[071], i[072], i[073], i[074], i[075], i[076], i[077], i[078], i[079],
                  i[096], i[097], i[098], i[099], i[100], i[101], i[102], i[103], i[104], i[105], i[106], i[107], i[108], i[109], i[110], i[111],
                  i[128], i[129], i[130], i[131], i[132], i[133], i[134], i[135], i[136], i[137], i[138], i[139], i[140], i[141], i[142], i[143],
                  i[160], i[161], i[162], i[163], i[164], i[165], i[166], i[167], i[168], i[169], i[170], i[171], i[172], i[173], i[174], i[175],
                  i[192], i[193], i[194], i[195], i[196], i[197], i[198], i[199], i[200], i[201], i[202], i[203], i[204], i[205], i[206], i[207],
                  i[224], i[225], i[226], i[227], i[228], i[229], i[230], i[231], i[232], i[233], i[234], i[235], i[236], i[237], i[238], i[239]};

assign ht70[5] = |{i[000], i[001], i[002], i[003], i[004], i[005], i[006], i[007], i[008], i[009], i[010], i[011], i[012], i[013], i[014], i[015], 
                  i[016], i[017], i[018], i[019], i[020], i[021], i[022], i[023], i[024], i[025], i[026], i[027], i[028], i[029], i[030], i[031],
                  i[064], i[065], i[066], i[067], i[068], i[069], i[070], i[071], i[072], i[073], i[074], i[075], i[076], i[077], i[078], i[079],
                  i[080], i[081], i[082], i[083], i[084], i[085], i[086], i[087], i[088], i[089], i[090], i[091], i[092], i[093], i[094], i[095],
                  i[128], i[129], i[130], i[131], i[132], i[133], i[134], i[135], i[136], i[137], i[138], i[139], i[140], i[141], i[142], i[143],
                  i[144], i[145], i[146], i[147], i[148], i[149], i[150], i[151], i[152], i[153], i[154], i[155], i[156], i[157], i[158], i[159], 
                  i[192], i[193], i[194], i[195], i[196], i[197], i[198], i[199], i[200], i[201], i[202], i[203], i[204], i[205], i[206], i[207],
                  i[208], i[209], i[210], i[211], i[212], i[213], i[214], i[215], i[216], i[217], i[218], i[219], i[220], i[221], i[222], i[223]};

assign ht70[6] = |{i[000], i[001], i[002], i[003], i[004], i[005], i[006], i[007], i[008], i[009], i[010], i[011], i[012], i[013], i[014], i[015], 
                  i[016], i[017], i[018], i[019], i[020], i[021], i[022], i[023], i[024], i[025], i[026], i[027], i[028], i[029], i[030], i[031],
                  i[032], i[033], i[034], i[035], i[036], i[037], i[038], i[039], i[040], i[041], i[042], i[043], i[044], i[045], i[046], i[047], 
                  i[048], i[049], i[050], i[051], i[052], i[053], i[054], i[055], i[056], i[057], i[058], i[059], i[060], i[061], i[062], i[063],
                  i[128], i[129], i[130], i[131], i[132], i[133], i[134], i[135], i[136], i[137], i[138], i[139], i[140], i[141], i[142], i[143],
	              i[144], i[145], i[146], i[147], i[148], i[149], i[150], i[151], i[152], i[153], i[154], i[155], i[156], i[157], i[158], i[159],
		          i[160], i[161], i[162], i[163], i[164], i[165], i[166], i[167], i[168], i[169], i[170], i[171], i[172], i[173], i[174], i[175],
		          i[176], i[177], i[178], i[179], i[180], i[181], i[182], i[183], i[184], i[185], i[186], i[187], i[188], i[189], i[190], i[191]};

assign ht70[7] = |{i[000], i[001], i[002], i[003], i[004], i[005], i[006], i[007], i[008], i[009], i[010], i[011], i[012], i[013], i[014], i[015], 
                  i[016], i[017], i[018], i[019], i[020], i[021], i[022], i[023], i[024], i[025], i[026], i[027], i[028], i[029], i[030], i[031],
                  i[032], i[033], i[034], i[035], i[036], i[037], i[038], i[039], i[040], i[041], i[042], i[043], i[044], i[045], i[046], i[047], 
                  i[048], i[049], i[050], i[051], i[052], i[053], i[054], i[055], i[056], i[057], i[058], i[059], i[060], i[061], i[062], i[063],
                  i[064], i[065], i[066], i[067], i[068], i[069], i[070], i[071], i[072], i[073], i[074], i[075], i[076], i[077], i[078], i[079],
                  i[080], i[081], i[082], i[083], i[084], i[085], i[086], i[087], i[088], i[089], i[090], i[091], i[092], i[093], i[094], i[095],
                  i[096], i[097], i[098], i[099], i[100], i[101], i[102], i[103], i[104], i[105], i[106], i[107], i[108], i[109], i[110], i[111],
                  i[112], i[113], i[114], i[115], i[116], i[117], i[118], i[119], i[120], i[121], i[122], i[123], i[124], i[125], i[126], i[127]}; 
endmodule

module yik149nqborvh6gofa51(
  
  input q_qkwqh5r,
  input clquq5nu,
  input ift60y9fnl2pw,
  input ktomwnwy0sxt8v,
  input [2:0] upi6iqvpb6svcz,
  input [63:0] zmjel5h70,
  input [63:0] lsgnmve7k1t,
  input [63:0] jj_j64pej,
  
  
  

  output [64-1:0]p0hjj76jp60rmlw, 
  output [4:0] bvdcuoqal71qlv60,
  output kv4pn5p7ocrk0,
  
  input  [64*2+5-1:0] m2k7jy,
  output [64*2+5-1:0] z2skz3wz,

  output i_mp1b_6j232kg,
  output bu481v83k29d,
  output asl_urmofi7s,
  output gh04xjbwykw9wd,
  output g4rmwbt0yslq,
  output p7fye2zf1aei,

  output wfoni28cogo3bhl,
  output rx_r34dltk5,
  output rux2i8zs5tg1l,
  output n2md11vbhgzi,
  output sslv1dv_v95mes2,
  output zu56_23__pyx62,
  
  output c597cob4z48yqld,
  output imknll0c6w2vjs,
  output clexjop8gcyt7i,
  output ug4q2r7d88wb9_,
  output ckzjjyyqsk_igo0q,
  output p23w6dm80pq0,
  
  input nyxl3jayn42b,
  input i0twiyq2wbmlvd6,
  input ql50zn__j2hmc8re,
  input ba0penccyqijkya4,

  input gf33atgy ,
  input ru_wi 
);


wire [31:0] fwknegmn = jj_j64pej[63:32];
wire [31:0] pu0_qq = jj_j64pej[31:00];
wire [31:0] ahdfbec41y = lsgnmve7k1t[63:32];
wire [31:0] b04cwa = lsgnmve7k1t[31:00];
wire [31:0] u49yq8sp = zmjel5h70[63:32];
wire [31:0] g91ks = zmjel5h70[31:0];


wire [5:0] qednpoi4d24hqegp;
assign bvdcuoqal71qlv60 = {qednpoi4d24hqegp[0],qednpoi4d24hqegp[1],qednpoi4d24hqegp[2],qednpoi4d24hqegp[3],qednpoi4d24hqegp[4]}; 

bh42kwltcb6jmjdg4k yo_63gowvnf2m3x9mw_o8d(
    .u49yq8sp                      (u49yq8sp                      ),
    .g91ks                      (g91ks                      ),
    .ahdfbec41y                      (ahdfbec41y                      ),
    .b04cwa                      (b04cwa                      ),
    .fwknegmn                      (fwknegmn                     ),
    .pu0_qq                      (pu0_qq                     ),
    .b1t_fvsbzg                  (q_qkwqh5r   ),
    .ift60y9fnl2pw               (ift60y9fnl2pw),
    .ktomwnwy0sxt8v               (ktomwnwy0sxt8v),
    .utngq               (clquq5nu               ),
                                                            
    .ncf9rmc                     (upi6iqvpb6svcz        ),
    .nyxl3jayn42b                (nyxl3jayn42b),
    .i0twiyq2wbmlvd6                (i0twiyq2wbmlvd6),
    .ql50zn__j2hmc8re                (ql50zn__j2hmc8re),
    .ba0penccyqijkya4                (ba0penccyqijkya4),
                                                            
    .g2gmxy0taet_c61t              (qednpoi4d24hqegp              ),
    .ynvgxkg9tf                  (p0hjj76jp60rmlw[31:0]),
    .ve6waju1kxdtbu                  (p0hjj76jp60rmlw[63:32]),
    .odq8ih2_pvx_6              (kv4pn5p7ocrk0),
    
    .m2k7jy                      (m2k7jy),
    .z2skz3wz                      (z2skz3wz),
    .i_mp1b_6j232kg                 (i_mp1b_6j232kg),
    .bu481v83k29d                 (bu481v83k29d),
    .asl_urmofi7s                 (asl_urmofi7s),
    .gh04xjbwykw9wd                 (gh04xjbwykw9wd),
    .g4rmwbt0yslq                 (g4rmwbt0yslq),
    .p7fye2zf1aei                 (p7fye2zf1aei),

    .wfoni28cogo3bhl                (wfoni28cogo3bhl),
    .rx_r34dltk5                (rx_r34dltk5),
    .rux2i8zs5tg1l                (rux2i8zs5tg1l),
    .n2md11vbhgzi                (n2md11vbhgzi),
    .sslv1dv_v95mes2                (sslv1dv_v95mes2),
    .zu56_23__pyx62                (zu56_23__pyx62),
  
    .c597cob4z48yqld                (c597cob4z48yqld),
    .imknll0c6w2vjs                (imknll0c6w2vjs),
    .clexjop8gcyt7i                (clexjop8gcyt7i),
    .ug4q2r7d88wb9_                (ug4q2r7d88wb9_),
    .ckzjjyyqsk_igo0q                (ckzjjyyqsk_igo0q),
    .p23w6dm80pq0                (p23w6dm80pq0),
  
    .gf33atgy                       (gf33atgy  ),
    .ru_wi                   (ru_wi ) 
) ;

endmodule

module bh42kwltcb6jmjdg4k(
    input [31:0] u49yq8sp ,
    input [31:0] g91ks ,

    input [31:0] ahdfbec41y ,
    input [31:0] b04cwa ,
    input [31:0] fwknegmn ,
    input [31:0] pu0_qq ,
    input utngq ,
    input ktomwnwy0sxt8v,
    input [2:0] ncf9rmc ,

    output [31:0] ve6waju1kxdtbu,
    output [31:0] ynvgxkg9tf,
    output [6-1:0] g2gmxy0taet_c61t ,
    output odq8ih2_pvx_6,



    input  [64*2+5-1:0] m2k7jy,
    output [64*2+5-1:0] z2skz3wz,
    output i_mp1b_6j232kg,
    output bu481v83k29d,
    output asl_urmofi7s,
    output gh04xjbwykw9wd,
    output g4rmwbt0yslq,
    output p7fye2zf1aei,

    output wfoni28cogo3bhl,
    output rx_r34dltk5,
    output rux2i8zs5tg1l,
    output n2md11vbhgzi,
    output sslv1dv_v95mes2,
    output zu56_23__pyx62,

    output c597cob4z48yqld,
    output imknll0c6w2vjs,
    output clexjop8gcyt7i,
    output ug4q2r7d88wb9_,
    output ckzjjyyqsk_igo0q,
    output p23w6dm80pq0,

    input nyxl3jayn42b,
    input i0twiyq2wbmlvd6,
    input ql50zn__j2hmc8re,
    input ba0penccyqijkya4,

    input b1t_fvsbzg,
    input ift60y9fnl2pw,
    input gf33atgy ,
    input ru_wi 
) ;


wire a3q6tl0i5iuy = nyxl3jayn42b ;
wire d0evt768bc = i0twiyq2wbmlvd6;
wire xpqt2l625a3 = 1'b1;
wire ywro5vq2yino = ql50zn__j2hmc8re;
wire e97gdk7jw4ev = ba0penccyqijkya4;
wire p1xybnd9a = 1'b1;

wire m7s5rkmh;
wire gma5v70c;
wire mb8pmo37pwn;
wire nftpir1zs;
wire wo1nm8zgf6;
wire mj9r0qdcj;

wire kp3n0pwlaqgh;
wire mjcsl_c3dwtdp6;
wire zk65zkc8xko9ebz_;
wire yai82tv8en1jptsp;
wire sbnvbrzm2242zu82;
wire pfrrs7z9swy5vf;

wire [2:0] dx22d5r9g2vd;
wire [2:0] dlv8z4devpq45;
wire [2:0] vnqm46gumvwx;
wire [2:0] rfxycz8syti7h;
wire [2:0] ach5cwxikdp;

wire [64*2+5-1:0] vr7175mt1g;
wire [64*2+5-1:0] t28xspeeyv;
wire [64*2+5-1:0] svl_gmw;
wire [64*2+5-1:0] yef02erc;
wire [64*2+5-1:0] myqiiy_cpkk;
wire [64*2+5-1:0] p9je8hjc;

wire [18-1:0] ygvkqdhr3wl;
wire [18-1:0] u5_4mgyu0a;
wire [18-1:0] s7nm7w5ep2a;
wire [18-1:0] a28ll7e7x;
wire [18-1:0] tsz7elf8cv;
wire [18-1:0] m_qz0i0513;

wire t8nr0xyjm88kch7l;
wire ckwgdt4l67va;
wire t6bx6zcifoc03dk;
wire fv3vyybkh98eba;
wire auj_3mt9a3wlbcyh;
wire g3ubkkn59kc;

wire fhqh1rdjxepeirvc1;
wire oxnijj3cb_5w;
wire ag79ahc9003tjfw;
wire hyp1jmmm6umhihlz;
wire e5g0gz5pr513gc;
wire iaoj1beeb4un1;

wire qxbi5ya_x3iyq;
wire ow9a1nk6tcubsc0;
wire zn79hxvf49003;
wire vur92j3awscoy3c;
wire clk6_twfdf0y;
wire l7t9rpi03xnwcm;

wire ks5rw5y1tx3;
wire kbjfvasuqsn4g;
wire ljz2siay0_;
wire d0z44bwpp5;
wire bop_ca3wk7;

wire tqert0u9oxp5tq2j7f;
wire dg4dhucjpo5xzo4_qpxw;
wire g3izwxx_mo1ghg7;
wire gc7v9_vi47psze_7640t;
wire j1l5j73k_gend8nlm;
wire hfzrr01xek2w6k6q8;
wire zh45pxgz_p2t5jp0u;
wire j_af3lmvq39fmm38;
wire vstyiobwn29fmatxc53;
wire l8dp94mozhdlxmr43;
wire x_vjfqyby9ywowiy2u3;

wire mnwum_pdiuo;
wire eu4746dfcv63;
wire uc1umghn15g19b;

wire yunzqdsnvu2whivp;
wire t5bfoq7ke3iipt_2;
wire p4n5_8jz95lf5a_;
wire sk_hgye1w_624w_;
wire m6wrb1i20poe2z7_wtnk;

wire aq_ibj5uwgvmvpubeu;
wire uzw0q1vxxy2cg;
wire dg5d0rszkwioqupp;
wire eoqybvzdtc5hh;
wire n75p3l63agiq3tuy;
wire dcd4ih54y76fim;
wire cfyrb77ier93zex;
wire bw5l8ov4grr29galln;
wire nunpqy34d5rby3u2c;
wire x7034mgujddxpm19suz;


wire[106-1:0] z7z1y_k7;
wire[106-1:0] sxo8i0fku66y;

wire[106-1:0] b_0ht;
wire[106-1:0] oazfr2ucb;
wire[106-1:0] p07jru;
wire[106-1:0] is4rk;
wire[106-1:0] h5w1j3;
wire[106-1:0] vs1z8;
wire[106-1:0] hk7neg5b6;
wire[106-1:0] x_5tn8w;
wire[106-1:0] xdzb4s0ejm;
wire[106-1:0] tr2ajiq;
wire[106-1:0] f0k2ir301f;
wire[106-1:0] n2fm6;
wire[106-1:0] cpkrdt;
wire[106-1:0] td137;
wire[106-1:0] kf_ejf;
wire[106-1:0] olreui;
wire[106-1:0] nh9i6q51r;
wire[106-1:0] zu59l2mmd;
wire[106-1:0] dtoeq;
wire[106-1:0] m5s6xnj;
wire[106-1:0] rzu745tt29;
wire[106-1:0] ca8pgl9;
wire[106-1:0] wqjzd4lir;
wire[106-1:0] aeeu2arrcv;
wire[106-1:0] aihp3cuom0;
wire[106-1:0] uucty;
wire[106-1:0] rwnza0fed;
wire[106-1:0] lfm5om4i85;

wire[106-1:0] zf2wuu6f;
wire[106-1:0] ipmcb4953;
wire[106-1:0] vje27h4vio;
wire[106-1:0] skablhb13q;
wire[106-1:0] cb_65dtz;
wire[106-1:0] mue2czm03;
wire[106-1:0] apzd3bocb0jlz;
wire[106-1:0] qsofrkqvi;
wire[106-1:0] tbqp2_p5b;
wire[106-1:0] vask7qpb;
wire[106-1:0] vkbk0udu;
wire[106-1:0] y9vjbgehnlld;
wire[106-1:0] snujns_17o;
wire[106-1:0] r49be1odf;
wire[106-1:0] fmmslemj9z9;
wire[106-1:0] tezkbiwpx10os;
wire[106-1:0] ezb1_13jolmi;
wire[106-1:0] vgfckvnmljw;
wire[106-1:0] ps3bgs1w;
wire[106-1:0] wbbij0elfpd;
wire[106-1:0] vm7box2gikw3;
wire[106-1:0] wxqo_7ac7g;
wire[106-1:0] ufo0585p;
wire[106-1:0] gyh98b_6jowgw;
wire[106-1:0] nqh156gtt8f;
wire[106-1:0] xjc8hz47unk4;
wire[106-1:0] crlqmi91i;
wire[106-1:0] xuugnk6md694i;

wire[106-1:0] fz5l6am6;
wire[106-1:0] fxx71cde0f;
wire[106-1:0] gizb4v58_bc;
wire[106-1:0] ydnoov3_7x;
wire[106-1:0] e9z05qhld0;
wire[106-1:0] uf8wgiec;
wire[106-1:0] sq4cj16ceo;
wire[106-1:0] dqlgpi77o;
wire[106-1:0] pw7_78ztt;
wire[106-1:0] k4g2t42mbrb;
wire[106-1:0] edqpyho0og;
wire[106-1:0] go2kpgsuttj;
wire[106-1:0] nc2dhbcdb26q;
wire[106-1:0] rcs83fuv1yxfs;

wire[106-1:0] at16xua1qxc;
wire[106-1:0] ai4n2ob_j7ocd;
wire[106-1:0] o0s11rb3;
wire[106-1:0] nzl699hjo;
wire[106-1:0] jqprtktb8qr8;
wire[106-1:0] frs3fk930avn;
wire[106-1:0] pk0153efgrg0;
wire[106-1:0] cpq3wxamh6ly;

wire[106-1:0] kaxkamth;
wire[106-1:0] vou_g00czb2;
wire[106-1:0] rbm2min6;
wire[106-1:0] qtui513wjhfz;

wire[106-1:0] mknydvsmn87;
wire[106-1:0] ga_yvggsogewp;
wire[106-1:0] z49e6oo_eurd;
wire[106-1:0] ttw8izs6;

wire e7hmnv0h1u8kjcw = (~kp3n0pwlaqgh) & a3q6tl0i5iuy;
wire enaanseli0es1 = (~mjcsl_c3dwtdp6) & d0evt768bc;
wire f4_3ig0unyv0i = (~zk65zkc8xko9ebz_) & xpqt2l625a3;
wire iue_ys441x03e_7n = (~yai82tv8en1jptsp) & ywro5vq2yino;
wire k5oz5augg717tkto = (~sbnvbrzm2242zu82) & e97gdk7jw4ev;
wire w9i0xdvu4_amoafu = (~pfrrs7z9swy5vf) & p1xybnd9a;

wire imq1k9bcch57k6w = utngq    ? kp3n0pwlaqgh :1'b0;
wire xocqwg27spn = m7s5rkmh ? mjcsl_c3dwtdp6 :1'b0;
wire zhppkn5dtqw = gma5v70c ? zk65zkc8xko9ebz_ :1'b0;
wire hlou4w_6e93mojh = mb8pmo37pwn ? yai82tv8en1jptsp :1'b0;
wire bi_6lyh1go = nftpir1zs ? sbnvbrzm2242zu82 :1'b0;
wire vaovag0tfaw2r = wo1nm8zgf6 ? pfrrs7z9swy5vf :1'b0;

wire qkv0nlfisqqas0 = kp3n0pwlaqgh;
wire stbn1nqzc00f = mjcsl_c3dwtdp6;
wire ybp58h03sal_ = zk65zkc8xko9ebz_;
wire hkc58ciovfj8f = yai82tv8en1jptsp;
wire iu4_c773tsqx = sbnvbrzm2242zu82;
wire o6xo7iacb14nta9 = pfrrs7z9swy5vf;

wire j04tei231k0topjtp = imq1k9bcch57k6w & a3q6tl0i5iuy;
wire qcxfzz_taf0uuvgpi = xocqwg27spn & d0evt768bc;
wire iefflu1iikpd9jjc = zhppkn5dtqw & xpqt2l625a3;
wire cv8vshys52pxuhd0n = hlou4w_6e93mojh & ywro5vq2yino;
wire apgiwgv4bubvui1j = bi_6lyh1go & e97gdk7jw4ev;
wire obkyh6cqeeh_i = vaovag0tfaw2r & p1xybnd9a;

wire g5jlqz0uszu2tl2 = qkv0nlfisqqas0 & a3q6tl0i5iuy;
wire x97f4cgxzyq9tb = stbn1nqzc00f & d0evt768bc;
wire r1555lotjfob = ybp58h03sal_ & xpqt2l625a3;
wire vsd4e757l2_bb = hkc58ciovfj8f & ywro5vq2yino;
wire mnchfusd_pal_g = iu4_c773tsqx & e97gdk7jw4ev;
wire lvibl7p2cgbe71k = o6xo7iacb14nta9 & p1xybnd9a;

assign ygvkqdhr3wl = {
                          t8nr0xyjm88kch7l,
                          ckwgdt4l67va,
                          t6bx6zcifoc03dk,
                          fv3vyybkh98eba,
                          auj_3mt9a3wlbcyh,
                          g3ubkkn59kc, 
                          fhqh1rdjxepeirvc1,
                          oxnijj3cb_5w,
                          ag79ahc9003tjfw,
                          hyp1jmmm6umhihlz,
                          e5g0gz5pr513gc,
                          iaoj1beeb4un1, 
                          qxbi5ya_x3iyq,
                          ow9a1nk6tcubsc0,
                          zn79hxvf49003,
                          vur92j3awscoy3c,
                          clk6_twfdf0y,
                          l7t9rpi03xnwcm 
                        };


assign {
                          i_mp1b_6j232kg,
                          bu481v83k29d,
                          asl_urmofi7s,
                          gh04xjbwykw9wd,
                          g4rmwbt0yslq,
                          p7fye2zf1aei,
                          wfoni28cogo3bhl,
                          rx_r34dltk5,
                          rux2i8zs5tg1l,
                          n2md11vbhgzi,
                          sslv1dv_v95mes2,
                          zu56_23__pyx62, 
                          c597cob4z48yqld,
                          imknll0c6w2vjs,
                          clexjop8gcyt7i,
                          ug4q2r7d88wb9_,
                          ckzjjyyqsk_igo0q,
                          p23w6dm80pq0 
                        } = m_qz0i0513;

assign z2skz3wz = p9je8hjc;
wire el96tsan45rrpod0r = utngq ? ((u49yq8sp[31] ^ ahdfbec41y[31]) ^ ktomwnwy0sxt8v) : ((g91ks[31] ^ b04cwa[31]) ^ ktomwnwy0sxt8v);
wire w628i27t5rsmxho = utngq ? (fwknegmn[31] ^ ift60y9fnl2pw) : (pu0_qq[31] ^ ift60y9fnl2pw);
wire jlx9c2o3yzo  = (el96tsan45rrpod0r ^ w628i27t5rsmxho);


wire [7-1:0] z5377lopdyjs6g;
wire [31:0] a52vuclb86uofcv7qqc;
wire [31:0] vra8744pgx17_zwuy6;


wire i48mlnnyzur = utngq ? (u49yq8sp[30:20] == 11'h000)      : (g91ks[30:23] == 8'h00);
wire td1glnmfo2 = utngq ? (ahdfbec41y[30:20] == 11'h000)      : (b04cwa[30:23] == 8'h00);
wire fut03jb6c4 = utngq ? (fwknegmn[30:20] == 11'h000)      : (pu0_qq[30:23] == 8'h00);
wire m23r0kqbby  = utngq ? ({fwknegmn[19:0],pu0_qq} == 52'b0) : (pu0_qq[22:0] == 23'b0);

assign mnwum_pdiuo = i48mlnnyzur;
assign eu4746dfcv63 = td1glnmfo2;
assign uc1umghn15g19b = fut03jb6c4 & ~m23r0kqbby;


wire wijmhrmp5iul;
wire cz7maz0fnx72thc;

b6d95x1xv7_zr3t2ebk sx7r9qgwm5ludj_2o(
    .hfzrr01xek2w6k6q8            (hfzrr01xek2w6k6q8),
    .uaeb8t1ovp              (zh45pxgz_p2t5jp0u),
    .y18h0qaenz              (j_af3lmvq39fmm38),
    .tqert0u9oxp5tq2j7f         (tqert0u9oxp5tq2j7f),
    .dg4dhucjpo5xzo4_qpxw         (dg4dhucjpo5xzo4_qpxw),
    .u49yq8sp                    (u49yq8sp),
    .g91ks                    (g91ks),
    .ahdfbec41y                    (ahdfbec41y),
    .b04cwa                    (b04cwa),
    .fwknegmn                    (fwknegmn),
    .pu0_qq                    (pu0_qq),
    .dx22d5r9g2vd               (dx22d5r9g2vd),
    .utngq             (utngq    ),
    .m7s5rkmh         (m7s5rkmh),
    .gma5v70c         (gma5v70c),
    .nxirove5d1                (wijmhrmp5iul   ),
    .oxto21kj774l      (cz7maz0fnx72thc),
    .acl1oms948eb26          (vra8744pgx17_zwuy6),
    .t0wz63jpdmeq4e          (a52vuclb86uofcv7qqc),
    .gzvyqzlwpz            (z5377lopdyjs6g),
    .kxfk1t4l2_39m7a7            (e7hmnv0h1u8kjcw),
    .su7v8qw44q19            (x97f4cgxzyq9tb),
    .t8nr0xyjm88kch7l             (t8nr0xyjm88kch7l),
    .ckwgdt4l67va             (ckwgdt4l67va),
    .t6bx6zcifoc03dk             (t6bx6zcifoc03dk),
    .fv3vyybkh98eba             (fv3vyybkh98eba),
    .auj_3mt9a3wlbcyh             (auj_3mt9a3wlbcyh),
    .g3ubkkn59kc             (g3ubkkn59kc),
    .fhqh1rdjxepeirvc1            (fhqh1rdjxepeirvc1),
    .oxnijj3cb_5w            (oxnijj3cb_5w),
    .ag79ahc9003tjfw            (ag79ahc9003tjfw),
    .hyp1jmmm6umhihlz            (hyp1jmmm6umhihlz),
    .e5g0gz5pr513gc            (e5g0gz5pr513gc),
    .iaoj1beeb4un1            (iaoj1beeb4un1),
    .qxbi5ya_x3iyq            (qxbi5ya_x3iyq),
    .ow9a1nk6tcubsc0            (ow9a1nk6tcubsc0),
    .zn79hxvf49003            (zn79hxvf49003),
    .vur92j3awscoy3c            (vur92j3awscoy3c),
    .clk6_twfdf0y            (clk6_twfdf0y),
    .l7t9rpi03xnwcm            (l7t9rpi03xnwcm),
    .ru_wi                 (ru_wi),
    .gf33atgy                     (gf33atgy)
);


assign kp3n0pwlaqgh = 1'b0;
assign mjcsl_c3dwtdp6 = cz7maz0fnx72thc;
assign zk65zkc8xko9ebz_ = kbjfvasuqsn4g;
assign yai82tv8en1jptsp = ljz2siay0_;
assign sbnvbrzm2242zu82 = d0z44bwpp5;
assign pfrrs7z9swy5vf = bop_ca3wk7;


wire[31:0] s6102_hpsio4ve;
wire[31:0] u5gxirwoddu54_;
wire[31:0] pfbn0r50hqi;
wire[31:0] a_vhiehymx7da1hco = vra8744pgx17_zwuy6;
wire[31:0] bn7gxjodtjqv9q5qd = s6102_hpsio4ve;
wire[31:0] k4x1lk0_vv_0ki1gtj = u5gxirwoddu54_;

wire[31:0] bcw8lurc42z;
wire[31:0] xgs6vgfhby7;
wire[31:0] fjo4qiwyjs8;
wire[31:0] wdskaz5d6p9ismr1j = gma5v70c ? a52vuclb86uofcv7qqc :32'b0;
wire[31:0] qqbg0l90wg42et = bcw8lurc42z;
wire[31:0] qz1zeyajzdmhr5vv6 = xgs6vgfhby7;
                       
wire[7-1:0] z80wawc634pnw8u;
wire[7-1:0] xqjlst8d7p1gb;
wire[7-1:0] gcl5p_j91agj;
wire[7-1:0] a5qzn5s78uj02pe = z5377lopdyjs6g;
wire[7-1:0] gj0mcve6t3a1peo = z80wawc634pnw8u;
wire[7-1:0] cv00o83d94urbkwcu = xqjlst8d7p1gb;

wire[11:0] zpl5t2pi8pm = utngq ? (mnwum_pdiuo ? 12'b1: {1'b0,u49yq8sp[30:20]}) :12'b0;
wire[11:0] y9qm_wv3pox4c1 = utngq ? (eu4746dfcv63 ? 12'b1: {1'b0,ahdfbec41y[30:20]}) :12'b0;
wire[11:0] q4n_ns9xf8f9z = utngq ? (uc1umghn15g19b ? 12'b1: {1'b0,fwknegmn[30:20]}) :12'b0;

wire[11:0] vnyip75m0u8z = (~utngq) ? (mnwum_pdiuo ? 12'b1: {4'b0,g91ks[30:23]}) :12'b0;
wire[11:0] ejb5jf8at329q8 = (~utngq) ? (eu4746dfcv63 ? 12'b1: {4'b0,b04cwa[30:23]}) :12'b0;
wire[11:0] whafz8l2nomw_0 = (~utngq) ? (uc1umghn15g19b ? 12'b1: {4'b0,pu0_qq[30:23]}) :12'b0;


wire[52:0] o94ohpc33fy_edaky = {53{utngq}}  & {~uc1umghn15g19b,fwknegmn[19:0],pu0_qq[31:0]};
wire[23:0] sw2iq_k_3ykq6l36 = {24{~utngq}} & {~uc1umghn15g19b, pu0_qq[22:0]};


wire vb_j3t59zgyb7r05r;
wire[12:0] duxpze1m6dlz2rx;
wire[12:0] crtsq13_r9b5_i8j;
wire[12:0] xrc71n3kb03z2;
wire b7x36_v4z0jlprnsb8vmn2;
wire[161-1:0] wfjl06kozsl7u3d95drhv8;
wire[74-1:0] gbyt7t2vj0c3ymg7p6dqxz;
wire fi2z120absus4g;

wire [12:0] v46v_ikm00k;
wire [12:0] pk01ktquuo1;
wire [12:0] mlgzk0dlchiy;

wire [12:0] not1kzp34m717_xrz3_;
wire [12:0] m4bd_iyv30v8ins0qb;

wire [12:0] u7v1l8233z7v63;
wire [12:0] vfz3yrokggbpc0b1b4;

wire [12:0] bv1krzrvrnk8hdr;
wire [12:0] ogkix3lj2m4hbon35a;
wire [12:0] c5g6edg75opsh985r;

wire [12:0] e8_x96sdkot60an7gl;
wire [12:0] k4weigq4ziemgtsb8c;

wire aed9k35_92eftqn4tu_nv;


wire [11:0] m69yhryw = utngq ? zpl5t2pi8pm : vnyip75m0u8z;
wire [11:0] rhd1sc8doent = utngq ? y9qm_wv3pox4c1 : ejb5jf8at329q8;
wire [11:0] zq3hfen = utngq ? q4n_ns9xf8f9z : whafz8l2nomw_0;


wire [12:0] vvtb10ccg215rrzm37t = vb_j3t59zgyb7r05r ? mlgzk0dlchiy : e8_x96sdkot60an7gl;

wire [12:0] u0owxonpqsp8  = m7s5rkmh ? 13'd967 : 13'd100;
wire [12:0] ntg11u8x4ichcr = m7s5rkmh ? 13'd968 : 13'd101;
wire [12:0] ya7uq7fuidy9 = m7s5rkmh ? 13'd970 : 13'd103;

xpl5poo_wcl1vxzty7q #(13) nt3lt6m53qdwz66yue(
    .ii (v46v_ikm00k), 
    .fij51v (pk01ktquuo1), 
    .cuzhl9 (~u0owxonpqsp8), 
    .c  (1'b1),
    .s  (e8_x96sdkot60an7gl)
);

xpl5poo_wcl1vxzty7q #(13) xqb_k4mgkbv_061( 
    .ii (v46v_ikm00k), 
    .fij51v (pk01ktquuo1),
    .cuzhl9 (~ntg11u8x4ichcr), 
    .c  (1'b1), 
    .s  (k4weigq4ziemgtsb8c)
);

xpl5poo_wcl1vxzty7q #(13) hjh3bjfmsdeqhve4g( 
    .ii (~v46v_ikm00k), 
    .fij51v (~pk01ktquuo1),
    .cuzhl9 (ya7uq7fuidy9),
    .c  (1'b0),
    .s  (bv1krzrvrnk8hdr)
);

wire [12:0] r6p8gd02fp8dbxt9j = mlgzk0dlchiy + 13'h1FFF;
wire [12:0] pa0vxwh5h1zrzt41cf     = vb_j3t59zgyb7r05r ? r6p8gd02fp8dbxt9j :
                                                 k4weigq4ziemgtsb8c[12] ? 13'b0 : k4weigq4ziemgtsb8c;


wire ri3iascff6a_jektfoqpz1b = (not1kzp34m717_xrz3_[12] | (not1kzp34m717_xrz3_ == 13'b0));

assign wfjl06kozsl7u3d95drhv8 = (
                             fi2z120absus4g ? (~{161'b0}) : 
                             (u7v1l8233z7v63[12:0] > 13'd160) ? 161'b0 :
                             ((~{161'b0}) >> u7v1l8233z7v63[7:0])
                           );

assign gbyt7t2vj0c3ymg7p6dqxz = fi2z120absus4g ? (~{74'b0}) :
                           (u7v1l8233z7v63[12:0] > 13'd73) ? 74'b0 :
                           ((~{74'b0}) >> u7v1l8233z7v63[6:0]);





wire ngn02441sf7gdrq30;
wire bf21b1jm9e5fpzs46pj4;
wire hahb3u6io9r35vs7a;
wire lyrxeddtp5exwibm;

wire zydb7odqtd2t5xehdt;
wire [162-1:0] hny7s8lqkaew1ht81;
wire [4-1:0] qz4o6968_5dqb5db3xgupbpl1;
wire ymtwckq9w36z4c;
wire [75-1:0] rdbo7d2_t715dy54ohz;
wire [4-1:0] stuv4gmzj7bpa1rm9df6woag;
wire k4rju_fn1hu;
wire gkh_mqfc5dvc;
wire a2iop2r7welh;
wire rdxa7brdak7c19s6;
wire md5qcqkyg3_k;

wire[12:0] h345ebh0vq = {2'b0,u49yq8sp[30:20]};
wire[12:0] vz7ad1k8gl = {2'b0,ahdfbec41y[30:20]};
wire[12:0] wr6ratxuyv = {2'b0,fwknegmn[30:20]};

wire[12:0] ps6tow7xumqnq69 = {5'b0,g91ks[30:23]};
wire[12:0] tb5ltp88utaxi_e = {5'b0,b04cwa[30:23]};
wire[12:0] mxhom0chw3b5o2 = {5'b0,pu0_qq[30:23]};

wire[52:0] rfcuzdq6uq3_k8v = {53{~(wijmhrmp5iul)}} & {53{ utngq}} & {~uc1umghn15g19b,fwknegmn[19:0],pu0_qq[31:0]};
wire[23:0] bm7h54zcw1xjwke = {24{~(wijmhrmp5iul)}} & {24{~utngq}} & {~uc1umghn15g19b, pu0_qq[22:0]};
wire[52:0] k6ydoqt3g9    = utngq ? rfcuzdq6uq3_k8v : {29'b0,bm7h54zcw1xjwke};

wire[12:0] cc9w1ghc8n = utngq ? h345ebh0vq : ps6tow7xumqnq69;
wire[12:0] wnw3w5n9j5i = utngq ? vz7ad1k8gl : tb5ltp88utaxi_e;
wire[12:0] fksw2fa96zbi = utngq ? wr6ratxuyv : mxhom0chw3b5o2;

wire [12:0] y1ck5xg3r1    = utngq ? 13'd1023: 13'd127;
wire [12:0] lsd7m09orucos = (cc9w1ghc8n + wnw3w5n9j5i + (~fksw2fa96zbi)) + (~(utngq ? 13'd966:13'd99)) + 1'b1;

wire [12:0] skjbk0pfgso_ = (cc9w1ghc8n + wnw3w5n9j5i + (~fksw2fa96zbi)) + (~(utngq ? 13'd965 : 13'd98) ) + 1'b1;
wire [12:0] mx2ztfgr0lzn = (cc9w1ghc8n + wnw3w5n9j5i + (~fksw2fa96zbi)) + (~(utngq ? 13'd967 : 13'd100)) + 1'b1;

wire ust6kl  = (mnwum_pdiuo ^ eu4746dfcv63) & (~uc1umghn15g19b);
wire sjgen2  = (~mnwum_pdiuo) & (~eu4746dfcv63) & (uc1umghn15g19b);
wire yxh7zvljyqqn = (~ust6kl) & (~sjgen2);

wire [12:0] d7zty5n83hwb7y;
wire [12:0] j9j9j7etnch5;
wire [12:0] yoysx5qs9zqcbwhf;

wire [12:0] x8n63zzgtm1 = ({13{k4rju_fn1hu }} & j9j9j7etnch5   ) 
                    | ({13{gkh_mqfc5dvc }} & yoysx5qs9zqcbwhf   )
	                | ({13{a2iop2r7welh}} & d7zty5n83hwb7y);

wire[52:0] l9zb_468vzbazfa6;
wire[23:0] aue5d6zocyk5kd3 = l9zb_468vzbazfa6[23:0];
wire[52:0] kw39fc_krl53t_d = l9zb_468vzbazfa6;

wire t6l_v4h7nke_u10 = x8n63zzgtm1[12];
wire [11:0] w6t4pgobkx_uhl = (m7s5rkmh ? 12'd163 : 12'd76);
wire cqhijr5kjq47ju8 = (~t6l_v4h7nke_u10) & (x8n63zzgtm1[11:0] > w6t4pgobkx_uhl);
wire eyrxcj62t1hhlhl5a    = (~t6l_v4h7nke_u10) & (~cqhijr5kjq47ju8);


wire [162+3+53-1:0] nr_k8g5yndryls = m7s5rkmh ? {1'b0,kw39fc_krl53t_d,108'b0,3'b0,53'b0} : 
                                              {1'b0,29'b0, aue5d6zocyk5kd3,108'b0,3'b0,53'b0};
wire [162+3+53-1:0] qxyuhl3_cfugo7n1xzi = m7s5rkmh ? {1'b0,53'b0,108'b0,3'b0,kw39fc_krl53t_d} :
                                                  {1'b0,53'b0,50'b0,3'b0,aue5d6zocyk5kd3,87'b0};
wire xvkeh6i41ok88w6 = (t6l_v4h7nke_u10 | cqhijr5kjq47ju8);

wire [162+3+53-1:0] mz1jva589d9eep1m5t = ({218{t6l_v4h7nke_u10}} & nr_k8g5yndryls) |
                                         ({218{cqhijr5kjq47ju8}} & qxyuhl3_cfugo7n1xzi);

wire [162+3+53-1:0] miz2cix1hgudijz739rzg95i = (nr_k8g5yndryls >> x8n63zzgtm1[7:0]);

wire uaj78s2_c4g_oj;

wire qcwfkcu7uqutzlw;

wire txe2dhitn770j9;
wire why9n7prff549n4;

wire [162+3+53-1:0] e6g87hojha93000xrh57dv;
wire [162+3+53-1:0] kfxmkdona0ind3vws9sfkn;

wire [162+3+53-1:0] sjebwuneqvcc = 
                          ({218{qcwfkcu7uqutzlw}} & kfxmkdona0ind3vws9sfkn) |
                          ({218{uaj78s2_c4g_oj}} & e6g87hojha93000xrh57dv);
wire [162+3+53-1:0] wlo72ilxg7lggpt = 
                          uzw0q1vxxy2cg ? (~sjebwuneqvcc) :
                                          sjebwuneqvcc;
assign zydb7odqtd2t5xehdt = uzw0q1vxxy2cg & 
                      ((~(|e6g87hojha93000xrh57dv[53+3-1:0])) & (~txe2dhitn770j9) | why9n7prff549n4 | md5qcqkyg3_k);


wire xv27tgo8wlbjoon2r_pla6qw8 = (&wlo72ilxg7lggpt[53-1:0]);
wire[3-1:0] inx58ut6yn0m9u8ddxgp1dzs = 
               uzw0q1vxxy2cg ? (wlo72ilxg7lggpt[53+3-1:53]+xv27tgo8wlbjoon2r_pla6qw8) :
                               wlo72ilxg7lggpt[53+3-1:53];
wire ynqs9guegsjl6wrn0lxbfm6 = 
               uzw0q1vxxy2cg ? (~xv27tgo8wlbjoon2r_pla6qw8) : (|wlo72ilxg7lggpt[53-1:0]);

assign qz4o6968_5dqb5db3xgupbpl1 = {inx58ut6yn0m9u8ddxgp1dzs, ynqs9guegsjl6wrn0lxbfm6};
assign hny7s8lqkaew1ht81 = wlo72ilxg7lggpt[162+3+53-1:53+3];
assign ngn02441sf7gdrq30 = t6l_v4h7nke_u10;

wire [75+3+24-1:0] k10u9kcpcjcbxjyv6ioeyes2v = {1'b0,e6g87hojha93000xrh57dv[(53+3+106+2+24-1):(53+3+106-48-24-3)]};
wire [75+3+24-1:0] txmbq5kkkg_43kcbeg = {1'b0,sjebwuneqvcc[(53+3+106+2+24-1):(53+3+106-48-24-3)]};

wire [75+3+24-1:0] oikeb907ubhp1wcadwcx = 
                    uzw0q1vxxy2cg ? (~txmbq5kkkg_43kcbeg) : txmbq5kkkg_43kcbeg;

assign ymtwckq9w36z4c = uzw0q1vxxy2cg & 
            ((~(|k10u9kcpcjcbxjyv6ioeyes2v[24+3-1:0])) & (~txe2dhitn770j9) | why9n7prff549n4 | md5qcqkyg3_k);

wire zqf__y5ie9otzt0zxfoyvd5m = (&oikeb907ubhp1wcadwcx[24-1:0]);

wire[3-1:0] mgeggocpknygj4oi61t8md35ey =
            uzw0q1vxxy2cg ? (oikeb907ubhp1wcadwcx[24+3-1:24] + zqf__y5ie9otzt0zxfoyvd5m) :
                            oikeb907ubhp1wcadwcx[24+3-1:24];

wire ketsbdosd29xg5aexr6mbz1pg = uzw0q1vxxy2cg ? (~zqf__y5ie9otzt0zxfoyvd5m) :
                            (|oikeb907ubhp1wcadwcx[24-1:0]);

assign stuv4gmzj7bpa1rm9df6woag = {mgeggocpknygj4oi61t8md35ey, ketsbdosd29xg5aexr6mbz1pg};
assign rdbo7d2_t715dy54ohz = oikeb907ubhp1wcadwcx[75+3+24-1:3+24];
assign hahb3u6io9r35vs7a = t6l_v4h7nke_u10;

assign bf21b1jm9e5fpzs46pj4 = why9n7prff549n4;
assign lyrxeddtp5exwibm = why9n7prff549n4;



assign vb_j3t59zgyb7r05r = m7s5rkmh ? ngn02441sf7gdrq30 : hahb3u6io9r35vs7a;
assign fi2z120absus4g = gma5v70c ? bf21b1jm9e5fpzs46pj4 : lyrxeddtp5exwibm;

wire [4-1:0] e_rkipm90ja1ygckb24b;
wire [4-1:0] iug5igicvl8jmztpzbzfkdvsb;
wire [4-1:0] vouwjch3wz7_qviomah6acriq;
wire [4-1:0] shh3tjbryqx94tx3p0bhj65rap;

wire [4-1:0] lu_owv4hd65jbek_fpn9r=gma5v70c ? qz4o6968_5dqb5db3xgupbpl1 : 4'b0;


wire [52:0] vwqwpqljff = {1'b0,u49yq8sp[19:0],g91ks[31:0]};

wire [52:0] t_5y5n4r = utngq ? {1'b0,u49yq8sp[19:0],g91ks[31:0]} :
                          {1'b0,23'b0,5'b0,1'b0, g91ks[22:0]} ;

wire [52:0] wj1f27njk3 = utngq ? {1'b0,u49yq8sp[19:0],g91ks[31:0]} :
                           {1'b0,23'b0,5'b0,1'b0,23'b0} ;

wire [52:0] i1 = utngq ? {1'b0,ahdfbec41y[19:0],b04cwa[31:0]} :
                       {1'b0,ahdfbec41y[22:0],5'b0,1'b0,b04cwa[22:0]} ;

wire [52:00] e2ry8ni = {53{~mnwum_pdiuo}} & {1'b0,23'b0,5'b0,(~eu4746dfcv63),b04cwa[22:0]};
wire [52:00] xyh6dubifq3 = {53{~eu4746dfcv63}} & {1'b0,23'b0,5'b0,1'b0,g91ks[22:0]};

wire [52:00] vim5vejcn = {53{~mnwum_pdiuo}} & {(~eu4746dfcv63),ahdfbec41y[19:0],b04cwa[31:0]} ;
wire [52:00] a8f6wteiequ6 = {53{~eu4746dfcv63}} & {1'b0,u49yq8sp[19:0],g91ks[31:0]} ;

wire [105:00] ms94p2owy = {53'b0, t_5y5n4r & {53{i1[00]}}       } ;
wire [105:00] x3cf2koq = {52'b0, t_5y5n4r & {53{i1[01]}}, 01'b0} ;
wire [105:00] pvq3jnz0 = {51'b0, t_5y5n4r & {53{i1[02]}}, 02'b0} ;
wire [105:00] ppqw59 = {50'b0, t_5y5n4r & {53{i1[03]}}, 03'b0} ;

wire [105:00] ugotq = {49'b0, t_5y5n4r & {53{i1[04]}}, 04'b0} ;
wire [105:00] eb1qolio5 = {48'b0, t_5y5n4r & {53{i1[05]}}, 05'b0} ;
wire [105:00] sq6nuqord = {47'b0, t_5y5n4r & {53{i1[06]}}, 06'b0} ;
wire [105:00] b9ol = {46'b0, t_5y5n4r & {53{i1[07]}}, 07'b0} ;

wire [105:00] piduv_l8m = {45'b0, t_5y5n4r & {53{i1[08]}}, 08'b0} ;
wire [105:00] nrousi = {44'b0, t_5y5n4r & {53{i1[09]}}, 09'b0} ;
wire [105:00] de2yw = {43'b0, t_5y5n4r & {53{i1[10]}}, 10'b0} ;
wire [105:00] lqr6n54ds = {42'b0, t_5y5n4r & {53{i1[11]}}, 11'b0} ;

wire [105:00] flkp4gvn4 = {41'b0, t_5y5n4r & {53{i1[12]}}, 12'b0} ;
wire [105:00] aa4a26a = {40'b0, t_5y5n4r & {53{i1[13]}}, 13'b0} ;
wire [105:00] w_2qgra2 = {39'b0, t_5y5n4r & {53{i1[14]}}, 14'b0} ;
wire [105:00] sdxfgz = {38'b0, t_5y5n4r & {53{i1[15]}}, 15'b0} ;

wire [105:00] ski6a = {37'b0, t_5y5n4r & {53{i1[16]}}, 16'b0} ;
wire [105:00] n0rxyxxr = {36'b0, t_5y5n4r & {53{i1[17]}}, 17'b0} ;
wire [105:00] ho9l9u21 = {35'b0, t_5y5n4r & {53{i1[18]}}, 18'b0} ;
wire [105:00] zuqqb4 = {34'b0, t_5y5n4r & {53{i1[19]}}, 19'b0} ;

wire [105:00] snpg9b = {33'b0, t_5y5n4r & {53{i1[20]}}, 20'b0} ;
wire [105:00] y_6xawz = {32'b0, t_5y5n4r & {53{i1[21]}}, 21'b0} ;
wire [105:00] gsm_x9kx = {31'b0, t_5y5n4r & {53{i1[22]}}, 22'b0} ;
wire [105:00] i2eoxni0c = {27'b0, t_5y5n4r & {53{i1[26]}}, 26'b0} ;

wire [105:00] vksr23hyn = utngq ? {30'b0, vwqwpqljff & {53{i1[23]}}, 23'b0} :{30'b0, e2ry8ni, 23'b0};
wire [105:00] o7myx = utngq ? {29'b0, vwqwpqljff & {53{i1[24]}}, 24'b0} :{30'b0, xyh6dubifq3, 23'b0};
wire [105:00] odvgzr = {28'b0, t_5y5n4r & {53{i1[25]}}, 25'b0} ;

wire [105:00] u4s5xf2f = {26'b0, t_5y5n4r & {53{i1[27]}}, 27'b0} ;
wire [105:00] tr8s9f = {25'b0, t_5y5n4r & {53{i1[28]}}, 28'b0} ;
wire [105:00] rb1s7rjun = {24'b0, wj1f27njk3 & {53{i1[29]}}, 29'b0} ;
wire [105:00] t9xi9g = {23'b0, wj1f27njk3 & {53{i1[30]}}, 30'b0} ;

wire [105:00] z4ivp = {22'b0, wj1f27njk3 & {53{i1[31]}}, 31'b0} ;
wire [105:00] mhyyf = {21'b0, wj1f27njk3 & {53{i1[32]}}, 32'b0} ;
wire [105:00] vovj = {20'b0, wj1f27njk3 & {53{i1[33]}}, 33'b0} ;
wire [105:00] rzjy = {19'b0, wj1f27njk3 & {53{i1[34]}}, 34'b0} ;

wire [105:00] nzxc = {18'b0, wj1f27njk3 & {53{i1[35]}}, 35'b0} ;
wire [105:00] jbo1 = {17'b0, wj1f27njk3 & {53{i1[36]}}, 36'b0} ;
wire [105:00] kt1r = {16'b0, wj1f27njk3 & {53{i1[37]}}, 37'b0} ;
wire [105:00] odf33uwsh = {15'b0, wj1f27njk3 & {53{i1[38]}}, 38'b0} ;

wire [105:00] zwhdwdts = {14'b0, wj1f27njk3 & {53{i1[39]}}, 39'b0} ;
wire [105:00] trlg2irc = {13'b0, wj1f27njk3 & {53{i1[40]}}, 40'b0} ;
wire [105:00] saaizm = {12'b0, wj1f27njk3 & {53{i1[41]}}, 41'b0} ;
wire [105:00] ti1yrg0n = {11'b0, wj1f27njk3 & {53{i1[42]}}, 42'b0} ;

wire [105:00] r1ynup = {10'b0, wj1f27njk3 & {53{i1[43]}}, 43'b0} ;
wire [105:00] uj7bx = {09'b0, wj1f27njk3 & {53{i1[44]}}, 44'b0} ;
wire [105:00] r2lj = {08'b0, wj1f27njk3 & {53{i1[45]}}, 45'b0} ;
wire [105:00] xn29hxzbi = {07'b0, wj1f27njk3 & {53{i1[46]}}, 46'b0} ;

wire [105:00] rbftzd = {06'b0, wj1f27njk3 & {53{i1[47]}}, 47'b0} ;
wire [105:00] lata8p_ = {05'b0, wj1f27njk3 & {53{i1[48]}}, 48'b0} ;
wire [105:00] om5py = {04'b0, wj1f27njk3 & {53{i1[49]}}, 49'b0} ;
wire [105:00] q7uoa = {03'b0, wj1f27njk3 & {53{i1[50]}}, 50'b0} ;

wire [105:00] tlo5ayfb3 = {02'b0, wj1f27njk3 & {53{i1[51]}}, 51'b0} ;
wire [105:00] lrlu4qd = utngq ? {01'b0, vim5vejcn, 52'b0} :{01'b0, 53'b0, 52'b0};
wire [105:00] tp0q8a9 = utngq ? {01'b0, a8f6wteiequ6, 52'b0} :{01'b0, 53'b0, 52'b0};

assign pk0153efgrg0 = nc2dhbcdb26q;
assign cpq3wxamh6ly = rcs83fuv1yxfs;

ikddk6f6fc0_2t0g5wt #(106) h_z_kq_953d61a(.frgfco(ms94p2owy), .ii(x3cf2koq), .fij51v(pvq3jnz0), .cuzhl9(ppqw59), .c(b_0ht), .s(oazfr2ucb));
ikddk6f6fc0_2t0g5wt #(106) bwm1_sh8ecm96koc6(.frgfco(ugotq), .ii(eb1qolio5), .fij51v(sq6nuqord), .cuzhl9(b9ol), .c(p07jru), .s(is4rk));
ikddk6f6fc0_2t0g5wt #(106) sf6r8y8jn2fp2m(.frgfco(piduv_l8m), .ii(nrousi), .fij51v(de2yw), .cuzhl9(lqr6n54ds), .c(h5w1j3), .s(vs1z8));
ikddk6f6fc0_2t0g5wt #(106) y0l52hfl3d_m92jn(.frgfco(flkp4gvn4), .ii(aa4a26a), .fij51v(w_2qgra2), .cuzhl9(sdxfgz), .c(hk7neg5b6), .s(x_5tn8w));
ikddk6f6fc0_2t0g5wt #(106) zeatop9zhu_ktn(.frgfco(ski6a), .ii(n0rxyxxr), .fij51v(ho9l9u21), .cuzhl9(zuqqb4), .c(xdzb4s0ejm), .s(tr2ajiq));
ikddk6f6fc0_2t0g5wt #(106) tjk53xfhdy2csr1k(.frgfco(snpg9b), .ii(y_6xawz), .fij51v(gsm_x9kx), .cuzhl9(i2eoxni0c), .c(f0k2ir301f), .s(n2fm6));
ikddk6f6fc0_2t0g5wt #(106) phvgwjbqn6nbmx(.frgfco(u4s5xf2f), .ii(tr8s9f), .fij51v(rb1s7rjun), .cuzhl9(t9xi9g), .c(kf_ejf), .s(olreui));
ikddk6f6fc0_2t0g5wt #(106) klo99kt0yecyq(.frgfco(z4ivp), .ii(mhyyf), .fij51v(vovj), .cuzhl9(rzjy), .c(nh9i6q51r), .s(zu59l2mmd));
ikddk6f6fc0_2t0g5wt #(106) u8nbojg6_i8m1(.frgfco(nzxc), .ii(jbo1), .fij51v(kt1r), .cuzhl9(odf33uwsh), .c(dtoeq), .s(m5s6xnj));
ikddk6f6fc0_2t0g5wt #(106) cqu3wqyv2zg07c(.frgfco(zwhdwdts), .ii(trlg2irc), .fij51v(saaizm), .cuzhl9(ti1yrg0n), .c(rzu745tt29), .s(ca8pgl9));
ikddk6f6fc0_2t0g5wt #(106) a_lyni_fs_rf573(.frgfco(r1ynup), .ii(uj7bx), .fij51v(r2lj), .cuzhl9(xn29hxzbi), .c(wqjzd4lir), .s(aeeu2arrcv));
ikddk6f6fc0_2t0g5wt #(106) o_yfzp5lbbgkn5g(.frgfco(rbftzd), .ii(lata8p_), .fij51v(om5py), .cuzhl9(q7uoa), .c(aihp3cuom0), .s(uucty));

j3aa8h4yagvjsr416mg #(106) agwu0uf8jew62x1(.frgfco(vksr23hyn), .ii(o7myx), .fij51v(odvgzr), .c(cpkrdt), .s(td137));
j3aa8h4yagvjsr416mg #(106) nwqo8cl2_md6kj(.frgfco(tlo5ayfb3), .ii(lrlu4qd), .fij51v(tp0q8a9), .c(rwnza0fed), .s(lfm5om4i85));


ikddk6f6fc0_2t0g5wt #(106) u6sgcgjiq33_uf(.frgfco(zf2wuu6f), .ii(ipmcb4953), .fij51v(vje27h4vio), .cuzhl9(skablhb13q), .c(fz5l6am6), .s(fxx71cde0f));
ikddk6f6fc0_2t0g5wt #(106) ozf9flh2yrvt(.frgfco(cb_65dtz), .ii(mue2czm03), .fij51v(apzd3bocb0jlz), .cuzhl9(qsofrkqvi), .c(gizb4v58_bc), .s(ydnoov3_7x));
ikddk6f6fc0_2t0g5wt #(106) m9qv8ygeiptdo(.frgfco(tbqp2_p5b), .ii(vask7qpb), .fij51v(vkbk0udu), .cuzhl9(y9vjbgehnlld), .c(e9z05qhld0), .s(uf8wgiec));
ikddk6f6fc0_2t0g5wt #(106) c_0cyk1r8q0hqat(.frgfco(snujns_17o), .ii(r49be1odf), .fij51v(fmmslemj9z9), .cuzhl9(tezkbiwpx10os), .c(sq4cj16ceo), .s(dqlgpi77o));
ikddk6f6fc0_2t0g5wt #(106) c0qeqi8sp_yk(.frgfco(ezb1_13jolmi), .ii(vgfckvnmljw), .fij51v(ps3bgs1w), .cuzhl9(wbbij0elfpd), .c(pw7_78ztt), .s(k4g2t42mbrb));
ikddk6f6fc0_2t0g5wt #(106) jmnnwewzh7mr9(.frgfco(vm7box2gikw3), .ii(wxqo_7ac7g), .fij51v(ufo0585p), .cuzhl9(gyh98b_6jowgw), .c(edqpyho0og), .s(go2kpgsuttj));
ikddk6f6fc0_2t0g5wt #(106) cl9r_064dvyo9(.frgfco(nqh156gtt8f), .ii(xjc8hz47unk4), .fij51v(crlqmi91i), .cuzhl9(xuugnk6md694i), .c(nc2dhbcdb26q), .s(rcs83fuv1yxfs));

ikddk6f6fc0_2t0g5wt #(106) hdz6o7o41zs7c(.frgfco(fz5l6am6), .ii(fxx71cde0f), .fij51v(gizb4v58_bc), .cuzhl9(ydnoov3_7x), .c(at16xua1qxc), .s(ai4n2ob_j7ocd));
ikddk6f6fc0_2t0g5wt #(106) iuekexy9l8owwrsvr(.frgfco(e9z05qhld0), .ii(uf8wgiec), .fij51v(sq4cj16ceo), .cuzhl9(dqlgpi77o), .c(o0s11rb3), .s(nzl699hjo));
ikddk6f6fc0_2t0g5wt #(106) mfzx4qx276e3(.frgfco(pw7_78ztt), .ii(k4g2t42mbrb), .fij51v(edqpyho0og), .cuzhl9(go2kpgsuttj), .c(jqprtktb8qr8), .s(frs3fk930avn));

ikddk6f6fc0_2t0g5wt #(106) daedh1f38p5y(.frgfco(at16xua1qxc), .ii(ai4n2ob_j7ocd), .fij51v(o0s11rb3), .cuzhl9(nzl699hjo), .c(kaxkamth), .s(vou_g00czb2));
ikddk6f6fc0_2t0g5wt #(106) r6p84hobtibxo2s7(.frgfco(jqprtktb8qr8), .ii(frs3fk930avn), .fij51v(pk0153efgrg0), .cuzhl9(cpq3wxamh6ly), .c(rbm2min6), .s(qtui513wjhfz));

ikddk6f6fc0_2t0g5wt #(106) xg5_6kqnhhavvt(.frgfco(mknydvsmn87), .ii(ga_yvggsogewp), .fij51v(z49e6oo_eurd), .cuzhl9(ttw8izs6), .c(z7z1y_k7), .s(sxo8i0fku66y));

wire [49-1:0] aeq24nddlbz7ivtqpajs;
wire [49-1:0] t30tnjjxkq990ukxik  ;
wire [9-1:0]  dhporcw1lcehxqjz0gujrc6c;
wire [49-1:0] ds6eargsa5f6nd7lwc37bed3js;
wire [49-1:0] do3dp95tfex0l3octe3jt  ;
wire [9-1:0]  tyaslfzhg2fu2p6m6x6;
wire [107-1:0] h2a5ydn7s_8l_gns9rz4hy9;
wire [107-1:0] cf738tb7h4toemtbbo0;

wire[106-1:0] dzjz6ib3 = z7z1y_k7;
wire[106-1:0] hlk5nd7kmyw77 = sxo8i0fku66y;


wire [107-1:0] dm1r_d8yslyd5itzw15 = {1'b0,dzjz6ib3};
wire [107-1:0] kupue75e6nzmbuw1wb3 = {1'b0,hlk5nd7kmyw77};
wire [107-1:0] anmdrteg214tvjess = {1'b0,hny7s8lqkaew1ht81[106-1:0]};

wire [49-1:0] z87rew964zzvrlg6iw = {1'b0,dzjz6ib3[47:0]};
wire [49-1:0] ca0ia87tlz4rigmk1 = {1'b0,hlk5nd7kmyw77[47:0]};
wire [49-1:0] sdw5ph6ql8ph8uefuk = {1'b0,rdbo7d2_t715dy54ohz[48-1:0]};


wire [107-1:0] d6627emd0xqqrn049 = gma5v70c ? dm1r_d8yslyd5itzw15 :{49'b0, 9'b0, z87rew964zzvrlg6iw};
wire [107-1:0] hf3p6bpo8sps667y2kdtd = gma5v70c ? kupue75e6nzmbuw1wb3 :{49'b0, 9'b0, ca0ia87tlz4rigmk1};
wire [107-1:0] h5xr9til85y0zw4d8w = gma5v70c ? anmdrteg214tvjess :{49'b0, 9'b0, sdw5ph6ql8ph8uefuk};



j3aa8h4yagvjsr416mg #(107) z22or8aiq2en4fhnqm1(
    .frgfco(d6627emd0xqqrn049), 
    .ii(hf3p6bpo8sps667y2kdtd), 
    .fij51v(h5xr9til85y0zw4d8w),
    .c(h2a5ydn7s_8l_gns9rz4hy9), 
    .s(cf738tb7h4toemtbbo0)
);
wire [107-1:0] xfeqb_2mh_vxx6vtn5cg0i = h2a5ydn7s_8l_gns9rz4hy9;
wire [107-1:0] f94g6z8m66ha1otod98   = cf738tb7h4toemtbbo0  ;


assign {ds6eargsa5f6nd7lwc37bed3js, dhporcw1lcehxqjz0gujrc6c, aeq24nddlbz7ivtqpajs} = h2a5ydn7s_8l_gns9rz4hy9;
assign {do3dp95tfex0l3octe3jt,   tyaslfzhg2fu2p6m6x6,   t30tnjjxkq990ukxik}   = cf738tb7h4toemtbbo0;

wire itl_t4bnss1vfv = uzw0q1vxxy2cg;
wire zvpmtk3x6t7gadtlw9x = uzw0q1vxxy2cg;


wire [163-1:0] ms697g8rg351b9m = {hny7s8lqkaew1ht81[162-1:106],f94g6z8m66ha1otod98[106-1:0],zydb7odqtd2t5xehdt};
wire [163-1:0] xvl5c9bnddhc9g = {55'b0,xfeqb_2mh_vxx6vtn5cg0i[107-1:0],itl_t4bnss1vfv};

wire [76-1:0] kgtwswp5fbffo = {76{~kbjfvasuqsn4g}} & 
    {rdbo7d2_t715dy54ohz[75-1:48],t30tnjjxkq990ukxik[48-1:0],ymtwckq9w36z4c};
wire [76-1:0] xqd_yyuw_5nzslx6wf = {76{~kbjfvasuqsn4g}} &
    {26'b0,aeq24nddlbz7ivtqpajs[49-1:0],zvpmtk3x6t7gadtlw9x};

wire [164-1:0] cdut53tpwkh302 = gma5v70c ? {ms697g8rg351b9m[163-1],ms697g8rg351b9m} 
                              : {77'b0,10'b0, kgtwswp5fbffo[76-1],kgtwswp5fbffo};
wire [164-1:0] bpzk76nrkskhqgqeym = gma5v70c ? {xvl5c9bnddhc9g[163-1],xvl5c9bnddhc9g} 
                              : {77'b0,10'b0, xqd_yyuw_5nzslx6wf[76-1],xqd_yyuw_5nzslx6wf};

wire vfoky1zddkg25vwisss4;
wire [163-1:0] b5wkg2i72jl6_5a;

wire [164-1:0] u_1lz3gy_x6_ha5hckf;
wire [164-1:0] mzs3mhha1mu673a02e;

assign {b5wkg2i72jl6_5a,vfoky1zddkg25vwisss4} = (u_1lz3gy_x6_ha5hckf + mzs3mhha1mu673a02e);


wire xah621mzhwehgh8q2k05;
wire dbbae0augcbydoflecfu8282_;
wire [76-1:0] pl8amgmncf10p418ylg;
wire [76-1:0] nxflth7__8qg2yxpps;
wire [10-1:0] qqob49t7jt82sljhfv8;

assign {nxflth7__8qg2yxpps, 
        dbbae0augcbydoflecfu8282_,
        qqob49t7jt82sljhfv8,
        pl8amgmncf10p418ylg,
        xah621mzhwehgh8q2k05}
        = {b5wkg2i72jl6_5a,vfoky1zddkg25vwisss4};

wire w5apvcv2k2460m846kcm2wn = vfoky1zddkg25vwisss4;
wire [163-1:0] uiy_h8mivw_xmbn8e =  b5wkg2i72jl6_5a;
wire ihnqe0vmp0coywgoq4xj1m = mb8pmo37pwn ? w5apvcv2k2460m846kcm2wn : xah621mzhwehgh8q2k05;
wire [163-1:0] jrdafd333s5adeh15 = mb8pmo37pwn ? uiy_h8mivw_xmbn8e : {pl8amgmncf10p418ylg,vouwjch3wz7_qviomah6acriq,83'b0};


wire[8-1:0] w770780rlqi6;

wire[255:0] o_q0p_iqbc1vaaavo9u2z4 = gma5v70c ? {ms697g8rg351b9m[163-1],ms697g8rg351b9m,2'b01,{(256-164-2){1'b0}}}
                                : {kgtwswp5fbffo[76-1],kgtwswp5fbffo,2'b01,{(256-77-2){1'b0}}};
wire[255:0] iugf352komlvpzztjw1 = gma5v70c ? {xvl5c9bnddhc9g[163-1],xvl5c9bnddhc9g,2'b00,{(256-164-2){1'b0}}}
                                : {xqd_yyuw_5nzslx6wf[76-1],xqd_yyuw_5nzslx6wf,2'b00,{(256-77-2){1'b0}}};

wire[255:0] k8uhevn2sa7r2v83o3l = gma5v70c ? {2'b0,wfjl06kozsl7u3d95drhv8,{(256-163){1'b1}}}
                                : {2'b0,gbyt7t2vj0c3ymg7p6dqxz,{(256-76){1'b1}}};

wire[256-1:0] djohwtsa;
wire [256-1:0] hzc1y = (djohwtsa | k8uhevn2sa7r2v83o3l);
wire [256-1:0] gzevpqks4ek;

genvar i;

generate
  for (i=0;i<256;i=i+1) begin: k521v71_bypqy
    if(i==0) begin:l9j7mf
      ggzvoy2zvu8ryca4ylw0 opkdldl0emb7 (
           .jq6ebmv({o_q0p_iqbc1vaaavo9u2z4[i+1:i],1'b0}),
           .f7rj({iugf352komlvpzztjw1[i+1:i],1'b0}),
           .uriczc(djohwtsa[i])
       );
    end
    else if(i==(256-1)) begin:w8m0qhqxdv9nq
      ggzvoy2zvu8ryca4ylw0 opkdldl0emb7 (
          .jq6ebmv({o_q0p_iqbc1vaaavo9u2z4[i],o_q0p_iqbc1vaaavo9u2z4[i:i-1]}), 
          .f7rj({iugf352komlvpzztjw1[i],iugf352komlvpzztjw1[i:i-1]}),
          .uriczc(djohwtsa[i])
      );
    end
    else begin:r9bggk8u55
      ggzvoy2zvu8ryca4ylw0 opkdldl0emb7 (
          .jq6ebmv(o_q0p_iqbc1vaaavo9u2z4[i+1:i-1]),
          .f7rj(iugf352komlvpzztjw1[i+1:i-1]),
          .uriczc(djohwtsa[i])
      );
    end
  end
endgenerate



uwtp9d4cv1y3gqfa7u3jo #(.onr7l(256), .hw3qvr(8)) w5ocjz3zbd5(.bjh(gzevpqks4ek), .ht70(w770780rlqi6));


wire[8-1:0] hlmjo66nn_vl0tc;



wire dhjwqosv4ycmcnx50oozvu;
wire q58jwqackb28ri3ianjbm5;
wire oystrf6qb5s0k8;

wire ghwsivxem72r_3m__sye = jrdafd333s5adeh15[163-1];

wire [163-1:0] m_n4zvnbl0boxtgug8;
wire wxy_rmva3xpos0 = (~sk_hgye1w_624w_ & nunpqy34d5rby3u2c & m_n4zvnbl0boxtgug8[163-1])
                | (sk_hgye1w_624w_ & (~nunpqy34d5rby3u2c) & (~m_n4zvnbl0boxtgug8[163-1]))
                | (~sk_hgye1w_624w_ & (~nunpqy34d5rby3u2c) & m_n4zvnbl0boxtgug8[163-1])
                | (sk_hgye1w_624w_ & nunpqy34d5rby3u2c & (~m_n4zvnbl0boxtgug8[163-1]));

wire [162-1:0] clkxpqou7ir6og;
wire [12:0] ivv694h2frwdqy0wg;
wire [12:0] rlmpudbadjn3njp6t3pg;
wire [12:0] ugxsstwfs7ud2ujj76;
wire [5:0] j_59k0vdcyzjg4dx9zjnwu1t;
wire w9teop0xh2jhgpg7iq_e;


wire [162-1:0] s2ojaltbql2 = m_n4zvnbl0boxtgug8[162-1:0];

wire sdalsx = b7x36_v4z0jlprnsb8vmn2;

wire [162-1:0] l951bdmlxqvlspmq7r  = {162{dhjwqosv4ycmcnx50oozvu}} ^ s2ojaltbql2;
wire [4-1:0] n0donsvsxqqra_u_1jj61 = {4{dhjwqosv4ycmcnx50oozvu}} ^ iug5igicvl8jmztpzbzfkdvsb;

wire l67y6vh9y51_i70 = (|xrc71n3kb03z2[12:6]);

wire [64-1:0] o_n5znqhy2;
wire [64-1:0] l3tc4muxpuaq0qp;
assign {o_n5znqhy2, l3tc4muxpuaq0qp} = l67y6vh9y51_i70 ? 128'b0 : 
    ({l951bdmlxqvlspmq7r[(162-1):(162-64)], {64{dhjwqosv4ycmcnx50oozvu}}} >> xrc71n3kb03z2[5:0]);

wire cdaynisyl0uvoktybe746  = (|s2ojaltbql2[162-64-1:0]);
wire vx_r1bmaww2bn4_312222 = (|s2ojaltbql2[161:98]) | cdaynisyl0uvoktybe746;

wire senhojkui8cidnqn2x3 = sdalsx &
                      (
                      l67y6vh9y51_i70 ? (vx_r1bmaww2bn4_312222 | (|iug5igicvl8jmztpzbzfkdvsb))
                                      : (|{cdaynisyl0uvoktybe746,iug5igicvl8jmztpzbzfkdvsb})
                      );

wire gn57dcv7d1vnwydmbqxgj8c1r8qc  = (&l951bdmlxqvlspmq7r[162-64-1:0]);
wire wqjtbrwyic68dlri5wvlgo3gufd1y = (&l951bdmlxqvlspmq7r[161:98]) & gn57dcv7d1vnwydmbqxgj8c1r8qc;

wire momttpny95s75_yad3b=sdalsx &
                      (
                      l67y6vh9y51_i70 ? (wqjtbrwyic68dlri5wvlgo3gufd1y & (&n0donsvsxqqra_u_1jj61))
                                       : (&{gn57dcv7d1vnwydmbqxgj8c1r8qc,n0donsvsxqqra_u_1jj61})
                      );

wire [162-1:0] q69e44l8s = {o_n5znqhy2,
                         l3tc4muxpuaq0qp,
                         (dhjwqosv4ycmcnx50oozvu ? momttpny95s75_yad3b : senhojkui8cidnqn2x3),
                         {33{dhjwqosv4ycmcnx50oozvu}}};

wire tusk45 = ~sdalsx;

wire [162-1:0] jvpxh7o;
wire [5:0] kwmsnzpbngxnqic88k;


u6rhkw924ptxmc8p5wde #(.onr7l(162+6)) wm3aijsc1tbqt0(
    .bjh     ({2'b0,s2ojaltbql2,iug5igicvl8jmztpzbzfkdvsb}),
    .a856yvdz (dhjwqosv4ycmcnx50oozvu),
    .w40py     (hlmjo66nn_vl0tc[7:0]),
    .adqhji    ({jvpxh7o, kwmsnzpbngxnqic88k}) 
);

wire md5368bgnloobe7ue9s5t7 = ({5'b0,hlmjo66nn_vl0tc} == (crtsq13_r9b5_i8j + 2'd2));

wire sq8tpegqmuekghx= (~md5368bgnloobe7ue9s5t7) & tusk45 & (~jvpxh7o[161]) & (~jvpxh7o[160]);

wire [12:0] a4zgmbptgvt41 = duxpze1m6dlz2rx + (~{5'b0,hlmjo66nn_vl0tc}) + 2'd3;

wire [12:0] laqt92c1184ni2n = duxpze1m6dlz2rx + (~{5'b0,hlmjo66nn_vl0tc}) + 2'd2;

wire [12:0] z48eqfoi7usg91y = duxpze1m6dlz2rx + (~{5'b0,hlmjo66nn_vl0tc}) + 3'd4;

wire [6-1:0] xsd5n8eqwh_b0n2vvvcup = ({6{tusk45}} & kwmsnzpbngxnqic88k)
			                   | ({6{sdalsx}} & 6'b0);

wire [162-1:0] pf46x9eq8b = ({162{tusk45}} & jvpxh7o)
			              | ({162{sdalsx}} & q69e44l8s);

wire [12:0] n0_3jdbndqe18 = ({13{tusk45}} & (a4zgmbptgvt41))
			         | ({13{sdalsx}} & 13'b1);

wire [12:0] gk6mz5clwkmam2g5 = ({13{tusk45}} & (laqt92c1184ni2n))
			            | ({13{sdalsx}} & 13'h0);

wire [12:0] e32ykab5wzwl8tnz = ({13{tusk45}} & (z48eqfoi7usg91y))
			            | ({13{sdalsx}} & 13'h2);

wire [63:0] ejo3ojh7m47_vp7sji6u_1;
wire [31:0] ei1aqk1e3hxolgk4w5xi_;
wire [7-1:0] ttnbtbp7drj;
wire [7-1:0] br_f61q6qczmz8;


wire ily0succ6y;
wire [162-1:0] gnbywwrr_k;
wire [162-1:0] zjk41qe_zcaealqo17u;
wire [162-1:0] rfia5mjpt09_4q8;
wire [162-1:0] n4vek2gzjekymw9k;
wire [162-1:0] n44e3s18fws7;
wire [6-1:0] obuwrw7em1vneml6md5g4tosu83;
wire rpt9_hjj40vp;

assign {n44e3s18fws7,obuwrw7em1vneml6md5g4tosu83} = 
    q58jwqackb28ri3ianjbm5 ? 
    (~{clkxpqou7ir6og,j_59k0vdcyzjg4dx9zjnwu1t} + 1'b1) :
    {clkxpqou7ir6og,j_59k0vdcyzjg4dx9zjnwu1t};

wire [162-1:0] ixu6irynjvjq6e =
    w9teop0xh2jhgpg7iq_e ? {n44e3s18fws7[162-2:0],obuwrw7em1vneml6md5g4tosu83[5]} : clkxpqou7ir6og;

wire [6-1:0] v9629b224rm418t6dl_2zdsn11 =
    w9teop0xh2jhgpg7iq_e ? {obuwrw7em1vneml6md5g4tosu83[4:0],q58jwqackb28ri3ianjbm5} :obuwrw7em1vneml6md5g4tosu83;

wire [24:0] so9eltti3mebugoo1myjy = ixu6irynjvjq6e[162-1:137];
wire [53:0] v4vz09_wnzl9u5octk7fx = ixu6irynjvjq6e[162-1:108]; 

wire [162-1:0] e9le = clkxpqou7ir6og;

wire [6-1:0] q0hij14o4y9qz6jhd = j_59k0vdcyzjg4dx9zjnwu1t;

wire k2jhucqujtuxh9bypblm = (|e9le[104:0]) | (|q0hij14o4y9qz6jhd);
wire iw957u8bwe3p0p11u = (&e9le[104:0]) & (&q0hij14o4y9qz6jhd);
wire jqafgdyih6p5y   = q58jwqackb28ri3ianjbm5 & iw957u8bwe3p0p11u;
assign n4vek2gzjekymw9k[108:105] = jqafgdyih6p5y ? (e9le[108:105] + 1'b1) : e9le[108:105];

wire mupaafv3dcalham02 = (&e9le[108:105]) & iw957u8bwe3p0p11u;
wire f022xf7q2yd19v4lbr1 = q58jwqackb28ri3ianjbm5 & mupaafv3dcalham02;
wire [4:0] ep5x4fv842l1sidj_keaw6v3t = 
    jqafgdyih6p5y ? ({1'b0,e9le[108:105]} + (w9teop0xh2jhgpg7iq_e ? {1'b0,1'b0,1'b1,1'b0,1'b1} : {1'b0,1'b1,1'b0,1'b0,1'b1}))
                    : ({1'b0,e9le[108:105]} + (w9teop0xh2jhgpg7iq_e ? {1'b0,1'b0,1'b1,1'b0,1'b0} : {1'b0,1'b1,1'b0,1'b0,1'b0}));

wire z9s1fu2p0vnmcm180v = ep5x4fv842l1sidj_keaw6v3t[4] & rpt9_hjj40vp;

wire l723_8vel4l18ye2 = (f022xf7q2yd19v4lbr1 | z9s1fu2p0vnmcm180v);

assign rfia5mjpt09_4q8[162-1:109]   = l723_8vel4l18ye2     ? (e9le[162-1:109] + 1'b1) : e9le[162-1:109];
assign n4vek2gzjekymw9k[162-1:109] = f022xf7q2yd19v4lbr1 ? (e9le[162-1:109] + 1'b1) : e9le[162-1:109];

wire hyagjmt16a_zstxtwf8jm = q58jwqackb28ri3ianjbm5 & (~iw957u8bwe3p0p11u) | (~q58jwqackb28ri3ianjbm5) & k2jhucqujtuxh9bypblm;
assign rfia5mjpt09_4q8[108:105] = rpt9_hjj40vp ? ep5x4fv842l1sidj_keaw6v3t[3:0] : n4vek2gzjekymw9k[108:105];
assign rfia5mjpt09_4q8[104:0]   = {hyagjmt16a_zstxtwf8jm,104'b0};
assign n4vek2gzjekymw9k[104:0] = {hyagjmt16a_zstxtwf8jm,104'b0};


wire u__9eqy_i2jtqaunig = (|e9le[133:0]) | (|q0hij14o4y9qz6jhd);
wire lghj4qt884nyzzs68fn = (&e9le[133:0]) & (&q0hij14o4y9qz6jhd);
wire ypiwt5rii6ld68i   = q58jwqackb28ri3ianjbm5 & lghj4qt884nyzzs68fn;
assign zjk41qe_zcaealqo17u[137:134] = ypiwt5rii6ld68i ? (e9le[137:134] + 1'b1) : e9le[137:134];

wire qzmmowot_ypheq7p = (&e9le[137:134]) & lghj4qt884nyzzs68fn;
wire za4u9g1m8rh3gbyu9b4k = q58jwqackb28ri3ianjbm5 & qzmmowot_ypheq7p;
wire [4:0] ejjy3t_onreouaxmzmtxqqnx = 
    ypiwt5rii6ld68i ? 
    {1'b0,e9le[137:134]} + (w9teop0xh2jhgpg7iq_e ? {1'b0,1'b0,1'b1,1'b0,1'b1} : {1'b0,1'b1,1'b0,1'b0,1'b1})
   :{1'b0,e9le[137:134]} + (w9teop0xh2jhgpg7iq_e ? {1'b0,1'b0,1'b1,1'b0,1'b0} : {1'b0,1'b1,1'b0,1'b0,1'b0});

wire x8tab32xn3zbroe5qqfqd = ejjy3t_onreouaxmzmtxqqnx[4] & ily0succ6y;

wire wtdg3rn2yqda2cp0 = za4u9g1m8rh3gbyu9b4k | x8tab32xn3zbroe5qqfqd;

wire i8jcp8i0jtrqr2nntrq4 = 
    (q58jwqackb28ri3ianjbm5 & (~lghj4qt884nyzzs68fn)) | 
    ((~q58jwqackb28ri3ianjbm5) & u__9eqy_i2jtqaunig);

assign gnbywwrr_k[133:0]       = {i8jcp8i0jtrqr2nntrq4,133'b0};
assign zjk41qe_zcaealqo17u[133:0] = gnbywwrr_k[133:0];

assign gnbywwrr_k[137:134] = ily0succ6y ? ejjy3t_onreouaxmzmtxqqnx[3:0] : zjk41qe_zcaealqo17u[137:134];

assign gnbywwrr_k[162-1:138] = wtdg3rn2yqda2cp0 ? (e9le[162-1:138] + 1'b1) : e9le[162-1:138];
assign zjk41qe_zcaealqo17u[162-1:138] = za4u9g1m8rh3gbyu9b4k ? (e9le[162-1:138] + 1'b1) : e9le[162-1:138];

wire v0yrssab8j= (w9teop0xh2jhgpg7iq_e ? n4vek2gzjekymw9k[107]      : n4vek2gzjekymw9k[108]     );
wire lh6unwr3hep  = (w9teop0xh2jhgpg7iq_e ? n4vek2gzjekymw9k[106]      : n4vek2gzjekymw9k[107]     );
wire rl79o_xu  = (w9teop0xh2jhgpg7iq_e ? n4vek2gzjekymw9k[105]      : n4vek2gzjekymw9k[106]     );
wire u2n0m_qrom5l  = (w9teop0xh2jhgpg7iq_e ? (|n4vek2gzjekymw9k[104:0]) : (|n4vek2gzjekymw9k[105:0]));

el7n_zz16sk_ntvue9v yh51n3oxckg3yvuobud ( 
                 .l     (v0yrssab8j), 
                 .g     (lh6unwr3hep),
                 .r     (rl79o_xu),
                 .s     (u2n0m_qrom5l), 
                 .ly53de  (oystrf6qb5s0k8),
                 .nfj6b    (ach5cwxikdp),
                 .f6dc_rhcaz(rpt9_hjj40vp) 
             );

wire w4z2jjbw0dlao = w9teop0xh2jhgpg7iq_e ? zjk41qe_zcaealqo17u[136]      : zjk41qe_zcaealqo17u[137]     ;
wire ew042ocnt   = w9teop0xh2jhgpg7iq_e ? zjk41qe_zcaealqo17u[135]      : zjk41qe_zcaealqo17u[136]     ;
wire oy6dz1dkg4cz   = w9teop0xh2jhgpg7iq_e ? zjk41qe_zcaealqo17u[134]      : zjk41qe_zcaealqo17u[135]     ;
wire v9x3wim2co7eb   = w9teop0xh2jhgpg7iq_e ? (|zjk41qe_zcaealqo17u[133:0]) : (|zjk41qe_zcaealqo17u[134:0]);

el7n_zz16sk_ntvue9v k7oond8b7ihic4auo ( 
                 .l     (w4z2jjbw0dlao), 
                 .g     (ew042ocnt),
                 .r     (oy6dz1dkg4cz),
                 .s     (v9x3wim2co7eb), 
                 .ly53de  (oystrf6qb5s0k8),
                 .nfj6b    (ach5cwxikdp),
                 .f6dc_rhcaz(ily0succ6y) );

wire [24:0] uo557q_42160ch = zjk41qe_zcaealqo17u[162-1:137];
wire [24:0] mmhfmsr3zdjrk2     = gnbywwrr_k[162-1:137];
wire yf80w6zpsarvnsrd5cnj3etc  = gnbywwrr_k[136];

wire [53:0] t_t7vy1dpix0yv7cp = n4vek2gzjekymw9k[162-1:108]; 
wire [53:0] fvonvyekztwxw4     = rfia5mjpt09_4q8[162-1:108];
wire ckpku1ypqvuy811tcixg  = rfia5mjpt09_4q8[107];

wire gi2lnto4gl0sc9      = (~(|{e9le,q0hij14o4y9qz6jhd})) & (~q58jwqackb28ri3ianjbm5);
wire co3mgjjdm6kydzn01y2wdjd = (ach5cwxikdp == 3'b10);

wire if0armmro_9a3439fyk6erutd6o   = l723_8vel4l18ye2 & (e9le[162-1-2:109] == (~(51'b0)));
wire rdrrbb27q9ldjkeiukgt5kthnq   = wtdg3rn2yqda2cp0 & (e9le[162-1-2:138] == (~(22'b0)));

wire kf48fwg3pjcnaeqo70skmm4ok = l723_8vel4l18ye2 & (e9le[162-1-1:109] == (~(52'b0)));
wire g5xi2zag08ihplpf5qzve6rd3ar4w = wtdg3rn2yqda2cp0 & (e9le[162-1-1:138] == (~(23'b0)));

wire atm4upf52hg3l87yr     = w9teop0xh2jhgpg7iq_e & (~if0armmro_9a3439fyk6erutd6o);
wire j384788dhg6btg4     = w9teop0xh2jhgpg7iq_e & (~rdrrbb27q9ldjkeiukgt5kthnq);

wire hq1a13ibszmpmt0aun = (~w9teop0xh2jhgpg7iq_e) & kf48fwg3pjcnaeqo70skmm4ok;
wire mt90aszfju_i2zee = (~w9teop0xh2jhgpg7iq_e) & g5xi2zag08ihplpf5qzve6rd3ar4w;

wire wy5xxr8o4e6 = (~hq1a13ibszmpmt0aun) & (~atm4upf52hg3l87yr);
wire ox0usqzivjky70 = (~mt90aszfju_i2zee) & (~j384788dhg6btg4);

wire v0k68izxc00gi8fsnfdw3rars6 = hq1a13ibszmpmt0aun | (atm4upf52hg3l87yr ? fvonvyekztwxw4[51] : fvonvyekztwxw4[52]); 
wire zmr0v5rhc9a6i2_ocf5gsr = mt90aszfju_i2zee | (j384788dhg6btg4 ? mmhfmsr3zdjrk2[22] : mmhfmsr3zdjrk2[23]); 

wire ue06qtglud650ghtx3rja2qw = atm4upf52hg3l87yr ? t_t7vy1dpix0yv7cp[51] : t_t7vy1dpix0yv7cp[52];
wire ld7oztlybql21_i8z999dw = j384788dhg6btg4 ? uo557q_42160ch[22] : uo557q_42160ch[23];

wire n4uew15tqtrctk4ucjxbd6 = (~v0k68izxc00gi8fsnfdw3rars6);
wire ojdi_fe_n7vgpm43st = (~zmr0v5rhc9a6i2_ocf5gsr);

wire g_awm2kdbu3xwua3s5h3lm = (~ue06qtglud650ghtx3rja2qw) & (ugxsstwfs7ud2ujj76==13'b1);
wire d5pok3w4j712te3kg = (~ld7oztlybql21_i8z999dw) & (ugxsstwfs7ud2ujj76==13'b1);

wire [51:0] dd3wknjfiqcua5zo47 = atm4upf52hg3l87yr ? {fvonvyekztwxw4[50:0],ckpku1ypqvuy811tcixg} : fvonvyekztwxw4[51:0]; 
wire [22:0] dkblcqwfc3rgjt = j384788dhg6btg4 ? {mmhfmsr3zdjrk2[21:0],yf80w6zpsarvnsrd5cnj3etc} : mmhfmsr3zdjrk2[22:0]; 

wire [12:0] vxmmbs2zogdgdg1a9w6= (n4uew15tqtrctk4ucjxbd6) ? 13'b0 :( 
                                  ({13{atm4upf52hg3l87yr}} & rlmpudbadjn3njp6t3pg    )
                                | ({13{hq1a13ibszmpmt0aun}} & ivv694h2frwdqy0wg) 
                                | ({13{wy5xxr8o4e6}} & ugxsstwfs7ud2ujj76        )
                             );

wire [12:0] xjmsngtqb2pofjyr62= (ojdi_fe_n7vgpm43st) ? 13'b0 :(
                                 ({13{j384788dhg6btg4}} & rlmpudbadjn3njp6t3pg    )
                               | ({13{mt90aszfju_i2zee}} & ivv694h2frwdqy0wg)
                               | ({13{ox0usqzivjky70}} & ugxsstwfs7ud2ujj76        )
                             );


wire d3k1qwoh84axi739q    = ((|ugxsstwfs7ud2ujj76[12:8]) | (&ugxsstwfs7ud2ujj76[7:0]))  & (~gi2lnto4gl0sc9);
wire gri8ix9g1pbxav6sg9u5    = ((|ugxsstwfs7ud2ujj76[12:11])| (&ugxsstwfs7ud2ujj76[10:0])) & (~gi2lnto4gl0sc9);

wire g7mzxj5gtyr15rwi0j = ((|rlmpudbadjn3njp6t3pg[12:8])  | (&rlmpudbadjn3njp6t3pg[7:0]))  & (~gi2lnto4gl0sc9);
wire z70kxcvmh__193m6hm54 = ((|rlmpudbadjn3njp6t3pg[12:11]) | (&rlmpudbadjn3njp6t3pg[10:0])) & (~gi2lnto4gl0sc9);

wire e_r09ivj7uw6jdsnewaowel = ((|ivv694h2frwdqy0wg[12:8])  | (&ivv694h2frwdqy0wg[7:0]))  & (~gi2lnto4gl0sc9);
wire g0xhc18bxv0d4rde99q = ((|ivv694h2frwdqy0wg[12:11]) | (&ivv694h2frwdqy0wg[10:0])) & (~gi2lnto4gl0sc9);

wire a80_azyei_zb7iz= (atm4upf52hg3l87yr & z70kxcvmh__193m6hm54)     
              |  (hq1a13ibszmpmt0aun & g0xhc18bxv0d4rde99q) 
              |  (wy5xxr8o4e6 & gri8ix9g1pbxav6sg9u5);

wire sx_hyu1_u6skpw= (j384788dhg6btg4 & g7mzxj5gtyr15rwi0j) 
              |  (mt90aszfju_i2zee & e_r09ivj7uw6jdsnewaowel) 
              |  (ox0usqzivjky70 & d3k1qwoh84axi739q);


wire w_nxipv295r = (lh6unwr3hep | rl79o_xu | u2n0m_qrom5l | a80_azyei_zb7iz) & (~gi2lnto4gl0sc9);
wire im2_gxx2wf1 = (ew042ocnt | oy6dz1dkg4cz | v9x3wim2co7eb | sx_hyu1_u6skpw) & (~gi2lnto4gl0sc9);

wire xukc0_vjn4mdb = (g_awm2kdbu3xwua3s5h3lm & (w_nxipv295r) & (~gi2lnto4gl0sc9));
wire u4lrnczx1k51 = (d5pok3w4j712te3kg & (im2_gxx2wf1) & (~gi2lnto4gl0sc9));


wire [7-1:0] iexsh3osgpw30cn9;
assign iexsh3osgpw30cn9[6] = 1'b0 ;
assign iexsh3osgpw30cn9[5]  = 1'b0;
assign iexsh3osgpw30cn9[4]  = im2_gxx2wf1;
assign iexsh3osgpw30cn9[3]  = u4lrnczx1k51;
assign iexsh3osgpw30cn9[2]  = sx_hyu1_u6skpw;
assign iexsh3osgpw30cn9[1]  = 1'b0 ;
assign iexsh3osgpw30cn9[0]  = 1'b0 ;

wire [7-1:0] h8hqm6t244wmwkos;
assign h8hqm6t244wmwkos[6] = 1'b0 ;
assign h8hqm6t244wmwkos[5]  = 1'b0;
assign h8hqm6t244wmwkos[4]  = w_nxipv295r;
assign h8hqm6t244wmwkos[3]  = xukc0_vjn4mdb;
assign h8hqm6t244wmwkos[2]  = a80_azyei_zb7iz;
assign h8hqm6t244wmwkos[1]  = 1'b0 ;
assign h8hqm6t244wmwkos[0]  = 1'b0 ;

assign br_f61q6qczmz8 = (o6xo7iacb14nta9 ? gcl5p_j91agj :iexsh3osgpw30cn9);
assign ttnbtbp7drj = (o6xo7iacb14nta9 ? gcl5p_j91agj :h8hqm6t244wmwkos);

wire wgsc2tqzny = gi2lnto4gl0sc9 ? co3mgjjdm6kydzn01y2wdjd : oystrf6qb5s0k8;

wire hk695dd9rzq_4e = (gi2lnto4gl0sc9) & (~o6xo7iacb14nta9);
wire gh6qttj1pq3bhe08 = (gi2lnto4gl0sc9) & (~o6xo7iacb14nta9);

wire fj1yluer7kh = sx_hyu1_u6skpw & (
                   (ach5cwxikdp == 3'b000) 
                 | (ach5cwxikdp == 3'b100)
                 | ( oystrf6qb5s0k8 & (ach5cwxikdp == 3'b10))
                 | (~oystrf6qb5s0k8 & (ach5cwxikdp == 3'b11))
                ) & (~o6xo7iacb14nta9);

wire g8y1_xip90dr = a80_azyei_zb7iz & (
                   (ach5cwxikdp == 3'b000) 
                 | (ach5cwxikdp == 3'b100)
                 | ( oystrf6qb5s0k8 & (ach5cwxikdp == 3'b10))
                 | (~oystrf6qb5s0k8 & (ach5cwxikdp == 3'b11))
                ) & (~o6xo7iacb14nta9);

wire k2j4gc3kgtl84 =sx_hyu1_u6skpw & (
                             (ach5cwxikdp==3'b01)
                           | ( oystrf6qb5s0k8 & (ach5cwxikdp == 3'b11))
                           | (~oystrf6qb5s0k8 & (ach5cwxikdp == 3'b10))
                          ) & (~o6xo7iacb14nta9);

wire qllbkpzwfl8ak = a80_azyei_zb7iz & (  
                             (ach5cwxikdp == 3'b01)
                           | ( oystrf6qb5s0k8 & (ach5cwxikdp == 3'b11))
                           | (~oystrf6qb5s0k8 & (ach5cwxikdp == 3'b10))
                          ) & (~o6xo7iacb14nta9);

wire tvyothg8mrryb7oy = (gh6qttj1pq3bhe08 | fj1yluer7kh | k2j4gc3kgtl84 | o6xo7iacb14nta9);
wire khmfdx6fcnt6_z = (hk695dd9rzq_4e | g8y1_xip90dr | qllbkpzwfl8ak | o6xo7iacb14nta9);

wire[63:0] aoxd23svi2153u = ({64{hk695dd9rzq_4e}} & {wgsc2tqzny,3'b000, 60'h000000000000000}) 
                       | ({64{g8y1_xip90dr}} & {oystrf6qb5s0k8,3'b111,60'hff0000000000000}) 
                       | ({64{qllbkpzwfl8ak}} & {oystrf6qb5s0k8,3'b111,60'hfefffffffffffff})
                       | ({64{o6xo7iacb14nta9}} & {fjo4qiwyjs8,pfbn0r50hqi});

wire[31:0] laovtnt4fep = ({32{gh6qttj1pq3bhe08}} & {wgsc2tqzny,3'b000, 28'h0000000}) 
                       | ({32{fj1yluer7kh}} & {oystrf6qb5s0k8,3'b111,28'hf800000}) 
                       | ({32{k2j4gc3kgtl84}} & {oystrf6qb5s0k8,3'b111,28'hf7fffff}) 
                       | ({32{o6xo7iacb14nta9}} & pfbn0r50hqi);

assign ejo3ojh7m47_vp7sji6u_1 = (khmfdx6fcnt6_z ? aoxd23svi2153u : {oystrf6qb5s0k8,vxmmbs2zogdgdg1a9w6[10:0],dd3wknjfiqcua5zo47[51:0]});
assign ei1aqk1e3hxolgk4w5xi_ = (tvyothg8mrryb7oy ? laovtnt4fep : {oystrf6qb5s0k8,xjmsngtqb2pofjyr62[ 7:0],dkblcqwfc3rgjt[22:0]}); 


wire [6-1:0] kzswwpy14fd;
wire [32-1:0] sqax;
wire [32-1:0] p7mp;

wire [32-1:0] cks72w2dfx = wo1nm8zgf6 ? ejo3ojh7m47_vp7sji6u_1[31:00] : ei1aqk1e3hxolgk4w5xi_[31:0];
wire [32-1:0] hn1twhx_e_ = ejo3ojh7m47_vp7sji6u_1[63:32] ;
wire [ 6-1:0] w1x194igcmc_xp = wo1nm8zgf6 ? ttnbtbp7drj[5:0] : br_f61q6qczmz8[5:0];

    localparam jomrtsbx11r1wra7a4vh9uu = 1'b0; 
    localparam wwd9tvhgk1kmgl6gr4iivcm = 1'b1; 
    localparam vn_ecxrltje9136ruzvw5p = 1'b0; 
    localparam rwmxv1tt34liv5y_x1du1v = 1'b1; 
    localparam zmk1gz_q9asrgfy2pfvsqo8j = 1'b1; 
    localparam nbrafm9zuo4qwtazxiu8gntc4 = 1'b0; 
wjr2um7_i8ekzqst54wvn1f0 #(164, vn_ecxrltje9136ruzvw5p) yqpdot5dwc5v52ic313yre3rqk(f4_3ig0unyv0i, cdut53tpwkh302, u_1lz3gy_x6_ha5hckf, gf33atgy, ru_wi) ;
wjr2um7_i8ekzqst54wvn1f0 #(164, vn_ecxrltje9136ruzvw5p) qzzw60bvle_oc9nko6e7hj8njryi(f4_3ig0unyv0i, bpzk76nrkskhqgqeym, mzs3mhha1mu673a02e, gf33atgy, ru_wi) ;
wjr2um7_i8ekzqst54wvn1f0 #(256, vn_ecxrltje9136ruzvw5p) f3jep1u0n7e00r4fhluw7u8(f4_3ig0unyv0i, hzc1y, gzevpqks4ek, gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(8, rwmxv1tt34liv5y_x1du1v) bhdwreu9s3_be08233uyel5( iue_ys441x03e_7n, w770780rlqi6,hlmjo66nn_vl0tc, gf33atgy, ru_wi) ;
wjr2um7_i8ekzqst54wvn1f0 #(163, rwmxv1tt34liv5y_x1du1v)  bomiqxlw8gdnx9l9t34fyv96xy0( iue_ys441x03e_7n, jrdafd333s5adeh15,m_n4zvnbl0boxtgug8, gf33atgy, ru_wi) ;
wjr2um7_i8ekzqst54wvn1f0 #(1, rwmxv1tt34liv5y_x1du1v)  gw_zi9gg_tz8ok44ubhcun23k_al44mv( iue_ys441x03e_7n, ghwsivxem72r_3m__sye,dhjwqosv4ycmcnx50oozvu, gf33atgy, ru_wi) ;
wjr2um7_i8ekzqst54wvn1f0 #(1, zmk1gz_q9asrgfy2pfvsqo8j)  mi_9kntdwo77unt7tjurz0vcr4ew38l4( k5oz5augg717tkto, dhjwqosv4ycmcnx50oozvu,q58jwqackb28ri3ianjbm5, gf33atgy, ru_wi) ;
wjr2um7_i8ekzqst54wvn1f0 #(1, zmk1gz_q9asrgfy2pfvsqo8j) hu2fgpf8q_hqn91b8nubfsr( k5oz5augg717tkto, wxy_rmva3xpos0,oystrf6qb5s0k8, gf33atgy, ru_wi) ;
wjr2um7_i8ekzqst54wvn1f0 #(1, zmk1gz_q9asrgfy2pfvsqo8j)  ae35uvork_awgq9a8m5vzqn2oyov26za6(k5oz5augg717tkto, sq8tpegqmuekghx, w9teop0xh2jhgpg7iq_e, gf33atgy, ru_wi) ;
wjr2um7_i8ekzqst54wvn1f0 #(162, zmk1gz_q9asrgfy2pfvsqo8j)hxb1q7rr3bmjk3493w5cr7dqa3tg       (k5oz5augg717tkto, pf46x9eq8b,        clkxpqou7ir6og       , gf33atgy, ru_wi) ;
wjr2um7_i8ekzqst54wvn1f0 #(13, zmk1gz_q9asrgfy2pfvsqo8j) omny9r3xrhmbrdgg__rgsh2in76     (k5oz5augg717tkto, n0_3jdbndqe18,          ugxsstwfs7ud2ujj76         , gf33atgy, ru_wi) ;
wjr2um7_i8ekzqst54wvn1f0 #(13, zmk1gz_q9asrgfy2pfvsqo8j) alxpmkf_nq84buavxitudqvqxry570q  (k5oz5augg717tkto, gk6mz5clwkmam2g5,       rlmpudbadjn3njp6t3pg      , gf33atgy, ru_wi) ;
wjr2um7_i8ekzqst54wvn1f0 #(13, zmk1gz_q9asrgfy2pfvsqo8j) lzyoc5m96qsl2fjweo2nl0q1xxxc_xk_  (k5oz5augg717tkto, e32ykab5wzwl8tnz,       ivv694h2frwdqy0wg      , gf33atgy, ru_wi) ;
wjr2um7_i8ekzqst54wvn1f0 #(6, zmk1gz_q9asrgfy2pfvsqo8j)  c_nmhlb9bn79mvdh8cqqxserpoj073cbv_zxgfb(k5oz5augg717tkto, xsd5n8eqwh_b0n2vvvcup, j_59k0vdcyzjg4dx9zjnwu1t, gf33atgy, ru_wi) ;

wjr2um7_i8ekzqst54wvn1f0 #(106, jomrtsbx11r1wra7a4vh9uu) xsdresj_2dwh5r4_jag_(e7hmnv0h1u8kjcw, b_0ht, zf2wuu6f, gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(106, jomrtsbx11r1wra7a4vh9uu) s_011ko_4oo8_r9b_dl4eg(e7hmnv0h1u8kjcw, oazfr2ucb, ipmcb4953, gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(106, jomrtsbx11r1wra7a4vh9uu) s9_lqp1eqv5btqxi1kt(e7hmnv0h1u8kjcw, p07jru, vje27h4vio, gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(106, jomrtsbx11r1wra7a4vh9uu) hhkvgpdgurxuct63s25z6yr(e7hmnv0h1u8kjcw, is4rk, skablhb13q, gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(106, jomrtsbx11r1wra7a4vh9uu) jcp8plysfeuji6dp9vhdu(e7hmnv0h1u8kjcw, h5w1j3, cb_65dtz, gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(106, jomrtsbx11r1wra7a4vh9uu) ma0if9l7bs50r8phuj1xpwa2(e7hmnv0h1u8kjcw, vs1z8, mue2czm03, gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(106, jomrtsbx11r1wra7a4vh9uu) ovy0gf0pd6lfukqb7b2j(e7hmnv0h1u8kjcw, hk7neg5b6, apzd3bocb0jlz, gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(106, jomrtsbx11r1wra7a4vh9uu) whmnvmf29clafnikzg_0gkzh(e7hmnv0h1u8kjcw, x_5tn8w, qsofrkqvi, gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(106, jomrtsbx11r1wra7a4vh9uu) tkcy3rsvlvtclvtfq60t(e7hmnv0h1u8kjcw, xdzb4s0ejm, tbqp2_p5b, gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(106, jomrtsbx11r1wra7a4vh9uu) j0ssa99h3b_a94c03l16yr(e7hmnv0h1u8kjcw, tr2ajiq, vask7qpb, gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(106, jomrtsbx11r1wra7a4vh9uu) j72fxy02u28es7pzioq5ea(e7hmnv0h1u8kjcw, f0k2ir301f, vkbk0udu, gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(106, jomrtsbx11r1wra7a4vh9uu) qdur6d5gukqpmscjz5gv80(e7hmnv0h1u8kjcw, n2fm6, y9vjbgehnlld, gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(106, jomrtsbx11r1wra7a4vh9uu) o7ubb5hk92nd_cev6j8udfoc(e7hmnv0h1u8kjcw, cpkrdt, snujns_17o, gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(106, jomrtsbx11r1wra7a4vh9uu) gcojzs3h4fbxkhklvlv(e7hmnv0h1u8kjcw, td137, r49be1odf, gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(106, jomrtsbx11r1wra7a4vh9uu) quocts4cdynzpx2rbz2tc(e7hmnv0h1u8kjcw, kf_ejf, fmmslemj9z9, gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(106, jomrtsbx11r1wra7a4vh9uu) wrztpkdkub0aaqx044pleyn(e7hmnv0h1u8kjcw, olreui, tezkbiwpx10os, gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(106, jomrtsbx11r1wra7a4vh9uu) fxz79lsk0afxrxgs83pv0u2(e7hmnv0h1u8kjcw, nh9i6q51r, ezb1_13jolmi, gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(106, jomrtsbx11r1wra7a4vh9uu) vhejcuzfqqo96a7pgu3yi(e7hmnv0h1u8kjcw, zu59l2mmd, vgfckvnmljw, gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(106, jomrtsbx11r1wra7a4vh9uu) haahd05n84u4rl35zfdm(e7hmnv0h1u8kjcw, dtoeq, ps3bgs1w, gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(106, jomrtsbx11r1wra7a4vh9uu) rk60y51yhz3zsq4cd7_jmc(e7hmnv0h1u8kjcw, m5s6xnj, wbbij0elfpd, gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(106, jomrtsbx11r1wra7a4vh9uu) jp0bgbst_qq5c3ox224ef(e7hmnv0h1u8kjcw, rzu745tt29, vm7box2gikw3, gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(106, jomrtsbx11r1wra7a4vh9uu) utd86x16ggfyouwuxqh(e7hmnv0h1u8kjcw, ca8pgl9, wxqo_7ac7g, gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(106, jomrtsbx11r1wra7a4vh9uu) bo8f_7l8i2ro2oxn3435d(e7hmnv0h1u8kjcw, wqjzd4lir, ufo0585p, gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(106, jomrtsbx11r1wra7a4vh9uu) jm4cbxmoud8sal3hqhvl_a(e7hmnv0h1u8kjcw, aeeu2arrcv, gyh98b_6jowgw, gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(106, jomrtsbx11r1wra7a4vh9uu) ywjsc5jucyo0ojwq84y(e7hmnv0h1u8kjcw, aihp3cuom0, nqh156gtt8f, gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(106, jomrtsbx11r1wra7a4vh9uu) uwj_qo8n95tzzw_6_221rom(e7hmnv0h1u8kjcw, uucty, xjc8hz47unk4, gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(106, jomrtsbx11r1wra7a4vh9uu) bdn7xg_dy8mwggrcjyjymu(e7hmnv0h1u8kjcw, rwnza0fed, crlqmi91i, gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(106, jomrtsbx11r1wra7a4vh9uu) olli8q54jyy4ggfd1i5(e7hmnv0h1u8kjcw, lfm5om4i85, xuugnk6md694i, gf33atgy, ru_wi);

wjr2um7_i8ekzqst54wvn1f0 #(106, wwd9tvhgk1kmgl6gr4iivcm) x_9gqzk8xvbvsbizszwhded(enaanseli0es1, kaxkamth, mknydvsmn87, gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(106, wwd9tvhgk1kmgl6gr4iivcm) j7ybceixk5pe9m4k35jtqu9(enaanseli0es1, vou_g00czb2, ga_yvggsogewp, gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(106, wwd9tvhgk1kmgl6gr4iivcm) nl5_k9zyk6sfgwb3jhuymxl(enaanseli0es1, rbm2min6, z49e6oo_eurd, gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(106, wwd9tvhgk1kmgl6gr4iivcm) edtx318j5x5s9o5d_zsghm(enaanseli0es1, qtui513wjhfz, ttw8izs6, gf33atgy, ru_wi);


wjr2um7_i8ekzqst54wvn1f0 #(1, wwd9tvhgk1kmgl6gr4iivcm) ht9klhzgg91fwcmno08n6aq95xi(    enaanseli0es1, eyrxcj62t1hhlhl5a,    uaj78s2_c4g_oj,    gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(1, wwd9tvhgk1kmgl6gr4iivcm) z865mjfgfegjo2vgs8pxtrjsdsq76( enaanseli0es1, xvkeh6i41ok88w6, qcwfkcu7uqutzlw, gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(1, wwd9tvhgk1kmgl6gr4iivcm) mepxprtqabir8cbid560j1vavl(     enaanseli0es1, cqhijr5kjq47ju8,     txe2dhitn770j9,     gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(1, wwd9tvhgk1kmgl6gr4iivcm) rgrjvfx02vxwmer6alh79m_y8(     enaanseli0es1, t6l_v4h7nke_u10,     why9n7prff549n4,     gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(1, jomrtsbx11r1wra7a4vh9uu)  tu8qb8wyrwnc6sgzdddpt_(       e7hmnv0h1u8kjcw, ust6kl,          k4rju_fn1hu,       gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(1, jomrtsbx11r1wra7a4vh9uu)  pv3f74et9vk1yxsj7bx9(       e7hmnv0h1u8kjcw, sjgen2,          gkh_mqfc5dvc,       gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(1, jomrtsbx11r1wra7a4vh9uu)  pi81bwm73pnf8epph6kl51d(      e7hmnv0h1u8kjcw, yxh7zvljyqqn,         a2iop2r7welh,      gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(1, jomrtsbx11r1wra7a4vh9uu)  jzrylspma8s0ap96hrrvqx(     e7hmnv0h1u8kjcw, wijmhrmp5iul,     rdxa7brdak7c19s6,     gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(1, wwd9tvhgk1kmgl6gr4iivcm) k7p2qehpj0jlcm384awy2tkn(     enaanseli0es1, rdxa7brdak7c19s6,     md5qcqkyg3_k,     gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(13, jomrtsbx11r1wra7a4vh9uu) b0kowpxb8belhsrce3qn8eto(     e7hmnv0h1u8kjcw, skjbk0pfgso_,        j9j9j7etnch5,     gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(13, jomrtsbx11r1wra7a4vh9uu) jyvuswo41hoz2170i_obtj6fupa(     e7hmnv0h1u8kjcw, mx2ztfgr0lzn,        yoysx5qs9zqcbwhf,     gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(13, jomrtsbx11r1wra7a4vh9uu) w4qqc7masy5ko6ch56b0bs(     e7hmnv0h1u8kjcw, lsd7m09orucos,        d7zty5n83hwb7y,     gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(53, jomrtsbx11r1wra7a4vh9uu) ghsmjljids8_peeaqktnv5235i9(     e7hmnv0h1u8kjcw, k6ydoqt3g9,        l9zb_468vzbazfa6,     gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(162+3+53, wwd9tvhgk1kmgl6gr4iivcm) mp1jptl21594ynyou3r_q7f96xlkuvag(enaanseli0es1, miz2cix1hgudijz739rzg95i, e6g87hojha93000xrh57dv, gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(162+3+53, wwd9tvhgk1kmgl6gr4iivcm) cdh80exqlv_rbbcmr6aedkaiuvcua5 (enaanseli0es1, mz1jva589d9eep1m5t,  kfxmkdona0ind3vws9sfkn,  gf33atgy, ru_wi);

wjr2um7_i8ekzqst54wvn1f0 #(4, vn_ecxrltje9136ruzvw5p) u17qu6fye8ftst_javd30bs7alyiy53( f4_3ig0unyv0i, lu_owv4hd65jbek_fpn9r,e_rkipm90ja1ygckb24b, gf33atgy, ru_wi) ;
wjr2um7_i8ekzqst54wvn1f0 #(4, rwmxv1tt34liv5y_x1du1v) zqzvkkqgz6honoaxrl4itajb9pqd8xgtkzsy( iue_ys441x03e_7n, e_rkipm90ja1ygckb24b,iug5igicvl8jmztpzbzfkdvsb, gf33atgy, ru_wi) ;

wjr2um7_i8ekzqst54wvn1f0 #(4, vn_ecxrltje9136ruzvw5p) a3qjt6zo6s8zyeca9l5ugn2c7xfl8qzrn( f4_3ig0unyv0i, stuv4gmzj7bpa1rm9df6woag,vouwjch3wz7_qviomah6acriq, gf33atgy, ru_wi) ;
wjr2um7_i8ekzqst54wvn1f0 #(4, rwmxv1tt34liv5y_x1du1v) nqkz70oksz8_32esbxyor4vtaq0vz5zajt2r4( iue_ys441x03e_7n, vouwjch3wz7_qviomah6acriq,shh3tjbryqx94tx3p0bhj65rap, gf33atgy, ru_wi) ;

wjr2um7_i8ekzqst54wvn1f0 #(1, jomrtsbx11r1wra7a4vh9uu) mqu5zw4myw8vymwp9cmdku( a3q6tl0i5iuy, kp3n0pwlaqgh,ks5rw5y1tx3, gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(1, wwd9tvhgk1kmgl6gr4iivcm) srqom02mwv_phdvq1a_ib( d0evt768bc, mjcsl_c3dwtdp6,kbjfvasuqsn4g, gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(1, vn_ecxrltje9136ruzvw5p) vaz1blo_uefvp9qexcvplugz( xpqt2l625a3, zk65zkc8xko9ebz_,ljz2siay0_, gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(1, rwmxv1tt34liv5y_x1du1v) ep8bm59kh5d2x6uj4xt( ywro5vq2yino, yai82tv8en1jptsp,d0z44bwpp5, gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(1, zmk1gz_q9asrgfy2pfvsqo8j) w8e5itol_ao0nm7e_52vr( e97gdk7jw4ev, sbnvbrzm2242zu82,bop_ca3wk7, gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(32, vn_ecxrltje9136ruzvw5p) v4j8235_nam1fiu3zkab8xd_21c( r1555lotjfob, a_vhiehymx7da1hco,s6102_hpsio4ve, gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(32, rwmxv1tt34liv5y_x1du1v) v21tk7n7wev742fp55vf5xqqq( vsd4e757l2_bb, bn7gxjodtjqv9q5qd,u5gxirwoddu54_, gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(32, zmk1gz_q9asrgfy2pfvsqo8j) x8_jd81266p8z1fcj6iz21( mnchfusd_pal_g, k4x1lk0_vv_0ki1gtj,pfbn0r50hqi, gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(32, vn_ecxrltje9136ruzvw5p) dj0one9s3sab0x2gg5atzwx8zx( iefflu1iikpd9jjc, wdskaz5d6p9ismr1j,bcw8lurc42z, gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(32, rwmxv1tt34liv5y_x1du1v) yh3zpsmuf3ocnu3j10i9jpzvrf( cv8vshys52pxuhd0n, qqbg0l90wg42et,xgs6vgfhby7, gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(32, zmk1gz_q9asrgfy2pfvsqo8j) r1uz64fsasu8psrdxc6ufkxzg( apgiwgv4bubvui1j, qz1zeyajzdmhr5vv6,fjo4qiwyjs8, gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(7, vn_ecxrltje9136ruzvw5p) a2rls04jan9ancxr5ikjl1( r1555lotjfob, a5qzn5s78uj02pe,z80wawc634pnw8u, gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(7, rwmxv1tt34liv5y_x1du1v) uuyd9e0cho5a7khwjhhim( vsd4e757l2_bb, gj0mcve6t3a1peo,xqjlst8d7p1gb, gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(7, zmk1gz_q9asrgfy2pfvsqo8j) llp57zho26rwgezh7ywuoidp43( mnchfusd_pal_g, cv00o83d94urbkwcu,gcl5p_j91agj, gf33atgy, ru_wi);


wjr2um7_i8ekzqst54wvn1f0  #(13, jomrtsbx11r1wra7a4vh9uu) esi92o0_6ku0admufz11b2pr     (e7hmnv0h1u8kjcw, {1'b0,m69yhryw},     v46v_ikm00k,         gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0  #(13, jomrtsbx11r1wra7a4vh9uu) d59blow5popuk1d_yb4qsrkt     (e7hmnv0h1u8kjcw, {1'b0,rhd1sc8doent},     pk01ktquuo1,         gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0  #(13, jomrtsbx11r1wra7a4vh9uu) enms6tp3zcxrlhqty70l69qk     (e7hmnv0h1u8kjcw, {1'b0,zq3hfen},     mlgzk0dlchiy,         gf33atgy, ru_wi);

wjr2um7_i8ekzqst54wvn1f0 #(13, wwd9tvhgk1kmgl6gr4iivcm) n432ha8msvit_sdsktnz7ycw847    (enaanseli0es1, vvtb10ccg215rrzm37t,     not1kzp34m717_xrz3_,     gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0  #(13, vn_ecxrltje9136ruzvw5p) y7r0cficqvskm2tztl9o9l    (f4_3ig0unyv0i, not1kzp34m717_xrz3_,     m4bd_iyv30v8ins0qb,     gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(13, rwmxv1tt34liv5y_x1du1v) smvhgqh7arln7vlp8kf9zfp5pkk    (iue_ys441x03e_7n, m4bd_iyv30v8ins0qb,     duxpze1m6dlz2rx,     gf33atgy, ru_wi);

wjr2um7_i8ekzqst54wvn1f0 #(13, wwd9tvhgk1kmgl6gr4iivcm) nmduxya878sq1w468x76kib     (enaanseli0es1, pa0vxwh5h1zrzt41cf,      u7v1l8233z7v63,      gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0  #(13, vn_ecxrltje9136ruzvw5p) podpc9cypa3zha2ugyevyu3kcq     (f4_3ig0unyv0i, u7v1l8233z7v63,      vfz3yrokggbpc0b1b4,      gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(13, rwmxv1tt34liv5y_x1du1v) r2fnhhuigvxbd2y_vm79v6g0ln     (iue_ys441x03e_7n, vfz3yrokggbpc0b1b4,      crtsq13_r9b5_i8j,      gf33atgy, ru_wi);

wjr2um7_i8ekzqst54wvn1f0 #(13, wwd9tvhgk1kmgl6gr4iivcm) p03fp57ph6vri1nvwfppjlyxe     (enaanseli0es1, bv1krzrvrnk8hdr,      ogkix3lj2m4hbon35a,      gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0  #(13, vn_ecxrltje9136ruzvw5p) x7dhcs2rth1d3xj6en6rl4g     (f4_3ig0unyv0i, ogkix3lj2m4hbon35a,      c5g6edg75opsh985r,      gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(13, rwmxv1tt34liv5y_x1du1v) a5hssevjjtim7isikj98xeq8t     (iue_ys441x03e_7n, c5g6edg75opsh985r,      xrc71n3kb03z2,      gf33atgy, ru_wi);

wjr2um7_i8ekzqst54wvn1f0  #(1, vn_ecxrltje9136ruzvw5p) nam4wmuvwwhkg8lb8mw47y0jy9k (f4_3ig0unyv0i, ri3iascff6a_jektfoqpz1b, aed9k35_92eftqn4tu_nv, gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(1, rwmxv1tt34liv5y_x1du1v) e29c_rqf5ys4xfm_198jsnp96cci (iue_ys441x03e_7n, aed9k35_92eftqn4tu_nv, b7x36_v4z0jlprnsb8vmn2, gf33atgy, ru_wi);


wjr2um7_i8ekzqst54wvn1f0 #(64*2+5, jomrtsbx11r1wra7a4vh9uu) n9gw4kvlef6fsgczh( a3q6tl0i5iuy, m2k7jy,vr7175mt1g,   gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(64*2+5, wwd9tvhgk1kmgl6gr4iivcm) hyt2121spe8shyb0injmy( d0evt768bc, vr7175mt1g,t28xspeeyv, gf33atgy, ru_wi) ;
wjr2um7_i8ekzqst54wvn1f0 #(64*2+5, vn_ecxrltje9136ruzvw5p) z2an52kwp_mwkpkd6l7e( xpqt2l625a3, t28xspeeyv,svl_gmw, gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(64*2+5, rwmxv1tt34liv5y_x1du1v) g172piz9shi1xcr8cbl( ywro5vq2yino, svl_gmw,yef02erc, gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(64*2+5, zmk1gz_q9asrgfy2pfvsqo8j) pmr116eyr89ullb6f6vrf0( e97gdk7jw4ev, yef02erc,myqiiy_cpkk, gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(64*2+5, nbrafm9zuo4qwtazxiu8gntc4) wdaja7kthn8he9amclp( p1xybnd9a, myqiiy_cpkk,p9je8hjc, gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(3, jomrtsbx11r1wra7a4vh9uu) u3u9ybp55bvtfbg7k0wo5f9( a3q6tl0i5iuy, ncf9rmc,dx22d5r9g2vd,     gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(3, wwd9tvhgk1kmgl6gr4iivcm) rt16qq5cp02mtdcs05y68om61( d0evt768bc, dx22d5r9g2vd,dlv8z4devpq45, gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(3, vn_ecxrltje9136ruzvw5p) eamrgujcg8gi_o5oqt56le8( xpqt2l625a3, dlv8z4devpq45,vnqm46gumvwx, gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(3, rwmxv1tt34liv5y_x1du1v) iwf673qhus9mxuaz_fhyp6br( ywro5vq2yino, vnqm46gumvwx,rfxycz8syti7h, gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(3, zmk1gz_q9asrgfy2pfvsqo8j) ga6atmffsvxu84i7du_5dh15( e97gdk7jw4ev, rfxycz8syti7h,ach5cwxikdp, gf33atgy, ru_wi);

wjr2um7_i8ekzqst54wvn1f0 #(1, jomrtsbx11r1wra7a4vh9uu) mlc4wlz5hm_bhzae_6zv( a3q6tl0i5iuy, utngq,m7s5rkmh,     gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(1, wwd9tvhgk1kmgl6gr4iivcm) rmf_ul1770x7dysjum2( d0evt768bc, m7s5rkmh,gma5v70c, gf33atgy, ru_wi) ;
wjr2um7_i8ekzqst54wvn1f0 #(1, vn_ecxrltje9136ruzvw5p) ezm_tpxm9syegize863( xpqt2l625a3, gma5v70c,mb8pmo37pwn, gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(1, rwmxv1tt34liv5y_x1du1v) h5wpz3flxw8am6c0fkm01f( ywro5vq2yino, mb8pmo37pwn,nftpir1zs, gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(1, zmk1gz_q9asrgfy2pfvsqo8j) s6xwp8jiwnv0wg3wat1( e97gdk7jw4ev, nftpir1zs,wo1nm8zgf6, gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(1, nbrafm9zuo4qwtazxiu8gntc4) dbrdqztg7qkl88sk4y( p1xybnd9a, wo1nm8zgf6,mj9r0qdcj, gf33atgy, ru_wi);

wjr2um7_i8ekzqst54wvn1f0 #(18, wwd9tvhgk1kmgl6gr4iivcm) koinfs8fk_ecfgkjfbz28( d0evt768bc, ygvkqdhr3wl,u5_4mgyu0a, gf33atgy, ru_wi) ;
wjr2um7_i8ekzqst54wvn1f0 #(18, vn_ecxrltje9136ruzvw5p) b2a22neevsb27tmjjj46mzf( xpqt2l625a3, u5_4mgyu0a,s7nm7w5ep2a, gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(18, rwmxv1tt34liv5y_x1du1v) bqe9dhjhleig2ckjdk5s( ywro5vq2yino, s7nm7w5ep2a,a28ll7e7x, gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(18, zmk1gz_q9asrgfy2pfvsqo8j) sk8gdadzomnhqqh_t0e( e97gdk7jw4ev, a28ll7e7x,tsz7elf8cv, gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(18, nbrafm9zuo4qwtazxiu8gntc4) fefv0hrmuumovxqfzl3w( p1xybnd9a, tsz7elf8cv,m_qz0i0513, gf33atgy, ru_wi);

wjr2um7_i8ekzqst54wvn1f0 #(1, jomrtsbx11r1wra7a4vh9uu) uh1h7mkm1105ck3_tgv8w_js8e( a3q6tl0i5iuy, ktomwnwy0sxt8v,tqert0u9oxp5tq2j7f,     gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(1, wwd9tvhgk1kmgl6gr4iivcm) i5e8ut49me_ifqxyd97h3k5i_da5y( d0evt768bc, tqert0u9oxp5tq2j7f,dg4dhucjpo5xzo4_qpxw, gf33atgy, ru_wi) ;
wjr2um7_i8ekzqst54wvn1f0 #(1, vn_ecxrltje9136ruzvw5p) h7geuz6zut0kz2z82bpekih5ekjjv( xpqt2l625a3, dg4dhucjpo5xzo4_qpxw,g3izwxx_mo1ghg7, gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(1, rwmxv1tt34liv5y_x1du1v) d0yz8nh5gvijgnbbabg2fm42ulxug( ywro5vq2yino, g3izwxx_mo1ghg7,gc7v9_vi47psze_7640t, gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(1, zmk1gz_q9asrgfy2pfvsqo8j) hx5z55i_8b16i8av8sa733fl4319( e97gdk7jw4ev, gc7v9_vi47psze_7640t,j1l5j73k_gend8nlm, gf33atgy, ru_wi);

wjr2um7_i8ekzqst54wvn1f0 #(1, jomrtsbx11r1wra7a4vh9uu) g_wsv9zxufdohwbloobyk98c( a3q6tl0i5iuy, b1t_fvsbzg,hfzrr01xek2w6k6q8,     gf33atgy, ru_wi);

wjr2um7_i8ekzqst54wvn1f0 #(1, jomrtsbx11r1wra7a4vh9uu) dhx99ci3sv7gp444qupp3rbz34z9fwi( a3q6tl0i5iuy, ift60y9fnl2pw,zh45pxgz_p2t5jp0u,     gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(1, wwd9tvhgk1kmgl6gr4iivcm) fbzrph3bosz_guwohud1gk7v2_efq( d0evt768bc, zh45pxgz_p2t5jp0u,j_af3lmvq39fmm38, gf33atgy, ru_wi) ;
wjr2um7_i8ekzqst54wvn1f0 #(1, vn_ecxrltje9136ruzvw5p) eevlhap5oclo1v2qtzoquztl1e4f4( xpqt2l625a3, j_af3lmvq39fmm38,vstyiobwn29fmatxc53, gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(1, rwmxv1tt34liv5y_x1du1v) itn43d2i1hay7soiq372qyc21238( ywro5vq2yino, vstyiobwn29fmatxc53,l8dp94mozhdlxmr43, gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(1, zmk1gz_q9asrgfy2pfvsqo8j) ey8te4o0gcp39dkv0mpzd0kdzs21u( e97gdk7jw4ev, l8dp94mozhdlxmr43,x_vjfqyby9ywowiy2u3, gf33atgy, ru_wi);

wjr2um7_i8ekzqst54wvn1f0 #(1, jomrtsbx11r1wra7a4vh9uu) kwvooixkzy1a7vk3ydn1il3lbe0( e7hmnv0h1u8kjcw, el96tsan45rrpod0r,yunzqdsnvu2whivp,     gf33atgy, ru_wi) ;
wjr2um7_i8ekzqst54wvn1f0 #(1, wwd9tvhgk1kmgl6gr4iivcm) htjsgy2gs1br0z34j0i0qafi7as5( enaanseli0es1, yunzqdsnvu2whivp,t5bfoq7ke3iipt_2, gf33atgy, ru_wi) ;
wjr2um7_i8ekzqst54wvn1f0 #(1, vn_ecxrltje9136ruzvw5p) di8oxbzk6a0z3ee1i7d9w3ozkg5( f4_3ig0unyv0i, t5bfoq7ke3iipt_2,p4n5_8jz95lf5a_, gf33atgy, ru_wi) ;
wjr2um7_i8ekzqst54wvn1f0 #(1, rwmxv1tt34liv5y_x1du1v) bliyyrbovz_fegxu1ngqk5f2zfoxxql( iue_ys441x03e_7n, p4n5_8jz95lf5a_,sk_hgye1w_624w_, gf33atgy, ru_wi) ;
wjr2um7_i8ekzqst54wvn1f0 #(1, zmk1gz_q9asrgfy2pfvsqo8j) innby01ks655lm1xsr5eaamreni( k5oz5augg717tkto, sk_hgye1w_624w_,m6wrb1i20poe2z7_wtnk, gf33atgy, ru_wi) ;

wjr2um7_i8ekzqst54wvn1f0 #(1, jomrtsbx11r1wra7a4vh9uu) sxreukw2a38yxj1vzu1vg3zkspzltf( e7hmnv0h1u8kjcw, w628i27t5rsmxho,dcd4ih54y76fim,     gf33atgy, ru_wi) ;
wjr2um7_i8ekzqst54wvn1f0 #(1, wwd9tvhgk1kmgl6gr4iivcm) ajuj7ycychmhkpeae6arj4g8go( enaanseli0es1, dcd4ih54y76fim,cfyrb77ier93zex, gf33atgy, ru_wi) ;
wjr2um7_i8ekzqst54wvn1f0 #(1, vn_ecxrltje9136ruzvw5p) m6k7m8zge09z7ki4k9rd2bb24alvn1( f4_3ig0unyv0i, cfyrb77ier93zex,bw5l8ov4grr29galln, gf33atgy, ru_wi) ;
wjr2um7_i8ekzqst54wvn1f0 #(1, rwmxv1tt34liv5y_x1du1v) js6e7qa3_ask5a5p8oim5e17pn5( iue_ys441x03e_7n, bw5l8ov4grr29galln,nunpqy34d5rby3u2c, gf33atgy, ru_wi) ;
wjr2um7_i8ekzqst54wvn1f0 #(1, zmk1gz_q9asrgfy2pfvsqo8j) dyzbfe5u1ryewf900_2v64zz6u6fu2( k5oz5augg717tkto, nunpqy34d5rby3u2c,x7034mgujddxpm19suz, gf33atgy, ru_wi) ;
                                                                    
wjr2um7_i8ekzqst54wvn1f0 #(1, jomrtsbx11r1wra7a4vh9uu) hllh25_6ak80kz_p626pt1b3eyng( e7hmnv0h1u8kjcw, jlx9c2o3yzo,aq_ibj5uwgvmvpubeu,     gf33atgy, ru_wi) ;
wjr2um7_i8ekzqst54wvn1f0 #(1, wwd9tvhgk1kmgl6gr4iivcm) kqrknqfgez_o1ii8bcahz06tn( enaanseli0es1, aq_ibj5uwgvmvpubeu,uzw0q1vxxy2cg, gf33atgy, ru_wi) ;
wjr2um7_i8ekzqst54wvn1f0 #(1, vn_ecxrltje9136ruzvw5p) b7dnwfo1vxx8auvff9vujdvjt( f4_3ig0unyv0i, uzw0q1vxxy2cg,dg5d0rszkwioqupp, gf33atgy, ru_wi) ;
wjr2um7_i8ekzqst54wvn1f0 #(1, rwmxv1tt34liv5y_x1du1v) biop1kj9nbffbf7i25_hgex8d801( iue_ys441x03e_7n, dg5d0rszkwioqupp,eoqybvzdtc5hh, gf33atgy, ru_wi) ;
wjr2um7_i8ekzqst54wvn1f0 #(1, zmk1gz_q9asrgfy2pfvsqo8j) ojpeb9uw53c39tbrm9sy6qzm( k5oz5augg717tkto, eoqybvzdtc5hh,n75p3l63agiq3tuy, gf33atgy, ru_wi) ;

wjr2um7_i8ekzqst54wvn1f0 #( 6, nbrafm9zuo4qwtazxiu8gntc4) rapss6b5k3mp6gy2zamv(p1xybnd9a, w1x194igcmc_xp, kzswwpy14fd, gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(32, nbrafm9zuo4qwtazxiu8gntc4) rd4b9cusrzefed4h2(p1xybnd9a, cks72w2dfx, sqax, gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(32, nbrafm9zuo4qwtazxiu8gntc4) bwhl0udyl3iwnsdupp(p1xybnd9a, hn1twhx_e_, p7mp, gf33atgy, ru_wi);

assign ve6waju1kxdtbu     = (~mj9r0qdcj) ? 32'hFFFFFFFF : p7mp ;
assign ynvgxkg9tf     = sqax ;
assign odq8ih2_pvx_6    = mj9r0qdcj;
assign g2gmxy0taet_c61t   = (kzswwpy14fd[5:0]) ;

endmodule



module b6d95x1xv7_zr3t2ebk (
  input hfzrr01xek2w6k6q8,
  input tqert0u9oxp5tq2j7f,
  input dg4dhucjpo5xzo4_qpxw,
  input uaeb8t1ovp,
  input y18h0qaenz,
  input [31:0] u49yq8sp,
  input [31:0] g91ks,
  input [31:0] ahdfbec41y,
  input [31:0] b04cwa,
  input [31:0] fwknegmn,
  input [31:0] pu0_qq,
  input [2:0] dx22d5r9g2vd ,
  input utngq ,
  input m7s5rkmh ,
  input gma5v70c ,
  
  output t8nr0xyjm88kch7l,
  output ckwgdt4l67va,
  output t6bx6zcifoc03dk,
  output fv3vyybkh98eba,
  output auj_3mt9a3wlbcyh,
  output g3ubkkn59kc,
  
  output fhqh1rdjxepeirvc1,
  output oxnijj3cb_5w,
  output ag79ahc9003tjfw,
  output hyp1jmmm6umhihlz,
  output e5g0gz5pr513gc,
  output iaoj1beeb4un1,
  
  output qxbi5ya_x3iyq,
  output ow9a1nk6tcubsc0,
  output zn79hxvf49003,
  output vur92j3awscoy3c,
  output clk6_twfdf0y,
  output l7t9rpi03xnwcm,
  
  output nxirove5d1 ,
  output oxto21kj774l,
  output [31:0] acl1oms948eb26 ,
  output [31:0] t0wz63jpdmeq4e ,
  output [7-1:0] gzvyqzlwpz ,
  
  input kxfk1t4l2_39m7a7,
  input su7v8qw44q19,
  input ru_wi ,
  input gf33atgy  
  );


wire [31:0] mt0bi3g2wl_2;
wire [31:0] h689l51bk2k;

wire [31:0] b_rhlgz0cfwhf;
wire [31:0] n9tamm9rbvvd2;

wire [31:0] fpxnvciny4_je;
wire [31:0] lqa8ikv0j187;

wire a6kqj451bde_m9da;
wire lpq2v4qkyqwiqpk1;
wire o3t1dji3a613j_eg;

wire t36cy3ns2ez3o;
wire lmho8xlq6q0h1a;
wire zt2d4a4gr9ofq9w;

wire zt6rqsdhqw7;
wire d7hx9zg2wjjjv3;
wire taq_q07z9hph4lm;

wire a5awpldu3sw;
wire i7bly_eqd;
wire x33dmi0y5f;

wire b24ef5xnoqv_a46g2j;
wire hjlyfppei9kyzcapr;
wire nokg86mpgq__4694sz;
wire tyej7yh8gfcvs4dj1w  ;
wire r2biwz6ygpji3__ncb ;
wire e0jzbq9orhjkou9a;
wire k9vwrysqc_d2cn33;
wire woakhpb63o446mm22w1y;
wire nw92wf7xmkgeosan2n;
wire ntgyshbri715o;
wire ujp1gamygxctzf;
wire ukg68tnxk0h;
wire f_mfwjqmhcwre1vb;
wire x6epzzn2duf6wiq;
wire ukki6iv4rlzm8_rrgid0;
wire e536oan25joqghkgc;

wire [31:0] kjid_zdh41d;
wire [31:0] spxgcbmn;

wire [31:0] st3n5qhz5;
wire [31:0] et5qcvg1;
wire [31:0] lmvgg9tgob;
wire [31:0] pzenmagq6d;


wire ykyxq88ejhnm6z = utngq ? (u49yq8sp[30:20] == 11'h7FF) : (g91ks[30:23] == 8'hFF);
wire w4b2rs6pj6ol3 = utngq ? (ahdfbec41y[30:20] == 11'h7FF) : (b04cwa[30:23] == 8'hFF);
wire lhkgv064wpt039f17 = utngq ? (fwknegmn[30:20] == 11'h7FF) : (pu0_qq[30:23] == 8'hFF);
wire i48mlnnyzur     = utngq ? (u49yq8sp[30:20] == 11'h000) : (g91ks[30:23] == 8'h00);
wire td1glnmfo2     = utngq ? (ahdfbec41y[30:20] == 11'h000) : (b04cwa[30:23] == 8'h00);
wire fut03jb6c4     = utngq ? (fwknegmn[30:20] == 11'h000) : (pu0_qq[30:23] == 8'h00);
wire exiyz1djym8k      = utngq ? ({u49yq8sp[19:0],g91ks} == 52'b0) : (g91ks[22:0] == 23'b0);
wire plon1c5v      = utngq ? ({ahdfbec41y[19:0],b04cwa} == 52'b0) : (b04cwa[22:0] == 23'b0);
wire m23r0kqbby      = utngq ? ({fwknegmn[19:0],pu0_qq} == 52'b0) : (pu0_qq[22:0] == 23'b0);
wire b284for6       = i48mlnnyzur & ~exiyz1djym8k;
wire uojp70       = td1glnmfo2 & ~plon1c5v;
wire y2vvp2k7       = fut03jb6c4 & ~m23r0kqbby;

assign nxirove5d1 = (fut03jb6c4 & m23r0kqbby);

wire b3sg1s11lhapi4q = m7s5rkmh ? h689l51bk2k[19] : mt0bi3g2wl_2[22];
wire ziof6rqvpaefe = m7s5rkmh ? n9tamm9rbvvd2[19] : b_rhlgz0cfwhf[22];
wire oorjhvonl7str = m7s5rkmh ? lqa8ikv0j187[19] : fpxnvciny4_je[22];

wire d0zbta_ht31enzsv8 = ~a6kqj451bde_m9da & (~t36cy3ns2ez3o);
wire heiexihf5s0k7 = ~lpq2v4qkyqwiqpk1 & (~lmho8xlq6q0h1a);
wire c37f4710eknce = ~o3t1dji3a613j_eg & (~zt2d4a4gr9ofq9w);

assign t8nr0xyjm88kch7l = a6kqj451bde_m9da & (~zt6rqsdhqw7) & (~b3sg1s11lhapi4q);
assign ckwgdt4l67va = lpq2v4qkyqwiqpk1 & (~d7hx9zg2wjjjv3) & (~ziof6rqvpaefe);
assign t6bx6zcifoc03dk = o3t1dji3a613j_eg & (~taq_q07z9hph4lm) & (~oorjhvonl7str);

assign fv3vyybkh98eba = a6kqj451bde_m9da & (~zt6rqsdhqw7) & b3sg1s11lhapi4q;
assign auj_3mt9a3wlbcyh = lpq2v4qkyqwiqpk1 & (~d7hx9zg2wjjjv3) & ziof6rqvpaefe;
assign g3ubkkn59kc = o3t1dji3a613j_eg & (~taq_q07z9hph4lm) & oorjhvonl7str;

wire rgophzfjh0ho = fv3vyybkh98eba | t8nr0xyjm88kch7l;
wire o7iy4_tc2hu65t = auj_3mt9a3wlbcyh | ckwgdt4l67va;
wire rxyy07ikbt = g3ubkkn59kc | t6bx6zcifoc03dk;

wire ril5uexky_bdg9 = a6kqj451bde_m9da & zt6rqsdhqw7;
wire x2jdhp44r0pkrb = lpq2v4qkyqwiqpk1 & d7hx9zg2wjjjv3;
wire xu6v86lgdej = o3t1dji3a613j_eg & taq_q07z9hph4lm;

wire rq4agdh39okdn = (t36cy3ns2ez3o & zt6rqsdhqw7);
wire rb83u6yov8lrz_ = (lmho8xlq6q0h1a & d7hx9zg2wjjjv3);
wire rdxa7brdak7c19s6 = (zt2d4a4gr9ofq9w & taq_q07z9hph4lm);

wire nzuwbec7zp0mo_bx = (t36cy3ns2ez3o & zt6rqsdhqw7) ;
wire joqrj9cv8v26mk2oo5k = (lmho8xlq6q0h1a & d7hx9zg2wjjjv3) ;
wire li4g0y3dl4figakcq0vw4 = (zt2d4a4gr9ofq9w & taq_q07z9hph4lm) ;


wire [5:0] xgxlhpclxbyl={
    d0zbta_ht31enzsv8 ,
    t8nr0xyjm88kch7l ,
    fv3vyybkh98eba ,
    ril5uexky_bdg9 ,
    a5awpldu3sw ,
    nzuwbec7zp0mo_bx };


wire [5:0] k2zdqkj22eh2ia4={
    heiexihf5s0k7 ,
    ckwgdt4l67va ,
    auj_3mt9a3wlbcyh ,
    x2jdhp44r0pkrb ,
    i7bly_eqd ,
    joqrj9cv8v26mk2oo5k };


wire [5:0] nokj_nbrd0q05={
    c37f4710eknce ,
    t6bx6zcifoc03dk ,
    g3ubkkn59kc ,
    xu6v86lgdej ,
    x33dmi0y5f ,
    li4g0y3dl4figakcq0vw4 };

wire dzojfvwrzquzn7d6 = (m7s5rkmh ? h689l51bk2k[31] : mt0bi3g2wl_2[31]) ^ tqert0u9oxp5tq2j7f;
wire ieowm6034zip90t0 = m7s5rkmh ? n9tamm9rbvvd2[31] : b_rhlgz0cfwhf[31];
wire l_jl3if05f9mjl6a = (m7s5rkmh ? lqa8ikv0j187[31] : fpxnvciny4_je[31]) ^ uaeb8t1ovp;

wire xbdga3hmlirn3cewzibd = (m7s5rkmh ? h689l51bk2k[31] : mt0bi3g2wl_2[31]);
wire s7ar_mb5ellso_bve_c6h = m7s5rkmh ? n9tamm9rbvvd2[31] : b_rhlgz0cfwhf[31];
wire pwqonk9822kdltcv = (m7s5rkmh ? lqa8ikv0j187[31] : fpxnvciny4_je[31]);
 
assign fhqh1rdjxepeirvc1 = ril5uexky_bdg9 & (~xbdga3hmlirn3cewzibd);
assign oxnijj3cb_5w = x2jdhp44r0pkrb & (~s7ar_mb5ellso_bve_c6h);
assign ag79ahc9003tjfw = xu6v86lgdej & (~pwqonk9822kdltcv);
assign hyp1jmmm6umhihlz = ril5uexky_bdg9 & xbdga3hmlirn3cewzibd;
assign e5g0gz5pr513gc = x2jdhp44r0pkrb & s7ar_mb5ellso_bve_c6h;
assign iaoj1beeb4un1 = xu6v86lgdej & pwqonk9822kdltcv;

assign qxbi5ya_x3iyq = nzuwbec7zp0mo_bx & (~xbdga3hmlirn3cewzibd);
assign ow9a1nk6tcubsc0 = joqrj9cv8v26mk2oo5k & (~s7ar_mb5ellso_bve_c6h);
assign zn79hxvf49003 = li4g0y3dl4figakcq0vw4 & (~pwqonk9822kdltcv);
assign vur92j3awscoy3c = nzuwbec7zp0mo_bx & xbdga3hmlirn3cewzibd;
assign clk6_twfdf0y = joqrj9cv8v26mk2oo5k & s7ar_mb5ellso_bve_c6h;
assign l7t9rpi03xnwcm = li4g0y3dl4figakcq0vw4 & pwqonk9822kdltcv;


wire u3xqcj_py28df9  = (dzojfvwrzquzn7d6 ^ ieowm6034zip90t0);
wire pbpbgg80uk98rnp9zfx = ((ril5uexky_bdg9 & rb83u6yov8lrz_) | (x2jdhp44r0pkrb & rq4agdh39okdn));
wire yoxk7st79jftwmt_o2 = t8nr0xyjm88kch7l | (fv3vyybkh98eba & (~ckwgdt4l67va));
wire p19wl_tr43pzf7imv = (~t8nr0xyjm88kch7l & ckwgdt4l67va) | (~rgophzfjh0ho & o7iy4_tc2hu65t) ;

wire ienp93w9y35f9r25  = (~rgophzfjh0ho) & (~o7iy4_tc2hu65t) & (~pbpbgg80uk98rnp9zfx) &
                      (~rq4agdh39okdn) & (~rb83u6yov8lrz_) & (ril5uexky_bdg9 | x2jdhp44r0pkrb);

wire ih_33hnmrd1x25wm = (~rgophzfjh0ho) & (~o7iy4_tc2hu65t) & (~pbpbgg80uk98rnp9zfx) &
                      (rq4agdh39okdn | rb83u6yov8lrz_);

wire gg8hr1d2zuwtq = (yoxk7st79jftwmt_o2 & dzojfvwrzquzn7d6) | (p19wl_tr43pzf7imv & ieowm6034zip90t0) ;

wire nf5_c5h6r7vllybxvuu = gg8hr1d2zuwtq;

wire eb5fqt4uost_16mf = yoxk7st79jftwmt_o2;
wire luq2gbfh0vumhehg = p19wl_tr43pzf7imv;
wire zerc6s7sl7lgz6bfjcaq = pbpbgg80uk98rnp9zfx;
wire h2560eibf5_tuqp9   = ienp93w9y35f9r25 ;
wire nfaghphefo7yy5hs  = ih_33hnmrd1x25wm ;

wire mwgivovgemp = ((u3xqcj_py28df9 & (~pbpbgg80uk98rnp9zfx)));

wire no15q796c2oxnnuxtl = (t8nr0xyjm88kch7l | ckwgdt4l67va) ;

wire vicjxmadg79 = (~(dzojfvwrzquzn7d6 == ieowm6034zip90t0));
wire uukbk_zwab  = (ril5uexky_bdg9 | x2jdhp44r0pkrb);
wire hv39vgxm4phr4 = (rq4agdh39okdn | rb83u6yov8lrz_);

wire ejbhi3rm3nires8 = t6bx6zcifoc03dk;
wire hm7czuadxryogi = (~t6bx6zcifoc03dk) & t8nr0xyjm88kch7l;
wire pogtbc_ke0sv6b4 = (~t6bx6zcifoc03dk) & (~t8nr0xyjm88kch7l) & ckwgdt4l67va;

wire rc3re4a63xpu_yd1cj = (~t6bx6zcifoc03dk) & (~t8nr0xyjm88kch7l) & (~ckwgdt4l67va) & g3ubkkn59kc    
                    & (~((ril5uexky_bdg9 & rb83u6yov8lrz_) | (x2jdhp44r0pkrb & rq4agdh39okdn)));

wire xxjjvbtcrwl359isuj = (~t6bx6zcifoc03dk) & (~t8nr0xyjm88kch7l) & (~ckwgdt4l67va) & (~g3ubkkn59kc) & fv3vyybkh98eba;

wire sfs721gr_3wdz1pu = (~t6bx6zcifoc03dk) & (~t8nr0xyjm88kch7l) & (~ckwgdt4l67va) & (~g3ubkkn59kc) &
                      (~fv3vyybkh98eba) & auj_3mt9a3wlbcyh;

wire runz2969rm9ytn5 = (ejbhi3rm3nires8 | rc3re4a63xpu_yd1cj);
wire na5ta260eufikav = (hm7czuadxryogi | xxjjvbtcrwl359isuj);
wire tu02pqzszv_zv9c2 = (pogtbc_ke0sv6b4 | sfs721gr_3wdz1pu);

wire ab7mi1doeepthr01s = (t6bx6zcifoc03dk | t8nr0xyjm88kch7l | ckwgdt4l67va);
wire am60t4qi0th37rjlc9c6  = (rxyy07ikbt | rgophzfjh0ho | o7iy4_tc2hu65t);

wire ztbzwq0hgbh5o8q7e_t96mxqdft =
    ((ril5uexky_bdg9 & rb83u6yov8lrz_) | (x2jdhp44r0pkrb & rq4agdh39okdn)) & g3ubkkn59kc;

wire f25zu62g51s1ynp22du9nq43= 
    (~am60t4qi0th37rjlc9c6) & 
    ((ril5uexky_bdg9 & rb83u6yov8lrz_) 
      | (rq4agdh39okdn & x2jdhp44r0pkrb) 
      | (xu6v86lgdej & uukbk_zwab & (l_jl3if05f9mjl6a == (~vicjxmadg79))));

wire ot23kox8_pzhv0xe = (ztbzwq0hgbh5o8q7e_t96mxqdft | f25zu62g51s1ynp22du9nq43);

wire z4kutmt0nobh_hi = (~am60t4qi0th37rjlc9c6) & ((xu6v86lgdej & (~l_jl3if05f9mjl6a)) | (uukbk_zwab & (~vicjxmadg79)));
wire mvghsqk7dap4s3qu = (~am60t4qi0th37rjlc9c6) & (~z4kutmt0nobh_hi) & ((xu6v86lgdej & l_jl3if05f9mjl6a) | (uukbk_zwab & vicjxmadg79));

wire t4oq11fuhs57 = (~am60t4qi0th37rjlc9c6) & (~f25zu62g51s1ynp22du9nq43) & (z4kutmt0nobh_hi | mvghsqk7dap4s3qu);

wire bjpwwba6z94w_3 = (~am60t4qi0th37rjlc9c6) & (~f25zu62g51s1ynp22du9nq43) & (~t4oq11fuhs57) & (rdxa7brdak7c19s6 & hv39vgxm4phr4);

wire gm_dirlc3hew6819 = 
     hfzrr01xek2w6k6q8 ? vicjxmadg79 :
     (l_jl3if05f9mjl6a == vicjxmadg79) ? l_jl3if05f9mjl6a : (dx22d5r9g2vd==3'b10);


wire q_te3tclg66qe = (~am60t4qi0th37rjlc9c6)
                 & (~f25zu62g51s1ynp22du9nq43)
                 & (~t4oq11fuhs57)
                 & (~bjpwwba6z94w_3)
                 & (hv39vgxm4phr4);

wire oj_l5oxyqxmeyycvbk = (ot23kox8_pzhv0xe
                    | na5ta260eufikav
                    | tu02pqzszv_zv9c2
                    | runz2969rm9ytn5
                    | t4oq11fuhs57
                    | bjpwwba6z94w_3
                    | q_te3tclg66qe);

wire j113kyg9fv =(ab7mi1doeepthr01s 
               | ztbzwq0hgbh5o8q7e_t96mxqdft
               | f25zu62g51s1ynp22du9nq43 );

wire [7-1:0] mfht_5q8z4r;
assign mfht_5q8z4r[6] = 1'b0;
assign mfht_5q8z4r[5] = 1'b0 ;
assign mfht_5q8z4r[4] = 1'b0 ;
assign mfht_5q8z4r[3] = 1'b0 ;
assign mfht_5q8z4r[2] = 1'b0 ;
assign mfht_5q8z4r[1] = 1'b0 ;
assign mfht_5q8z4r[0] = j113kyg9fv ;

assign oxto21kj774l = (oj_l5oxyqxmeyycvbk);

wire [31:0] spmt41qn9y8c4ow = gma5v70c ? {(spxgcbmn[31]^dg4dhucjpo5xzo4_qpxw), spxgcbmn[30:20], 1'b1, spxgcbmn[18:0]} : 
                         {(spxgcbmn[31] ^ dg4dhucjpo5xzo4_qpxw), spxgcbmn[30:23], 1'b1, spxgcbmn[21:0]} ;
wire [31:0] m470gs4zsmzio89 = gma5v70c ? {kjid_zdh41d[31:0]} :
                         {(kjid_zdh41d[31] ^ dg4dhucjpo5xzo4_qpxw), kjid_zdh41d[30:23], 1'b1, kjid_zdh41d[21:0]} ;

wire [31:0] hp32gsbkr0r56l5 = gma5v70c ? {et5qcvg1[31:20], 1'b1, et5qcvg1[18:0]} : 
                         {et5qcvg1[31:23], 1'b1, et5qcvg1[21:0]} ;
wire [31:0] am7bark1491ab = gma5v70c ? {st3n5qhz5[31:0]} : 
                         {st3n5qhz5[31:23], 1'b1, st3n5qhz5[21:0]} ;

wire [31:0] bgc3eb6ihyzhdzmu = gma5v70c ? {(pzenmagq6d[31]^y18h0qaenz), pzenmagq6d[30:20], 1'b1, pzenmagq6d[18:0]} : 
                         {(pzenmagq6d[31] ^ y18h0qaenz), pzenmagq6d[30:23], 1'b1, pzenmagq6d[21:0]} ;
wire [31:0] kn9p5nbne0a6su5so = gma5v70c ? {lmvgg9tgob[31:0]} : 
                         {(lmvgg9tgob[31] ^ y18h0qaenz),lmvgg9tgob[30:23], 1'b1, lmvgg9tgob[21:0]} ;

wire [32-1:0] e5otgqgjkm78gyd = 32'h7FC00000;
wire [31:0] d5p6z8zb2f0jx4 =
      ({32{e0jzbq9orhjkou9a}} & e5otgqgjkm78gyd ) 
    | ({32{k9vwrysqc_d2cn33}} & e5otgqgjkm78gyd ) 
    | ({32{woakhpb63o446mm22w1y}} & e5otgqgjkm78gyd ) 
    | ({32{nw92wf7xmkgeosan2n}} & e5otgqgjkm78gyd ) 
    | ({32{ntgyshbri715o}} & {ukki6iv4rlzm8_rrgid0, 8'hFF, {23{1'b0}}} )  
    | ({32{ujp1gamygxctzf }} & {e536oan25joqghkgc, 8'h00, {23{1'b0}}} ) 
    | ({32{ukg68tnxk0h }} & {(lmvgg9tgob[31]^y18h0qaenz),lmvgg9tgob[30:0]} ) ;


wire [64-1:0] k7gcz3dfv8 = 64'h7FF80000_00000000;
wire [63:0] xdku8yqh6_4k2q0r0 =
      ({64{e0jzbq9orhjkou9a}} & k7gcz3dfv8 ) 
    | ({64{k9vwrysqc_d2cn33}} & k7gcz3dfv8 ) 
    | ({64{woakhpb63o446mm22w1y}} & k7gcz3dfv8 ) 
    | ({64{nw92wf7xmkgeosan2n}} & k7gcz3dfv8 ) 
    | ({64{ntgyshbri715o}} & {ukki6iv4rlzm8_rrgid0, 11'h7FF, {52{1'b0}}}  ) 
    | ({64{ujp1gamygxctzf }} & {e536oan25joqghkgc, 11'h00, {52{1'b0}}} ) 
    | ({64{ukg68tnxk0h }} & {(pzenmagq6d[31]^y18h0qaenz),pzenmagq6d[30:0],lmvgg9tgob} ) ;


assign t0wz63jpdmeq4e = gma5v70c ? xdku8yqh6_4k2q0r0[63:32] : 32'b0 ;
assign acl1oms948eb26 = gma5v70c ? xdku8yqh6_4k2q0r0[31:00] : d5p6z8zb2f0jx4;

    parameter jomrtsbx11r1wra7a4vh9uu = 1'b0; 
    parameter wwd9tvhgk1kmgl6gr4iivcm = 1'b1; 
    parameter vn_ecxrltje9136ruzvw5p = 1'b0; 
    parameter rwmxv1tt34liv5y_x1du1v = 1'b1; 
    parameter zmk1gz_q9asrgfy2pfvsqo8j = 1'b1; 
    parameter nbrafm9zuo4qwtazxiu8gntc4 = 1'b0; 

wjr2um7_i8ekzqst54wvn1f0 #(32, jomrtsbx11r1wra7a4vh9uu) nmzo32pyvc66wef5gvk(kxfk1t4l2_39m7a7, g91ks, mt0bi3g2wl_2, gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(32, jomrtsbx11r1wra7a4vh9uu) jelbuucaew_cgzlyb8n7t(kxfk1t4l2_39m7a7, u49yq8sp, h689l51bk2k, gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(32, jomrtsbx11r1wra7a4vh9uu) uubni3r18_6sayqvhdajn2u(kxfk1t4l2_39m7a7, b04cwa, b_rhlgz0cfwhf, gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(32, jomrtsbx11r1wra7a4vh9uu) bvaaztbtyba718kqmei9m(kxfk1t4l2_39m7a7, ahdfbec41y, n9tamm9rbvvd2, gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(32, jomrtsbx11r1wra7a4vh9uu) sfg7i6l63phfnpkl2pp_0o(kxfk1t4l2_39m7a7, pu0_qq, fpxnvciny4_je, gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(32, jomrtsbx11r1wra7a4vh9uu) ai53fzlz7hcur2ho_7ahak0g(kxfk1t4l2_39m7a7, fwknegmn, lqa8ikv0j187, gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(1, jomrtsbx11r1wra7a4vh9uu) eyeep_e3rri0fahnlo71hen36oq(kxfk1t4l2_39m7a7, ykyxq88ejhnm6z, a6kqj451bde_m9da, gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(1, jomrtsbx11r1wra7a4vh9uu) t8r5v2uwf1waa4v96sw96z8tyb(kxfk1t4l2_39m7a7, w4b2rs6pj6ol3, lpq2v4qkyqwiqpk1, gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(1, jomrtsbx11r1wra7a4vh9uu) gnnqz2hpob6azeco13vxzbbieujnnd3(kxfk1t4l2_39m7a7, lhkgv064wpt039f17, o3t1dji3a613j_eg, gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(1, jomrtsbx11r1wra7a4vh9uu) y7991x2uy1vhr88g42okei(kxfk1t4l2_39m7a7, i48mlnnyzur, t36cy3ns2ez3o, gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(1, jomrtsbx11r1wra7a4vh9uu) ahwwvqi6hf4wm64jc1e3wdm(kxfk1t4l2_39m7a7, td1glnmfo2, lmho8xlq6q0h1a, gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(1, jomrtsbx11r1wra7a4vh9uu) ij9_l04eczcv_gxk2evus1pd0(kxfk1t4l2_39m7a7, fut03jb6c4, zt2d4a4gr9ofq9w, gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(1, jomrtsbx11r1wra7a4vh9uu) hxg47jdrzzgrbzocg1gf4(kxfk1t4l2_39m7a7, exiyz1djym8k, zt6rqsdhqw7, gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(1, jomrtsbx11r1wra7a4vh9uu) geozx2st936cq6vnjue9z5n(kxfk1t4l2_39m7a7, plon1c5v, d7hx9zg2wjjjv3, gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(1, jomrtsbx11r1wra7a4vh9uu) c9oumub1edawp5wmtu9ram1a(kxfk1t4l2_39m7a7, m23r0kqbby, taq_q07z9hph4lm, gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(1, jomrtsbx11r1wra7a4vh9uu) hbq66srtxpudye4efb_o3c2hz(kxfk1t4l2_39m7a7, b284for6, a5awpldu3sw, gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(1, jomrtsbx11r1wra7a4vh9uu) n1r7m54_sq9r9er1uzgarxi(kxfk1t4l2_39m7a7, uojp70, i7bly_eqd, gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(1, jomrtsbx11r1wra7a4vh9uu) qwl3kax5iakt7gdsh3sh(kxfk1t4l2_39m7a7, y2vvp2k7, x33dmi0y5f, gf33atgy, ru_wi);

wjr2um7_i8ekzqst54wvn1f0 #(32, wwd9tvhgk1kmgl6gr4iivcm) ud6au_cgi6vayel7drfmx0ex(su7v8qw44q19, fpxnvciny4_je, lmvgg9tgob, gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(32, wwd9tvhgk1kmgl6gr4iivcm) xgink5yfz9zc04p184tyoz3a(su7v8qw44q19, lqa8ikv0j187, pzenmagq6d, gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(32, wwd9tvhgk1kmgl6gr4iivcm) jdskcstk76zv39re3f4b(su7v8qw44q19, mt0bi3g2wl_2, kjid_zdh41d, gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(32, wwd9tvhgk1kmgl6gr4iivcm) guhu28y2eykxj18fyxul9g67(su7v8qw44q19, h689l51bk2k, spxgcbmn, gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(32, wwd9tvhgk1kmgl6gr4iivcm) c90ekopwubbbojgwmdpk8dpz(su7v8qw44q19, b_rhlgz0cfwhf, st3n5qhz5, gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(32, wwd9tvhgk1kmgl6gr4iivcm) g39bg7n3vzhf7463zv0wo(su7v8qw44q19, n9tamm9rbvvd2, et5qcvg1, gf33atgy, ru_wi);

wjr2um7_i8ekzqst54wvn1f0 #(7, wwd9tvhgk1kmgl6gr4iivcm) ae2bvfb4f1o4_efu5vwlxig(su7v8qw44q19, mfht_5q8z4r, gzvyqzlwpz, gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(1, wwd9tvhgk1kmgl6gr4iivcm) kgoo8v3yoicb9rpjtzgqafvvvcwu(su7v8qw44q19, eb5fqt4uost_16mf, b24ef5xnoqv_a46g2j, gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(1, wwd9tvhgk1kmgl6gr4iivcm) bp3nhrloqsvsbj7_nz58jv2px2uue2(su7v8qw44q19, luq2gbfh0vumhehg, hjlyfppei9kyzcapr, gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(1, wwd9tvhgk1kmgl6gr4iivcm) y7w7zn3vomnrqd4_jut98ptawv4d48r5(su7v8qw44q19, zerc6s7sl7lgz6bfjcaq, nokg86mpgq__4694sz, gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(1, wwd9tvhgk1kmgl6gr4iivcm) cxjhc3o16q0sgtk_hcnin33seb(su7v8qw44q19, h2560eibf5_tuqp9, tyej7yh8gfcvs4dj1w  , gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(1, wwd9tvhgk1kmgl6gr4iivcm) loz9uduqfi0fp3apkko3mq5oqibtcn(su7v8qw44q19, nfaghphefo7yy5hs, r2biwz6ygpji3__ncb , gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(1, wwd9tvhgk1kmgl6gr4iivcm) a4dg1dyj3nnzjbksy67xr4ys(su7v8qw44q19, ot23kox8_pzhv0xe, e0jzbq9orhjkou9a, gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(1, wwd9tvhgk1kmgl6gr4iivcm) m1t7livs_ovdnd5j9chqmvxyni8rt9(su7v8qw44q19, na5ta260eufikav, k9vwrysqc_d2cn33, gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(1, wwd9tvhgk1kmgl6gr4iivcm) owu0_4ea7qquzw1vk2uir38cg7(su7v8qw44q19, tu02pqzszv_zv9c2, woakhpb63o446mm22w1y, gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(1, wwd9tvhgk1kmgl6gr4iivcm) yu39q9853vqq8enr6i18ydw1sr(su7v8qw44q19, runz2969rm9ytn5, nw92wf7xmkgeosan2n, gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(1, wwd9tvhgk1kmgl6gr4iivcm) kzkscujm7zyqt5btx9x7bp504(su7v8qw44q19, t4oq11fuhs57, ntgyshbri715o, gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(1, wwd9tvhgk1kmgl6gr4iivcm) efxbfrofaen3qxr2fhcpsil4f0(su7v8qw44q19, bjpwwba6z94w_3, ujp1gamygxctzf, gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(1, wwd9tvhgk1kmgl6gr4iivcm) ez0ky3xcoym1i30byu0n1s7v58(su7v8qw44q19, q_te3tclg66qe, ukg68tnxk0h, gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(1, wwd9tvhgk1kmgl6gr4iivcm) itpq8yk0_1w_gbzrus_jv6becmzxh6(su7v8qw44q19, nf5_c5h6r7vllybxvuu, f_mfwjqmhcwre1vb, gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(1, wwd9tvhgk1kmgl6gr4iivcm) c4xl8uyn6e7rbwct6rdd8o(su7v8qw44q19, mwgivovgemp, x6epzzn2duf6wiq, gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(1, wwd9tvhgk1kmgl6gr4iivcm) lr6zkeim0ap2e8gygduyf1pb3d(su7v8qw44q19, mvghsqk7dap4s3qu, ukki6iv4rlzm8_rrgid0, gf33atgy, ru_wi);
wjr2um7_i8ekzqst54wvn1f0 #(1, wwd9tvhgk1kmgl6gr4iivcm) g1kovjgl55_gmhiq476o62a5ng_5(su7v8qw44q19, gm_dirlc3hew6819, e536oan25joqghkgc, gf33atgy, ru_wi);

endmodule






module joupdqm1ityga9jgy(

 
  output  frfkcvpr3s1e,

  
  
  
  
  input  rj9pxiv3u3_pir,
  output b972jgf18d478vs1,

  input  [64-1:0] gurbf_74_clu,
  input  [64-1:0] d1egtw92y1cy,
  input  [64-1:0] h501hw2_6,
  input  [48-1:0] kiw03i3frj1_6,
  input  [4-1:0] lw3kfp2bybej9,
  input  [3-1:0] ndsh540w8qc1oph,

  
  
  
  output ct0b7_gmchg9rz, 
  input  xvcpof07ihp69zc, 
  output [64-1:0] y3a80wegnmcxvkiw09,
  output [5-1:0] qngaib4rx7i91p4y2vv,
  output [4 -1:0] bqcca4rpw2hdc6m1,
  output pjmhhc9l2dpz6y954 , 

  input  gf33atgy,
  input  ru_wi
  );

  
  wire jm8sn97g2 = kiw03i3frj1_6[11:11 ];
  wire zmu_037gb8ee = kiw03i3frj1_6[12:12 ];
  wire rcj3zne6zm = kiw03i3frj1_6[13:13];
  wire zh6xcagzy = kiw03i3frj1_6[14:14];
  wire hm3rl2  = kiw03i3frj1_6[15:15  ];
  wire hebytic  = kiw03i3frj1_6[16:16  ];
  wire zqb12c2vz  = kiw03i3frj1_6[17:17  ];
  wire fsb7d3b  = kiw03i3frj1_6[18:18  ];
  wire j7z6st  = kiw03i3frj1_6[19:19  ];
  wire ely1y4r   = kiw03i3frj1_6[20:20   ];
  wire jnxbsnbaz7   = kiw03i3frj1_6[21:21   ];
  wire zn9ww900k   = kiw03i3frj1_6[22:22   ];

  wire nn8hi7fy9 = kiw03i3frj1_6[23:23];

  wire mua3clml   = hm3rl2; 
  wire h20o6   = hebytic | fsb7d3b | j7z6st | ely1y4r | jnxbsnbaz7 | zn9ww900k; 
  wire b9_ew6   = zqb12c2vz;
  wire j1pdh0m0vwd = rcj3zne6zm;
  wire gj_3wro5 = zh6xcagzy;
  wire h19pbx3g = zmu_037gb8ee | h20o6;
  wire ltfdvur8ps = jm8sn97g2 | mua3clml | b9_ew6;
  
  
  
  
  wire slg6nsvuv = j1pdh0m0vwd | gj_3wro5;
  wire n7fjyanmcz = h19pbx3g  | gj_3wro5;


  assign pjmhhc9l2dpz6y954 = 1'b0; 

  
  wire [64-1:0] rbjhd36ql4z;

  wire [64-1:0] tcck0j = gurbf_74_clu;
  wire [64-1:0] onuou7_ = (mua3clml | h20o6) ? (
                                     nn8hi7fy9 ? 64'h3FF0000000000000 : 64'hFFFFFFFF_3F800000    
                             ) :
                                     d1egtw92y1cy ;
  wire [64-1:0] zyxzjxq6_0 = (mua3clml | h20o6) ? d1egtw92y1cy : b9_ew6 ? 64'b0 : h501hw2_6;
  wire [64-1:0] lnlkxa0j6_sskdk;
  wire [64-1:0] k_k63_2;
  wire [64-1:0] ltzccammu;
  wire [64*2+5-1:0] m2k7jy;
  wire [64*2+5-1:0] z2skz3wz;
  wire msm6acopl7;
  wire x5y3581fh7r;
  wire wx17e ;
  wire ydini_vx ;
  wire ztt7ua0 ;
  assign m2k7jy = {
                   tcck0j,
                   zyxzjxq6_0,
                   fsb7d3b,
                   j7z6st,
                   ely1y4r ,
                   jnxbsnbaz7 ,
                   zn9ww900k  
                 };
  assign {
                   k_k63_2,
                   ltzccammu,
                   msm6acopl7,
                   x5y3581fh7r,
                   wx17e ,
                   ydini_vx ,
                   ztt7ua0  
                 } = z2skz3wz;
  
  wire vipj5v4jp;
  wire [5-1:0] adnx9wgdt2;
  wire i_mp1b_6j232kg;
  wire bu481v83k29d;
  wire asl_urmofi7s;
  wire gh04xjbwykw9wd;
  wire g4rmwbt0yslq;
  wire p7fye2zf1aei;

  wire wfoni28cogo3bhl;
  wire rx_r34dltk5;
  wire rux2i8zs5tg1l;
  wire n2md11vbhgzi;
  wire sslv1dv_v95mes2;
  wire zu56_23__pyx62;

  wire c597cob4z48yqld;
  wire imknll0c6w2vjs;
  wire clexjop8gcyt7i;
  wire ug4q2r7d88wb9_;
  wire ckzjjyyqsk_igo0q;
  wire p23w6dm80pq0;



  wire nyxl3jayn42b;
  wire i0twiyq2wbmlvd6;
  wire ql50zn__j2hmc8re;
  wire ba0penccyqijkya4;


  yik149nqborvh6gofa51 hdj7ensq1ogl49j0njiyy (
    .p0hjj76jp60rmlw (rbjhd36ql4z),
    .bvdcuoqal71qlv60  (adnx9wgdt2),
    .kv4pn5p7ocrk0 (vipj5v4jp),

    .q_qkwqh5r (b9_ew6),
    .ift60y9fnl2pw (n7fjyanmcz),
    .ktomwnwy0sxt8v (slg6nsvuv),
    .upi6iqvpb6svcz (ndsh540w8qc1oph),
    .zmjel5h70(tcck0j),
    .lsgnmve7k1t(onuou7_),
    .jj_j64pej(zyxzjxq6_0),
    .clquq5nu (nn8hi7fy9),

    .nyxl3jayn42b    (nyxl3jayn42b),
    .i0twiyq2wbmlvd6    (i0twiyq2wbmlvd6),
    .ql50zn__j2hmc8re    (ql50zn__j2hmc8re),
    .ba0penccyqijkya4    (ba0penccyqijkya4),

    .m2k7jy       (m2k7jy),
    .z2skz3wz       (z2skz3wz),
    .i_mp1b_6j232kg  (i_mp1b_6j232kg),
    .bu481v83k29d  (bu481v83k29d),
    .asl_urmofi7s  (asl_urmofi7s),
    .gh04xjbwykw9wd  (gh04xjbwykw9wd),
    .g4rmwbt0yslq  (g4rmwbt0yslq),
    .p7fye2zf1aei  (p7fye2zf1aei),

    .wfoni28cogo3bhl  (wfoni28cogo3bhl),
    .rx_r34dltk5  (rx_r34dltk5),
    .rux2i8zs5tg1l  (rux2i8zs5tg1l),
    .n2md11vbhgzi  (n2md11vbhgzi),
    .sslv1dv_v95mes2  (sslv1dv_v95mes2),
    .zu56_23__pyx62  (zu56_23__pyx62),

    .c597cob4z48yqld  (c597cob4z48yqld),
    .imknll0c6w2vjs  (imknll0c6w2vjs),
    .clexjop8gcyt7i  (clexjop8gcyt7i),
    .ug4q2r7d88wb9_  (ug4q2r7d88wb9_),
    .ckzjjyyqsk_igo0q  (ckzjjyyqsk_igo0q),
    .p23w6dm80pq0  (p23w6dm80pq0),

    .gf33atgy           (gf33atgy),
    .ru_wi       (ru_wi) 
);



  wire uw10__8ugrmq = (~(|rbjhd36ql4z[63:32]));
  wire gbgcgcfnfxi = (~(|rbjhd36ql4z[31:0]));

  wire e3o4d7law = vipj5v4jp ? rbjhd36ql4z[63] : rbjhd36ql4z[31];

  wire [31:0] r56lhto7 = rbjhd36ql4z[63:32];
  wire [31:0] yka_eie89ig5s = rbjhd36ql4z[31:0];

  wire pcl9ui9 = vipj5v4jp ? (r56lhto7[30:20] == 11'h000) : (yka_eie89ig5s[30:23] == 8'h00);
  wire poa5nd  = vipj5v4jp ? ({r56lhto7[19:0],yka_eie89ig5s} == 52'b0) : (yka_eie89ig5s[22:0] == 23'b0);

  wire es9vn3z75r = (pcl9ui9 & poa5nd);

  wire a0fg2t9h6tq =  
                  i_mp1b_6j232kg 
                | gh04xjbwykw9wd;

  wire tbgd7r1xno7vm =  
                  asl_urmofi7s 
                | p7fye2zf1aei;

  wire dlosqsis7q80_ =  
                  a0fg2t9h6tq 
                | tbgd7r1xno7vm; 

  wire vtxlcvvq0nvajcrq4 =  
                   (wfoni28cogo3bhl | n2md11vbhgzi) | 
                   (rux2i8zs5tg1l | zu56_23__pyx62) ; 

  wire r5q3i07u_qjv_4rv =  
                   (c597cob4z48yqld & p23w6dm80pq0) | 
                   (clexjop8gcyt7i & ug4q2r7d88wb9_) ; 

  wire [64-1:0] iwp02pcdhcv0_r =
      vipj5v4jp ? 64'h7FF80000_00000000 : 64'hFFFFFFFF_7FC00000;
 
 
 
 
 
 
 
 
  wire [64-1:0] wie8936i2lu2reok65cmt = 
                   ({64{c597cob4z48yqld & p23w6dm80pq0}} & (x5y3581fh7r ? k_k63_2 : ltzccammu)) |
                   ({64{clexjop8gcyt7i & ug4q2r7d88wb9_}} & (x5y3581fh7r ? ltzccammu : k_k63_2)) ; 

  wire [64-1:0] jkr38ajp1z06936xom4 = 
                          wfoni28cogo3bhl ? k_k63_2 : 
                          rux2i8zs5tg1l ? ltzccammu : 
                          n2md11vbhgzi ? ltzccammu : 
                          zu56_23__pyx62 ? k_k63_2 : 64'b0;

  wire [64-1:0] zpgc60ujc9n_ze4p8hu = 
                          wfoni28cogo3bhl ? ltzccammu : 
                          rux2i8zs5tg1l ? k_k63_2 : 
                          n2md11vbhgzi ? k_k63_2 : 
                          zu56_23__pyx62 ? ltzccammu : 64'b0;

  wire [64-1:0] fofnxo6g_lgqgrtmx0 = 
                          (wfoni28cogo3bhl & rux2i8zs5tg1l) ? 64'd1 : 
                          (n2md11vbhgzi & zu56_23__pyx62) ? 64'd1 : 64'd0;

  wire [64-1:0] u08yfy5e6kk5a8 = (~fofnxo6g_lgqgrtmx0) & ((n2md11vbhgzi ) ? 64'd1 : 
                                                              (wfoni28cogo3bhl ) ? 64'd0 :
                                                              (zu56_23__pyx62 ) ? 64'd0 : 
                                                              (rux2i8zs5tg1l ) ? 64'd1 : 64'd0);

  wire [64-1:0] dmjno7nzrlaman = fofnxo6g_lgqgrtmx0 | u08yfy5e6kk5a8;

  wire [64-1:0] ww5sr98mowl5ywq3_ra = 
                   ({64{a0fg2t9h6tq & (~tbgd7r1xno7vm)}} & ltzccammu) |
                   ({64{tbgd7r1xno7vm & (~a0fg2t9h6tq)}} & k_k63_2) | 
                   ({64{a0fg2t9h6tq & tbgd7r1xno7vm}} & iwp02pcdhcv0_r);

  wire [5-1:0] nlcoync4_09qdzukzlg1ldd = ({5{i_mp1b_6j232kg | asl_urmofi7s}} & 5'b10000);

 
 
 
 
 
  wire [5-1:0] hw9ucazaipf6wqinslhyp3qu = 
                 ({5{(ydini_vx | ztt7ua0) & (a0fg2t9h6tq | tbgd7r1xno7vm)}} & 5'b10000) |
                 ({5{(wx17e) & (i_mp1b_6j232kg | asl_urmofi7s)}} & 5'b10000);
  wire [64-1:0] b2tzuhirihknqomwsj = 
                   ({64{a0fg2t9h6tq | tbgd7r1xno7vm}} & 64'b0);

  assign lnlkxa0j6_sskdk = 
             ({64{msm6acopl7}} & (dlosqsis7q80_ ? ww5sr98mowl5ywq3_ra : vtxlcvvq0nvajcrq4 ? zpgc60ujc9n_ze4p8hu : r5q3i07u_qjv_4rv ? wie8936i2lu2reok65cmt : e3o4d7law ? k_k63_2 : ltzccammu)) 
           | ({64{x5y3581fh7r}} & (dlosqsis7q80_ ? ww5sr98mowl5ywq3_ra : vtxlcvvq0nvajcrq4 ? jkr38ajp1z06936xom4 : r5q3i07u_qjv_4rv ? wie8936i2lu2reok65cmt : e3o4d7law ? ltzccammu : k_k63_2)) 
           | ({64{wx17e }} & (dlosqsis7q80_ ? b2tzuhirihknqomwsj : vtxlcvvq0nvajcrq4 ? fofnxo6g_lgqgrtmx0  : es9vn3z75r ? 64'd1 : 64'd0)) 
           | ({64{ydini_vx }} & (dlosqsis7q80_ ? b2tzuhirihknqomwsj : vtxlcvvq0nvajcrq4 ? u08yfy5e6kk5a8  : (e3o4d7law & (~es9vn3z75r)) ? 64'd1 : 64'd0)) 
           | ({64{ztt7ua0 }} & (dlosqsis7q80_ ? b2tzuhirihknqomwsj : vtxlcvvq0nvajcrq4 ? dmjno7nzrlaman  : (e3o4d7law | es9vn3z75r) ? 64'd1 : 64'd0)) 
             ; 

  wire [5-1:0] r0po1i47kks = 
             ({5{msm6acopl7|x5y3581fh7r}} & nlcoync4_09qdzukzlg1ldd) |
             ({5{wx17e|ydini_vx|ztt7ua0}} & hw9ucazaipf6wqinslhyp3qu) ;

  wire ndmoar5d7_k  = msm6acopl7 | x5y3581fh7r | wx17e | ydini_vx | ztt7ua0; 

  assign y3a80wegnmcxvkiw09  = ndmoar5d7_k ? lnlkxa0j6_sskdk : rbjhd36ql4z[64-1:0];
  assign qngaib4rx7i91p4y2vv = ndmoar5d7_k ? r0po1i47kks  : adnx9wgdt2;


  m4df8f44pc8gto0crv amm5wjm012bze0i7a1ikk(
    .rj9pxiv3u3_pir      (rj9pxiv3u3_pir   ),
    .b972jgf18d478vs1    (b972jgf18d478vs1 ),
    .lw3kfp2bybej9     (lw3kfp2bybej9  ),

    .ct0b7_gmchg9rz    (ct0b7_gmchg9rz    ),
    .xvcpof07ihp69zc    (xvcpof07ihp69zc    ),
    .bqcca4rpw2hdc6m1(bqcca4rpw2hdc6m1), 

    .nyxl3jayn42b    (nyxl3jayn42b),
    .i0twiyq2wbmlvd6    (i0twiyq2wbmlvd6),
    .ql50zn__j2hmc8re    (ql50zn__j2hmc8re),
    .ba0penccyqijkya4    (ba0penccyqijkya4),
     
    .frfkcvpr3s1e    (frfkcvpr3s1e),

    .gf33atgy            (gf33atgy),
    .ru_wi          (ru_wi) 
  );
endmodule




module w8pxut7bux607aof8nd6je #(
  parameter onr7l=8 
  )(
   input gf33atgy,
   input ru_wi,
   input bp_c30xz,
   input [onr7l-1:0] ii,
   input [onr7l-1:0] fij51v,
   input [onr7l-1:0] cuzhl9,
   input [onr7l-1:0] oho1e63,
   input [onr7l-1:0] hl69c,
   input [onr7l-1:0] mck7r06,
   output [onr7l-1:0] tsa1sag7  
  );

wire [onr7l-1:0] xu71ol6m;
wire [onr7l-1:0] pzfjpy9cyi;
wire [onr7l-1:0] n_kxkqf4v;
wire [onr7l-1:0] husl7u_7_j3;
wire [onr7l-1:0] hrib5mm9yr;
wire [onr7l-1:0] qfrx77e4yg;
wire [onr7l-1:0] ctog_xjo2ob;
wire [onr7l-1:0] etmlzc7qal0;

j3aa8h4yagvjsr416mg #(onr7l) youaa_7z41aka(.frgfco(ii),     .ii(fij51v),     .fij51v(cuzhl9),     .c(xu71ol6m), .s(pzfjpy9cyi));
j3aa8h4yagvjsr416mg #(onr7l) q_n1ieirpg4rsd(.frgfco(oho1e63),     .ii(hl69c),     .fij51v(mck7r06),     .c(n_kxkqf4v), .s(husl7u_7_j3));
j3aa8h4yagvjsr416mg #(onr7l) vp65y6zi18jrl12r(.frgfco(xu71ol6m ), .ii(pzfjpy9cyi ), .fij51v(n_kxkqf4v ), .c(hrib5mm9yr), .s(qfrx77e4yg));
j3aa8h4yagvjsr416mg #(onr7l) n5dt8y1hqv6jex38(.frgfco(husl7u_7_j3 ), .ii(qfrx77e4yg ), .fij51v(hrib5mm9yr ), .c(ctog_xjo2ob), .s(etmlzc7qal0));

wire [onr7l-1:0] j4_xgi95i0;
wire [onr7l-1:0] mvy2p19o_u;

ux607_gnrl_dffl #(onr7l) dgc7fphr8yy137b(bp_c30xz, ctog_xjo2ob, j4_xgi95i0, gf33atgy, ru_wi) ;
ux607_gnrl_dffl #(onr7l) v3de3jdo4ura_2nr(bp_c30xz, etmlzc7qal0, mvy2p19o_u, gf33atgy, ru_wi) ;

assign tsa1sag7 =(j4_xgi95i0 + mvy2p19o_u);

endmodule


module xh5dey_d_oxo365f0d85q3d #(
  parameter onr7l=64,
  parameter hw3qvr=6
)(
  input [onr7l-1:0] bjh,
  output [hw3qvr-1:0] ht70
);

wire [onr7l-1:0] cvf2uttd2wy;

assign cvf2uttd2wy[onr7l-1] = bjh[onr7l-1];

genvar j;
generate 
 for (j=onr7l-2; j>=0; j=j-1) begin: m_j0ywdyf2
    assign cvf2uttd2wy[j] = (|bjh[onr7l-1:j]);
 end
endgenerate

wire [onr7l-1:0] i = cvf2uttd2wy & {1'b1,~cvf2uttd2wy[onr7l-1:1]};

assign ht70[0]=( i[00] | i[02] | i[04] | i[06] | i[08] |
                i[10] | i[12] | i[14] | i[16] | i[18] |
                i[20] | i[22] | i[24] | i[26] | i[28] |
                i[30] | i[32] | i[34] | i[36] | i[38] |
                i[40] | i[42] | i[44] | i[46] | i[48] |
                i[50] | i[52] | i[54] | i[56] | i[58] |
                i[60] | i[62] );

assign ht70[1]=( i[00] | i[01] | i[04] | i[05] | 
                i[08] | i[09] | i[12] | i[13] | 
                i[16] | i[17] | i[20] | i[21] | 
                i[24] | i[25] | i[28] | i[29] | 
                i[32] | i[33] | i[36] | i[37] |
                i[40] | i[41] | i[44] | i[45] | 
                i[48] | i[49] | i[52] | i[53] | 
                i[56] | i[57] | i[60] | i[61] );

assign ht70[2]=( i[00] | i[01] | i[02] | i[03] | 
                i[08] | i[09] | i[10] | i[11] | 
                i[16] | i[17] | i[18] | i[19] | 
                i[24] | i[25] | i[26] | i[27] | 
                i[32] | i[33] | i[34] | i[35] |
                i[40] | i[41] | i[42] | i[43] | 
                i[48] | i[49] | i[50] | i[51] | 
                i[56] | i[57] | i[58] | i[59] );

assign ht70[3]=( i[00] | i[01] | i[02] | i[03] | i[04] | i[05] | i[06] | i[07] | 
                i[16] | i[17] | i[18] | i[19] | i[20] | i[21] | i[22] | i[23] | 
                i[32] | i[33] | i[34] | i[35] | i[36] | i[37] | i[38] | i[39] | 
                i[48] | i[49] | i[50] | i[51] | i[52] | i[53] | i[54] | i[55] );

assign ht70[4]=( i[00] | i[01] | i[02] | i[03] | i[04] | i[05] | i[06] | i[07] |
                i[08] | i[09] | i[10] | i[11] | i[12] | i[13] | i[14] | i[15] | 
                i[32] | i[33] | i[34] | i[35] | i[36] | i[37] | i[38] | i[39] |
                i[40] | i[41] | i[42] | i[43] | i[44] | i[45] | i[46] | i[47] );

assign ht70[5]=( i[00] | i[01] | i[02] | i[03] | i[04] | i[05] | i[06] | i[07] |
                i[08] | i[09] | i[10] | i[11] | i[12] | i[13] | i[14] | i[15] | 
                i[16] | i[17] | i[18] | i[19] | i[20] | i[21] | i[22] | i[23] |
                i[24] | i[25] | i[26] | i[27] | i[28] | i[29] | i[30] | i[31] );

endmodule


module k_f7ns0a54rui10fjf(
  input [56:0] f02vn4ah,
  input [56:0] gt_sq2dtwcr,
  input [56:0] lxff,
  input [56:0] c2u,
  input v2f5pmhic4,
  input ust6kl,
  input p2yjv_h8o,
  output [56:0] xphx,
  output [56:0] fap75
);
wire [56:0] frgfco;
wire [56:0] ii;

assign frgfco = {f02vn4ah[56-1:0], 1'b0} ;

assign ii [56:1] = gt_sq2dtwcr[56-1:0] ;
assign ii [0] = ust6kl ;

wire [56:0] fij51v = c2u & {57{ust6kl & ~p2yjv_h8o}} 
               | lxff & {57{~ust6kl & ~p2yjv_h8o} } ;

j3aa8h4yagvjsr416mg #(.onr7l(57)) q7bx0z96lxa4m2ew(
      .frgfco(frgfco), 
      .ii(ii), 
      .fij51v(fij51v), 
      .c(fap75),
      .s(xphx)
) ;
endmodule 

module j3rmuwv9gah_ceeqolq8gh(
  input [56:0] j0xu7nslfaf ,
  input [56:0] hh9u1ei_ ,
  input [56:0]  qnj9dtloi3,
  input [56:0]  vetlu9oe6w4uu,
  input [56:0]  bdl76yc6,
  input [56:0]  rpcdbj3xdniw,
  input ust6kl,
  input p2yjv_h8o ,
  input v2f5pmhic4,
  output [56:0] xphx,
  output [56:0] fap75
);

wire [56:0] xb50rkdb = {3'b111, ((~bdl76yc6[56:3] & j0xu7nslfaf[56:3]) | hh9u1ei_[56:3])} ;
wire [56:0] eamkigyzf = {3'b000, ((rpcdbj3xdniw[56:3] & j0xu7nslfaf[56:3]) | hh9u1ei_[56:3])} ;

wire [56:0] o_guu3_gbbxp0w = xb50rkdb ;
wire [56:0] tkh3ul4k7mwyk = eamkigyzf ;

wire [56:0] frgfco;
wire [56:0] ii;

assign frgfco = {qnj9dtloi3[56-1:0], 1'b0} ;

assign ii [56:1] = vetlu9oe6w4uu[56-1:0] ;
assign ii [0] = 1'b0 ;

wire [56:0] oz7_y5 = ust6kl ? o_guu3_gbbxp0w : tkh3ul4k7mwyk ;

wire [56:0] fij51v = oz7_y5 & {57{~p2yjv_h8o}};

j3aa8h4yagvjsr416mg #(.onr7l(57)) aq3g7s7q92egq_k0_(
      .frgfco(frgfco), 
      .ii(ii), 
      .fij51v(fij51v), 
      .c(fap75),
      .s(xphx)
) ;

endmodule








module ur945ax08pidlnz7_o24hdlr (
   output eypswghjg4a5o,
   
   input  yh0oeg399pvwaqg13,

   output jdo6mn_o05686d2cl ,
   input  baefqz_y6q1d7 ,
   output [4-1:0] ju_5ti46ayy7vdw ,

   output cl_ffrx4sh ,
   output bp_c30xz ,
   output rg10e3avkel ,
   output bhmxsiib6 ,
   output vawmftolubc5 ,
   output c6yo0on_3i ,
   output mg9we1s5d77ws ,

   input [4:0] gd2wkhivb2,
   output ilnqntxsop67,
   
   input  vwd0ug0ks5l ,
   output am_rltp_3w ,
   input [4-1:0] p_rmwvx8z ,
   input uu3yswtakfh,
   input y7s8lz156ibl,

   output q02bklc,
   output nv_meva_f5,
   output lzbquud,
   output y_zx8qolynd,
   output ux0s4l13o,
   
   input gf33atgy ,
   input ru_wi
);

  wire [4-1:0] cc3ge9cz7;
  wire [4-1:0] aiquiiki8;
  wire [4-1:0] e0p08_7j5;
  wire [4-1:0] qoebaecu92e79;
  wire [4-1:0] ht7rmsqp;

  wire nb1jr8lxfasu;
  wire s_0et5df8n3c;
  wire tvw8333v4r7;
  wire rcg7crpr5469;

  wire vz82rs1jwm_ss4fx;
  wire muuiv46mbw9;
  wire xkf1d_xedftb;
  wire agdfmofemj5l2p49;

  wire tw5jlr32l519o;
  wire o_9hw_8713p4h7z;
  wire il4krkgf7p5cxl;
  wire rxhar6hyxqjwvnz2;

  wire kmacljnxh7lvk5i;
  wire klms6kt2b_obz;
  wire h0wd8tmw_mo7;
  wire dvp51opx0833g;

  wire oigtqtxhcsu;
  wire pzoy0nmzgolij;
  wire zobwulnd9v0c;
  wire gw828d9uqkxqaje;


  ux607_gnrl_pipe_stage # (
    
    
   .CUT_READY(1),
   .DP(1),
   .DW(1)
  ) zq_q7kj7fywyb (
   .i_vld(nb1jr8lxfasu), 
   .i_rdy(s_0et5df8n3c), 
   .i_dat(1'b0),
   .o_vld(tvw8333v4r7), 
   .o_rdy(rcg7crpr5469), 
   .o_dat(),
 
   .clk  (gf33atgy  ),
   .rst_n(ru_wi)  
  ); 
  
  ux607_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(1)
  ) eiq3ggh0jsyp6 (
   .i_vld(vz82rs1jwm_ss4fx), 
   .i_rdy(muuiv46mbw9), 
   .i_dat(1'b0),
   .o_vld(xkf1d_xedftb), 
   .o_rdy(agdfmofemj5l2p49), 
   .o_dat(),
 
   .clk  (gf33atgy  ),
   .rst_n(ru_wi)  
  );

  ux607_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(1)
  ) lt55clin45_ (
   .i_vld(tw5jlr32l519o), 
   .i_rdy(o_9hw_8713p4h7z), 
   .i_dat(1'b0),
   .o_vld(il4krkgf7p5cxl), 
   .o_rdy(rxhar6hyxqjwvnz2), 
   .o_dat(),
 
   .clk  (gf33atgy  ),
   .rst_n(ru_wi)  
  );

  ux607_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(1)
  ) fq7ijeb38_v6 (
   .i_vld(kmacljnxh7lvk5i), 
   .i_rdy(klms6kt2b_obz), 
   .i_dat(1'b0),
   .o_vld(h0wd8tmw_mo7), 
   .o_rdy(dvp51opx0833g), 
   .o_dat(),
 
   .clk  (gf33atgy  ),
   .rst_n(ru_wi)  
  );

  ux607_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(1)
  ) gw200oyqgikg0v3 (
   .i_vld(oigtqtxhcsu), 
   .i_rdy(pzoy0nmzgolij), 
   .i_dat(1'b0),
   .o_vld(zobwulnd9v0c), 
   .o_rdy(gw828d9uqkxqaje), 
   .o_dat(),
 
   .clk  (gf33atgy  ),
   .rst_n(ru_wi)  
  );


  assign nb1jr8lxfasu = vwd0ug0ks5l;
  assign am_rltp_3w    = s_0et5df8n3c;

  wire rjtgb6qfj_;

  wire yugh1j8ln_hxn18mdugn7brp = xkf1d_xedftb | rjtgb6qfj_   |
                               il4krkgf7p5cxl | h0wd8tmw_mo7 | zobwulnd9v0c;

  wire i2s0_vxulj0ph;

  assign vz82rs1jwm_ss4fx = (~i2s0_vxulj0ph) & tvw8333v4r7;

  assign rcg7crpr5469 = 
                
                
                 (i2s0_vxulj0ph & (~yugh1j8ln_hxn18mdugn7brp) & pzoy0nmzgolij)  |  
                
                 ((~i2s0_vxulj0ph) & muuiv46mbw9)  ;  

  assign ilnqntxsop67 = i2s0_vxulj0ph & tvw8333v4r7 & (~yugh1j8ln_hxn18mdugn7brp);

  wire ke2zowu68b;
  wire u8osyypd4og = ke2zowu68b;

  assign tw5jlr32l519o = u8osyypd4og & xkf1d_xedftb;
  assign agdfmofemj5l2p49 = u8osyypd4og & o_9hw_8713p4h7z;

  assign kmacljnxh7lvk5i = il4krkgf7p5cxl;
  assign rxhar6hyxqjwvnz2 = klms6kt2b_obz;

  assign oigtqtxhcsu = (i2s0_vxulj0ph & (~yugh1j8ln_hxn18mdugn7brp) & tvw8333v4r7) | h0wd8tmw_mo7;
  assign dvp51opx0833g = pzoy0nmzgolij;

  assign gw828d9uqkxqaje = baefqz_y6q1d7;

  
  wire e195_h9mxm = nb1jr8lxfasu & s_0et5df8n3c;
  wire cd126jvcmhx = vz82rs1jwm_ss4fx & muuiv46mbw9;
  wire ilrjm2wqau48 = tw5jlr32l519o & o_9hw_8713p4h7z;
  wire yvfzn9cc11s74h = kmacljnxh7lvk5i & klms6kt2b_obz;
  wire i0xaobdc7iq_ = oigtqtxhcsu & pzoy0nmzgolij;
  
  
  
  assign mg9we1s5d77ws =   y7s8lz156ibl  & e195_h9mxm; 
  assign cl_ffrx4sh    = (~y7s8lz156ibl) & e195_h9mxm;
  assign bp_c30xz    = (~i2s0_vxulj0ph) & cd126jvcmhx;
  assign bhmxsiib6    = ilrjm2wqau48;
  assign vawmftolubc5    = yvfzn9cc11s74h;
  assign c6yo0on_3i    = i0xaobdc7iq_;
  
  
  wire [4-1:0] sqvxx0i7d92gx = ilnqntxsop67 ? cc3ge9cz7 : qoebaecu92e79;
  wire byww_uvpsuhkw = ilnqntxsop67 ? q02bklc : y_zx8qolynd;
  
  ux607_gnrl_dfflr #(4) qczvjv_7ny6223javex( e195_h9mxm, p_rmwvx8z ,    cc3ge9cz7, gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(4) zfr1dnozbtsz777r( cd126jvcmhx, cc3ge9cz7,    aiquiiki8, gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(4) s77xw6ck8e34d2me( ilrjm2wqau48, aiquiiki8,    e0p08_7j5, gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(4) ajwzga1ey41yyvii9e( yvfzn9cc11s74h, e0p08_7j5,    qoebaecu92e79, gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(4) gu3_h1avqa8a_v1b7ik( i0xaobdc7iq_, sqvxx0i7d92gx, ht7rmsqp, gf33atgy, ru_wi);
  
  ux607_gnrl_dfflr #(1) in_abkeq_j_llwdhb5( e195_h9mxm, uu3yswtakfh ,    q02bklc, gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1) xlw9u_vkflngtr8a97( cd126jvcmhx, q02bklc,    nv_meva_f5, gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1) zch8zga0frb96o9i6n( ilrjm2wqau48, nv_meva_f5,    lzbquud, gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1) m9t5keerkc36d_5i( yvfzn9cc11s74h, lzbquud,    y_zx8qolynd, gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1) kkuy_1at__pkh4ka9y( i0xaobdc7iq_, byww_uvpsuhkw, ux0s4l13o, gf33atgy, ru_wi);

  ux607_gnrl_dfflr #(1) rnl9n1hic4hho7_  (e195_h9mxm, y7s8lz156ibl, i2s0_vxulj0ph, gf33atgy, ru_wi);

  wire fh60_h952l3kq = bp_c30xz;
  wire wjxl3yibmrr = bhmxsiib6;
  wire uqzfldw8oiv = (fh60_h952l3kq | wjxl3yibmrr);
  wire e039cbo7i3ro = (fh60_h952l3kq | (~wjxl3yibmrr));

  ux607_gnrl_dfflr #(1) sp6s6aj1kxxf9(uqzfldw8oiv , e039cbo7i3ro, rjtgb6qfj_, gf33atgy, ru_wi);

  assign rg10e3avkel = (rjtgb6qfj_ & (~ke2zowu68b));

  wire t1jgrhr93g = (bp_c30xz | rg10e3avkel);
  wire [4:0] qa5i4r05;
  wire [4:0] kxo6gjxjsdo90 = bp_c30xz ? 5'b0 
                      : rjtgb6qfj_ ? (qa5i4r05 + 1'b1)
                      : qa5i4r05;
  
  wire v5413v6titvvqo9f = (bp_c30xz | bhmxsiib6) ? 1'b0
                  : (rjtgb6qfj_ & ((qa5i4r05 == gd2wkhivb2) | yh0oeg399pvwaqg13)) ? 1'b1 
                  : ke2zowu68b;
  
  ux607_gnrl_dfflr #(5) qt6et9tyn634  (t1jgrhr93g   , kxo6gjxjsdo90   , qa5i4r05,   gf33atgy, ru_wi);
  ux607_gnrl_dffr  #(1) eilo1x4kysxho7 (v5413v6titvvqo9f , ke2zowu68b  ,            gf33atgy, ru_wi);
  
  assign ju_5ti46ayy7vdw  = ht7rmsqp;
  assign jdo6mn_o05686d2cl = zobwulnd9v0c;

  assign eypswghjg4a5o = tvw8333v4r7 | yugh1j8ln_hxn18mdugn7brp;

endmodule

    


module jgdiavy4q4l1fecbof09xfij9(
  output [4:0] gd2wkhivb2,
  output [31:0] xptd3f_t3cg5 ,
  output [31:0] r4nxuj5xq_p ,
  output [5:0] g2gmxy0taet_c61t, 
  output yh0oeg399pvwaqg13,
  input [31:0] ie_pkh83p_8 ,
  input [31:0] e3oq_fn1szj61 ,
  input [31:0] r1pjdyql2t19 ,
  input [31:0] wswzu1c4y6et ,
  input [5:0] a0_2x3l9euvn1ixa6,
  input [5:0] dvmjxjsqko9mdgn,
  input m0e2_guluq90ndzyt,
  input tqpavw30 ,
  input kjauvty_w ,
  input j5crtzpyh ,
  input ilnqntxsop67,
  input [63:0] powr,
  input [5:0] ey7de2vqxx,
  input cl_ffrx4sh ,
  input bp_c30xz ,
  input rg10e3avkel ,
  input bhmxsiib6 ,
  input vawmftolubc5 ,
  input c6yo0on_3i ,
  input [2:0] n5900it0gq9hnv ,

  input q02bklc,
  input nv_meva_f5,
  input lzbquud,
  input y_zx8qolynd,
  input ux0s4l13o, 

  input gf33atgy ,
  input ru_wi
);

wire mb75fcy6;
wire op5chmv5;
wire jdnbsmmk7_x9;
wire ka66jgi;
wire bpeajju419;
wire [2:0] hmoqkhn1z1r_z ;
wire [2:0] vy74ohm_7sana1i ;
wire [2:0] muvr3ixctzt7xm ;
wire [2:0] ljxpmbsqoaz ;

wire ymxz08x0;
wire soxc9xw1gp;
wire fvz__7_m;

wire [51:00]i4ia5732yw;

wire [6:0] rvezutl8owb63ik2aznm;

wire [10:0] h1_vm6sos4nriqkv;
wire [10:0] a4meogg6iciznynf;


wire [51:00]dsr2v_ycsx8gw = (q02bklc) ?  {ie_pkh83p_8[19:00], e3oq_fn1szj61} :
                       {e3oq_fn1szj61[22:00], 29'b0} ;
wire [51:00]ohh5oui0c7_sw = (q02bklc) ?  {r1pjdyql2t19[19:00], wswzu1c4y6et} :
                       {wswzu1c4y6et[22:00], 29'b0} ;


wire [10:0] cs118t0ggohu0 = q02bklc ? ie_pkh83p_8[30:20] : {3'b0, e3oq_fn1szj61[30:23]} ;
wire [10:0] yruj_3_m8kmx8 = q02bklc ? r1pjdyql2t19[30:20] : {3'b0, wswzu1c4y6et[30:23]} ;

wire [6:0] j2vilqf6umhqi5cj = {1'b0,a0_2x3l9euvn1ixa6}+(~{1'b0,dvmjxjsqko9mdgn})+1'b1;

wire c6s9w3jn0hb6hlu8 = q02bklc ? ie_pkh83p_8[31] : e3oq_fn1szj61[31] ;
wire f9sel_gzzue0p = q02bklc ? r1pjdyql2t19[31] : wswzu1c4y6et[31] ;
wire tumgwa57fmq     = (c6s9w3jn0hb6hlu8 ^ f9sel_gzzue0p) & (~bpeajju419) ;

ux607_gnrl_dffl #(52) ej5m7cpak6j9n3emp_( bp_c30xz, ohh5oui0c7_sw,i4ia5732yw, gf33atgy, ru_wi) ;
ux607_gnrl_dffl #(11) bexpv42ix4ljbgehwcpz( bp_c30xz, cs118t0ggohu0,h1_vm6sos4nriqkv, gf33atgy, ru_wi) ;
ux607_gnrl_dffl #(11) p36ys77nbx56irpi98vkn( bp_c30xz, yruj_3_m8kmx8,a4meogg6iciznynf, gf33atgy, ru_wi) ;
ux607_gnrl_dffl #(7) mwx7rmqgffi2dllr_4h3_j( bp_c30xz, j2vilqf6umhqi5cj,rvezutl8owb63ik2aznm, gf33atgy, ru_wi) ;
ux607_gnrl_dffl #(1) jb2vg520hqqjrmjwtl( bp_c30xz, tumgwa57fmq,ymxz08x0,  gf33atgy, ru_wi) ;
ux607_gnrl_dffl #(1) utbbpnfgs40__oepmp( bhmxsiib6, ymxz08x0,soxc9xw1gp, gf33atgy, ru_wi) ;
ux607_gnrl_dffl #(1) rerytuhl64s93djaqy( vawmftolubc5, soxc9xw1gp,fvz__7_m, gf33atgy, ru_wi) ;
ux607_gnrl_dffl #(1) k96aigyhamjvtt( cl_ffrx4sh, kjauvty_w,mb75fcy6, gf33atgy, ru_wi) ;
ux607_gnrl_dffl #(1) j8ki25jgiim5x4( bp_c30xz, mb75fcy6,op5chmv5, gf33atgy, ru_wi) ;
ux607_gnrl_dffl #(1) yuzt_sczfb5le7b5( bhmxsiib6, op5chmv5,jdnbsmmk7_x9, gf33atgy, ru_wi) ;
ux607_gnrl_dffl #(1) ze3e_pvijtokd9hc( vawmftolubc5, jdnbsmmk7_x9,ka66jgi, gf33atgy, ru_wi) ;

ux607_gnrl_dffl #(1) yqjzc53wc7zvk( cl_ffrx4sh, j5crtzpyh,bpeajju419,     gf33atgy, ru_wi) ;

ux607_gnrl_dffl #(3) jg7q3ynjtdq99zsv( cl_ffrx4sh, n5900it0gq9hnv,hmoqkhn1z1r_z, gf33atgy, ru_wi) ;
ux607_gnrl_dffl #(3) p9_xcemge8tswownc( bp_c30xz, hmoqkhn1z1r_z,vy74ohm_7sana1i, gf33atgy, ru_wi) ;
ux607_gnrl_dffl #(3) wqqqmt_nblnha17atm( bhmxsiib6, vy74ohm_7sana1i,muvr3ixctzt7xm, gf33atgy, ru_wi) ;
ux607_gnrl_dffl #(3) ralzwkf31br1daal0c3( vawmftolubc5, muvr3ixctzt7xm,ljxpmbsqoaz, gf33atgy, ru_wi) ;




wire [56:0] f02vn4ah ;
wire [56:0] gt_sq2dtwcr ;
wire [56:0] qnj9dtloi3 ;
wire [56:0] vetlu9oe6w4uu ;




wire [56:0] hh9u1ei_ ;
wire [56:0] j0xu7nslfaf ;










wire [56:0] kpgls4tvuy_dq9a, xa5onwxrrff4hh, zbx4klyjkjk_39m, e9s410oe7si, ukt_9nlhm1d82lf;




wire [56:0] cwpbbg1e2nj0_4, akr00lq3hfph, auu79qzp63t0_cc0ru, qng6_z6rdlwu3, nm2k_djs2vlsf, tgw4pkh5equ6;

wire [56:0] egu8s6ddp42vmr_, y9y3ifqe7hc9;
wire [56:0] rdni7d46kfcdi42ua_u, en9y41nnuz2vzeawh, y7p07bro15sk6x, tmdz9eok35r5rqh372;
wire [56:0] b8yz7269cdmzraahb5fd, z6zj1f1qh0oelp37, ywljljk4a1d9jwh, k0irpzrxgjyru3yx4mp9k;

wire c2wxauj7al18yu52i = (~rg10e3avkel) & bpeajju419 & m0e2_guluq90ndzyt;
wire h_1o1ctw53rpnu = (~rg10e3avkel) & bpeajju419 & (~m0e2_guluq90ndzyt);
wire c6ljq5fny_e840w8 = (~c2wxauj7al18yu52i)&(~h_1o1ctw53rpnu);

wire [56:0] m12cj1uda_55q = {{57-53{1'b0}}, 1'b1, dsr2v_ycsx8gw} ;

wire [56:0] m2i1g5vbxt_66qc = rg10e3avkel ? rdni7d46kfcdi42ua_u : m12cj1uda_55q;

wire [56:0] xbafc6rtavt={57{c2wxauj7al18yu52i}}&{{57-52{1'b0}}, ohh5oui0c7_sw}
                           |{57{h_1o1ctw53rpnu }}&{{57-54{1'b0}}, ohh5oui0c7_sw[51], ~ohh5oui0c7_sw[51], ohh5oui0c7_sw[50:0], 1'b0} 
                           |{57{c6ljq5fny_e840w8 }}&b8yz7269cdmzraahb5fd;

wire [56:0] vikr4dkjqa  = {57{rg10e3avkel}} & en9y41nnuz2vzeawh ;
wire [56:0] rl03stxg_58y37 = {57{rg10e3avkel}} & z6zj1f1qh0oelp37 ;

ux607_gnrl_dffl #(57) sq7d6_w3q4d_( (bp_c30xz|rg10e3avkel), m2i1g5vbxt_66qc,f02vn4ah, gf33atgy, ru_wi) ;
ux607_gnrl_dffl #(57) zvtsw2kmy7cdj( (bp_c30xz|rg10e3avkel), vikr4dkjqa,gt_sq2dtwcr, gf33atgy, ru_wi) ;

ux607_gnrl_dffl #(57) doemfgbifhav91( (bp_c30xz|rg10e3avkel), xbafc6rtavt,qnj9dtloi3, gf33atgy, ru_wi) ;
ux607_gnrl_dffl #(57) cbip1swk1il6s( (bp_c30xz|rg10e3avkel), rl03stxg_58y37,vetlu9oe6w4uu, gf33atgy, ru_wi) ;


wire [56:0] mbdukyi7q31yfk ;
assign mbdukyi7q31yfk[56:0] = rg10e3avkel ? egu8s6ddp42vmr_[56:0] : {57{1'b0}} ;
ux607_gnrl_dffl #(57) d8gcnhha1qd( (bp_c30xz|rg10e3avkel), mbdukyi7q31yfk,j0xu7nslfaf, gf33atgy, ru_wi) ;

wire [56:0] ia0z1gm4t ;
assign ia0z1gm4t[56:0] = rg10e3avkel ? y9y3ifqe7hc9[56:0] : {2'b11, {56-1{1'b0}}} ;
ux607_gnrl_dffl #(57) bxifuvosuztpqot( (bp_c30xz|rg10e3avkel), ia0z1gm4t,hh9u1ei_, gf33atgy, ru_wi) ;


wire [56:0] frnl5v3o0_t7gza = {{57-54{1'b1}}, 1'b0, ~i4ia5732yw, 1'b1} ;
wire [56:0] xm8tp6rdhheq = {{57-54{1'b0}}, 1'b1, i4ia5732yw, 1'b0} ;

wire [56:0] r1n0w69_56r = frnl5v3o0_t7gza;
wire [56:0] jpsmvgay7 = xm8tp6rdhheq;

wire [56:0] zz7zrnav5  = rg10e3avkel ? {1'b0, y7p07bro15sk6x[(57-2):0]}  : {57{1'b0}} ; 
wire [56:0] hyfi70xcwvn = rg10e3avkel ? {1'b0, tmdz9eok35r5rqh372[(57-2):0]} : {57{1'b0}} ;

wire [56:0] qgb201ctaut  = rg10e3avkel ?  ywljljk4a1d9jwh  : {1'b1, {56{1'b0}}};
wire [56:0] kkszmj3b8q5hfov = rg10e3avkel ?  k0irpzrxgjyru3yx4mp9k : {57{1'b0}}      ;

wire [56:0] mt29_5butm72e = (rg10e3avkel ? (op5chmv5) : (mb75fcy6) )
                                ?  zz7zrnav5 :qgb201ctaut ;
wire [56:0] of1i8e_jw529exo =(rg10e3avkel ? (op5chmv5) : (mb75fcy6) )
                                ?  hyfi70xcwvn:kkszmj3b8q5hfov ;

wire [56:0] y0wrqy7l2h51920o898g ;
wire [56:0] whoml6jvz_49h7juvthtlt;

ux607_gnrl_dffl #(57) qwd66orrfap8jt_tkovsbnu( (bp_c30xz|rg10e3avkel), mt29_5butm72e,y0wrqy7l2h51920o898g, gf33atgy, ru_wi) ;
ux607_gnrl_dffl #(57) zftwu91_bzdepumvd7tjvghm0knn5( (bp_c30xz|rg10e3avkel), of1i8e_jw529exo,whoml6jvz_49h7juvthtlt, gf33atgy, ru_wi) ;

wire [56:0] l3sysfx =y0wrqy7l2h51920o898g;
wire [56:0] axhwk29y_ =whoml6jvz_49h7juvthtlt;

wire [56:0] bdl76yc6 =y0wrqy7l2h51920o898g;
wire [56:0] rpcdbj3xdniw =whoml6jvz_49h7juvthtlt;


wire [56:0] ojk8q0kqtxllaplj;
wire [56:0] b1pqez6o5omxzmfznu;

wire jdfz_dz2jhta5u1yf9gos;
wire n4jy7r9ysk_2d7ln1b ;
wire ltqug0zz86r6inrtrd3ka_;
wire [56:0] yr2h8vple3eqnb10komi;
wire [56:0] ga5vua0dxn26946fa8;

wire ryp5ontk__fndad_tb;
wire g6hanemcq58y1qbg9oq1 ;
wire s_71c29qisbvq8epzcgk;

wire [56:0] dj4yob34_3cd976v1j;
wire [56:0] z4a5yhlbtwxj9apjsyei;

wire g7cis5oe708ujt3x0cdwe;
wire hvel5rfcw7x9rm8cpg0fqk ;
wire p402yurs5fhwyc1_l05fyj;

wire [56:0] k8do2wvfeyicatk;
wire [56:0] rogttp_918epecp;
wire [56:0] dn_bzogydbhihkvzp ;
wire [56:0] x48yww8t6_;
wire [56:0] zzlnkkybj4u;

wire oyk2eu49b5f0eun1;
wire qx_3kns2zktoq89v ;
wire t6weyoe475iamw_a2s;

assign dn_bzogydbhihkvzp[56-1:0] = j0xu7nslfaf[56:1] ;
assign dn_bzogydbhihkvzp[56] = 1'b1 ;

assign x48yww8t6_  = (t6weyoe475iamw_a2s ? axhwk29y_ : l3sysfx) & dn_bzogydbhihkvzp | ~{57{qx_3kns2zktoq89v}} & ~dn_bzogydbhihkvzp ;
assign zzlnkkybj4u = (oyk2eu49b5f0eun1 ? l3sysfx : axhwk29y_) & dn_bzogydbhihkvzp | {57{qx_3kns2zktoq89v}} & ~dn_bzogydbhihkvzp ;

wire [56:0] lymqnwpqqd7eo     = k8do2wvfeyicatk;
wire [56:0] rem0ynapbt     = rogttp_918epecp;
wire [56:0] l7xy7kv51ktg8h13 = jpsmvgay7;
wire [56:0] rbi8qf9fn4a0egz = r1n0w69_56r;
wire [56:0] wdnl3il5muz    = dn_bzogydbhihkvzp;
wire [56:0] mab9c3nqmjs3     = x48yww8t6_;
wire [56:0] qpmqnbpmd_    = zzlnkkybj4u;

wire o50il7yxbt7z0x3d37 = (oyk2eu49b5f0eun1 & ryp5ontk__fndad_tb) | (t6weyoe475iamw_a2s & g7cis5oe708ujt3x0cdwe) | (qx_3kns2zktoq89v & jdfz_dz2jhta5u1yf9gos);
wire m635cj42noktlwru  = (oyk2eu49b5f0eun1 & g6hanemcq58y1qbg9oq1 ) | (t6weyoe475iamw_a2s & hvel5rfcw7x9rm8cpg0fqk ) | (qx_3kns2zktoq89v & n4jy7r9ysk_2d7ln1b );
wire alav2057kmm4ocdrj6p = (oyk2eu49b5f0eun1 & s_71c29qisbvq8epzcgk) | (t6weyoe475iamw_a2s & p402yurs5fhwyc1_l05fyj) | (qx_3kns2zktoq89v & ltqug0zz86r6inrtrd3ka_);

assign zbx4klyjkjk_39m[56-1:0] = wdnl3il5muz[56:1] ;
assign zbx4klyjkjk_39m[56] = 1'b1 ;

assign e9s410oe7si  = (alav2057kmm4ocdrj6p ? qpmqnbpmd_ : mab9c3nqmjs3) & zbx4klyjkjk_39m | ~{57{m635cj42noktlwru}} & ~zbx4klyjkjk_39m ;
assign ukt_9nlhm1d82lf = (o50il7yxbt7z0x3d37 ? mab9c3nqmjs3 : qpmqnbpmd_) & zbx4klyjkjk_39m | {57{m635cj42noktlwru}} & ~zbx4klyjkjk_39m ;

o_6c7gxntcc9ta0bisv_ m3aicq27z2xaq4zawr(
  .rydw         (f02vn4ah),
  .d4y         (gt_sq2dtwcr),
  .ust6kl      (oyk2eu49b5f0eun1),
  .p2yjv_h8o       (qx_3kns2zktoq89v ),
  .v2f5pmhic4      (t6weyoe475iamw_a2s)
);

k_f7ns0a54rui10fjf o8dihxfe89lavyttvyy(
  .f02vn4ah     (f02vn4ah),
  .gt_sq2dtwcr     (gt_sq2dtwcr),
  .lxff         (jpsmvgay7),
  .c2u         (r1n0w69_56r),
  .v2f5pmhic4      (t6weyoe475iamw_a2s),
  .ust6kl      (oyk2eu49b5f0eun1),
  .p2yjv_h8o       (qx_3kns2zktoq89v ),
  .xphx        (k8do2wvfeyicatk),
  .fap75        (rogttp_918epecp)
);

k_f7ns0a54rui10fjf de093bye1d40jtvon11ctzy0(
  .f02vn4ah     (f02vn4ah),
  .gt_sq2dtwcr     (gt_sq2dtwcr),
  .lxff         (jpsmvgay7),
  .c2u         (r1n0w69_56r),
  .v2f5pmhic4      (1'b0),
  .ust6kl      (1'b0),
  .p2yjv_h8o       (1'b1 ),
  .xphx    (ojk8q0kqtxllaplj),
  .fap75    (b1pqez6o5omxzmfznu)
);

o_6c7gxntcc9ta0bisv_ av5_ksyzfr_kxe8hh_qhos20h(
  .rydw     (ojk8q0kqtxllaplj),
  .d4y     (b1pqez6o5omxzmfznu),
  .ust6kl  (jdfz_dz2jhta5u1yf9gos),
  .p2yjv_h8o   (n4jy7r9ysk_2d7ln1b ),
  .v2f5pmhic4  (ltqug0zz86r6inrtrd3ka_)
);

k_f7ns0a54rui10fjf bvgqo389l506i5xifmx8p(
  .f02vn4ah  (f02vn4ah),
  .gt_sq2dtwcr  (gt_sq2dtwcr),
  .lxff      (jpsmvgay7),
  .c2u      (r1n0w69_56r),
  .v2f5pmhic4   (1'b0),
  .ust6kl   (1'b1),
  .p2yjv_h8o    (1'b0 ),
  .xphx     (yr2h8vple3eqnb10komi),
  .fap75     (ga5vua0dxn26946fa8)
);

o_6c7gxntcc9ta0bisv_ i7cl0g27ah_cth33swo469k94m5(
  .rydw     (yr2h8vple3eqnb10komi),
  .d4y     (ga5vua0dxn26946fa8),
  .ust6kl  (ryp5ontk__fndad_tb),
  .p2yjv_h8o   (g6hanemcq58y1qbg9oq1 ),
  .v2f5pmhic4  (s_71c29qisbvq8epzcgk)
);

k_f7ns0a54rui10fjf xm513tsl9asq0udbyda2c4x1(
  .f02vn4ah     (f02vn4ah),
  .gt_sq2dtwcr     (gt_sq2dtwcr),
  .lxff         (jpsmvgay7),
  .c2u         (r1n0w69_56r),
  .v2f5pmhic4      (1'b1),
  .ust6kl      (1'b0),
  .p2yjv_h8o       (1'b0 ),
  .xphx        (dj4yob34_3cd976v1j),
  .fap75        (z4a5yhlbtwxj9apjsyei)
);

o_6c7gxntcc9ta0bisv_ hxfjldgp8743mrsohpen0165g(
  .rydw     (dj4yob34_3cd976v1j),
  .d4y     (z4a5yhlbtwxj9apjsyei),
  .ust6kl  (g7cis5oe708ujt3x0cdwe),
  .p2yjv_h8o   (hvel5rfcw7x9rm8cpg0fqk ),
  .v2f5pmhic4  (p402yurs5fhwyc1_l05fyj)
);

k_f7ns0a54rui10fjf i5oohtdnevwj10_yw5d1b(
  .f02vn4ah    (lymqnwpqqd7eo),
  .gt_sq2dtwcr    (rem0ynapbt),
  .lxff        (l7xy7kv51ktg8h13),
  .c2u        (rbi8qf9fn4a0egz),
  .v2f5pmhic4     (alav2057kmm4ocdrj6p),
  .ust6kl     (o50il7yxbt7z0x3d37),
  .p2yjv_h8o      (m635cj42noktlwru ),
  .xphx       (kpgls4tvuy_dq9a),
  .fap75       (xa5onwxrrff4hh)
);

wire [56:0]  ttvgztn4ru160b   ;
wire [56:0]  oh1pxv8qcnplrgo3   ;
wire [56:0]  lovw9bfiau5   ;
wire [56:0]  mxitknpihbhrw5sww  ;
wire [56:0] gi76ah3kj_olhbn78 ;
wire [56:0] boaiq6wchz7i2 ;

wire bxnmrvfiby6xnqw;
wire a6kr5mct028pmi0y ;
wire g0vipqrmixsjij2hpqh;

wire [56:0] sgi9gzhjru8d892uvzal;
wire [56:0] zg60fn4x_hifd3tzr99ws5;
wire fach7g602cp5pfv495hxfsi2;
wire sttd9ltzewe96u0avin ;
wire tj3_m_2dk6y0ne3vsh3ny7h;

wire [56:0] dapzhiwux43bk048sk2eu;
wire [56:0] jk3enwxs2jgr01wut8k93c;

wire [56:0]  czepceb8cf30t  = ttvgztn4ru160b;
wire [56:0]  iemo64unuz  = oh1pxv8qcnplrgo3;
wire [56:0]  f9i_bkopj9l = gi76ah3kj_olhbn78;
wire [56:0]  ajtqi23mcudo = boaiq6wchz7i2;
wire [56:0]  jktrsmt_35  = lovw9bfiau5 ;
wire [56:0]  m90slbblo4kr = mxitknpihbhrw5sww;
wire x7vywfbj3dtfvtk9_u2ac_;
wire q18e0mz7vc6mig449yc3qqq ;
wire ak2yhshn8shq149lie4lvhbr;
wire [56:0] oyav5pb1eqa80315m9hson;
wire [56:0] ov_aksk53u0_umg1g;
wire dlk4u_9nr9jwdqouudg;
wire kk06y2e5djq5d3dqqga_ ;
wire xixvcz37its5hkaykvc;

assign gi76ah3kj_olhbn78[56-1:0] = j0xu7nslfaf[56:1] ;
assign gi76ah3kj_olhbn78[56] = 1'b1 ;

assign boaiq6wchz7i2[56-1:0] = hh9u1ei_[56:1] ;
assign boaiq6wchz7i2[56] = 1'b0 ;

assign lovw9bfiau5  = (g0vipqrmixsjij2hpqh ? rpcdbj3xdniw : bdl76yc6) & gi76ah3kj_olhbn78 | ~{57{a6kr5mct028pmi0y}} & ~gi76ah3kj_olhbn78 ;
assign mxitknpihbhrw5sww = (bxnmrvfiby6xnqw ? bdl76yc6 : rpcdbj3xdniw) & gi76ah3kj_olhbn78 | {57{a6kr5mct028pmi0y}} & ~gi76ah3kj_olhbn78 ;

wire z0nhfvlkven7d46k148 = (bxnmrvfiby6xnqw & dlk4u_9nr9jwdqouudg) | (g0vipqrmixsjij2hpqh & x7vywfbj3dtfvtk9_u2ac_) | (a6kr5mct028pmi0y & fach7g602cp5pfv495hxfsi2);
wire peilpz_ztgggjru81rx  = (bxnmrvfiby6xnqw & kk06y2e5djq5d3dqqga_ ) | (g0vipqrmixsjij2hpqh & q18e0mz7vc6mig449yc3qqq ) | (a6kr5mct028pmi0y & sttd9ltzewe96u0avin );
wire et0yen5jfo2lf2pc8ob = (bxnmrvfiby6xnqw & xixvcz37its5hkaykvc) | (g0vipqrmixsjij2hpqh & ak2yhshn8shq149lie4lvhbr) | (a6kr5mct028pmi0y & tj3_m_2dk6y0ne3vsh3ny7h);

assign auu79qzp63t0_cc0ru[56-1:0] = f9i_bkopj9l[56:1] ;
assign auu79qzp63t0_cc0ru[56] = 1'b1 ;

assign qng6_z6rdlwu3[56-1:0] = ajtqi23mcudo[56:1] ;
assign qng6_z6rdlwu3[56] = 1'b0 ;

assign nm2k_djs2vlsf  = (et0yen5jfo2lf2pc8ob ? m90slbblo4kr : jktrsmt_35) & auu79qzp63t0_cc0ru | ~{57{peilpz_ztgggjru81rx}} & ~auu79qzp63t0_cc0ru ;
assign tgw4pkh5equ6 = (z0nhfvlkven7d46k148 ? jktrsmt_35 : m90slbblo4kr) & auu79qzp63t0_cc0ru | {57{peilpz_ztgggjru81rx}} & ~auu79qzp63t0_cc0ru ;


o_6c7gxntcc9ta0bisv_ rc1u9jfq92zxwewd983(
  .rydw     (qnj9dtloi3),
  .d4y     (vetlu9oe6w4uu),
  .ust6kl(bxnmrvfiby6xnqw),
  .p2yjv_h8o (a6kr5mct028pmi0y ),
  .v2f5pmhic4(g0vipqrmixsjij2hpqh)
);

j3rmuwv9gah_ceeqolq8gh hcrebfd_hlyywllt8_fgxo(
  .j0xu7nslfaf  (gi76ah3kj_olhbn78  ),
  .hh9u1ei_  (boaiq6wchz7i2  ),
  .qnj9dtloi3     (qnj9dtloi3     ),
  .vetlu9oe6w4uu     (vetlu9oe6w4uu     ),
  .bdl76yc6     (bdl76yc6     ),
  .rpcdbj3xdniw    (rpcdbj3xdniw    ),
  .ust6kl(bxnmrvfiby6xnqw),
  .p2yjv_h8o (a6kr5mct028pmi0y ),
  .v2f5pmhic4(g0vipqrmixsjij2hpqh),
  .xphx    (ttvgztn4ru160b    ),
  .fap75    (oh1pxv8qcnplrgo3    )
);

j3rmuwv9gah_ceeqolq8gh he0ghe1fxooarbft880d2s_i(
  .j0xu7nslfaf  (gi76ah3kj_olhbn78  ),
  .hh9u1ei_  (boaiq6wchz7i2  ),
  .qnj9dtloi3     (qnj9dtloi3     ),
  .vetlu9oe6w4uu     (vetlu9oe6w4uu     ),
  .bdl76yc6     (bdl76yc6     ),
  .rpcdbj3xdniw    (rpcdbj3xdniw    ),
  .ust6kl(1'b0),
  .p2yjv_h8o (1'b1 ),
  .v2f5pmhic4(1'b0),
  .xphx    (sgi9gzhjru8d892uvzal    ),
  .fap75    (zg60fn4x_hifd3tzr99ws5    )
);

o_6c7gxntcc9ta0bisv_ kszarpk0ok6lgvq8n8ghcg3iooa(
  .rydw     (sgi9gzhjru8d892uvzal),
  .d4y     (zg60fn4x_hifd3tzr99ws5),
  .ust6kl(fach7g602cp5pfv495hxfsi2),
  .p2yjv_h8o (sttd9ltzewe96u0avin ),
  .v2f5pmhic4(tj3_m_2dk6y0ne3vsh3ny7h)
);

j3rmuwv9gah_ceeqolq8gh xsgsyy_qrazvmjprmqubxpoq7(
  .j0xu7nslfaf  (gi76ah3kj_olhbn78  ),
  .hh9u1ei_  (boaiq6wchz7i2  ),
  .qnj9dtloi3     (qnj9dtloi3     ),
  .vetlu9oe6w4uu     (vetlu9oe6w4uu     ),
  .bdl76yc6     (bdl76yc6     ),
  .rpcdbj3xdniw    (rpcdbj3xdniw    ),
  .ust6kl(1'b0),
  .p2yjv_h8o (1'b0 ),
  .v2f5pmhic4(1'b1),
  .xphx    (dapzhiwux43bk048sk2eu    ),
  .fap75    (jk3enwxs2jgr01wut8k93c    )
);

o_6c7gxntcc9ta0bisv_ pif2tnv84k6n7h42umga_r0yoo(
  .rydw     (dapzhiwux43bk048sk2eu),
  .d4y     (jk3enwxs2jgr01wut8k93c),
  .ust6kl(x7vywfbj3dtfvtk9_u2ac_),
  .p2yjv_h8o (q18e0mz7vc6mig449yc3qqq ),
  .v2f5pmhic4(ak2yhshn8shq149lie4lvhbr)
);

j3rmuwv9gah_ceeqolq8gh s_0se4um3s8lbue1099m17x4o5e(
  .j0xu7nslfaf  (gi76ah3kj_olhbn78  ),
  .hh9u1ei_  (boaiq6wchz7i2  ),
  .qnj9dtloi3     (qnj9dtloi3     ),
  .vetlu9oe6w4uu     (vetlu9oe6w4uu     ),
  .bdl76yc6     (bdl76yc6     ),
  .rpcdbj3xdniw    (rpcdbj3xdniw    ),
  .ust6kl(1'b1),
  .p2yjv_h8o (1'b0 ),
  .v2f5pmhic4(1'b0),
  .xphx    (oyav5pb1eqa80315m9hson    ),
  .fap75    (ov_aksk53u0_umg1g    )
);

o_6c7gxntcc9ta0bisv_ olq050kk4rmedzqu38cflesnar(
  .rydw     (oyav5pb1eqa80315m9hson),
  .d4y     (ov_aksk53u0_umg1g),
  .ust6kl(dlk4u_9nr9jwdqouudg),
  .p2yjv_h8o (kk06y2e5djq5d3dqqga_ ),
  .v2f5pmhic4(xixvcz37its5hkaykvc)
);

j3rmuwv9gah_ceeqolq8gh gzo6r385p3vaf5jkvqkb0n(
  .j0xu7nslfaf  (auu79qzp63t0_cc0ru  ),
  .hh9u1ei_  (qng6_z6rdlwu3  ),
  .qnj9dtloi3     (czepceb8cf30t     ),
  .vetlu9oe6w4uu     (iemo64unuz     ),
  .bdl76yc6     (jktrsmt_35     ),
  .rpcdbj3xdniw    (m90slbblo4kr    ),
  .ust6kl(z0nhfvlkven7d46k148),
  .p2yjv_h8o (peilpz_ztgggjru81rx ),
  .v2f5pmhic4(et0yen5jfo2lf2pc8ob),
  .xphx    (cwpbbg1e2nj0_4    ),
  .fap75    (akr00lq3hfph    )
);



wire [56:0] hwqvqv2vg878jbynag4ryrcx  = y0wrqy7l2h51920o898g;
wire [56:0] kn9671jc047ux3q9yah    = f02vn4ah;
wire [56:0] rar8x5t9fi4syd7i6uyk5s    = gt_sq2dtwcr;
wire [56:0] nrywq2tmp3g982cvvginuc7   = qnj9dtloi3;
wire [56:0] e8tzezf_thfz1km4te5u6fyx   = vetlu9oe6w4uu;
wire [56:0] kj26lnz73c8d__9na = (op5chmv5)? kn9671jc047ux3q9yah : nrywq2tmp3g982cvvginuc7;
wire [56:0] dlvkaeviq1zaag674rqh = (op5chmv5)? rar8x5t9fi4syd7i6uyk5s : e8tzezf_thfz1km4te5u6fyx;

assign y7p07bro15sk6x = e9s410oe7si ;
assign tmdz9eok35r5rqh372 = ukt_9nlhm1d82lf ;
assign ywljljk4a1d9jwh = nm2k_djs2vlsf ;
assign k0irpzrxgjyru3yx4mp9k = tgw4pkh5equ6 ;
assign rdni7d46kfcdi42ua_u =  kpgls4tvuy_dq9a ;
assign en9y41nnuz2vzeawh =  xa5onwxrrff4hh ;
assign b8yz7269cdmzraahb5fd = cwpbbg1e2nj0_4 ;
assign z6zj1f1qh0oelp37 = akr00lq3hfph ;
assign egu8s6ddp42vmr_ =    zbx4klyjkjk_39m ;
assign y9y3ifqe7hc9 =    qng6_z6rdlwu3;

wire dxxo5mff9x_pbcd;
wire [56:0] fi4wkjfu_s;
wire [56:0] lvp4vbfx0yanj2bx;
wire [56:0] jlegg9zaqp;

wire o2hwq7m3;
wire tpe8tof60d;
wire m0qhdqaf5;
wire g3p10kiz99y850a;
wire iapkhff31e8bvi;
wire x6zbixrb07sg20;
wire mvmgfmewg0eh3;
wire kwwz987lpvix_s;

wire [12:0] rs_sll4oetbhrkvo;
wire [12:0] huh3ueqh1jxsvjurg;
wire [12:0] to1yx1mxgbw;
wire [5:0] fyhrv__1qga;
wire pg6vffbz3lj1aqrks;
wire xmlpt3as21gtcu65s;

wire [56:0] fslbafh5 = kj26lnz73c8d__9na + dlvkaeviq1zaag674rqh ;
wire [56:0] rgl7v53v9fe4w = nv_meva_f5 ? {3'b000, hwqvqv2vg878jbynag4ryrcx[56:9], 6'b10_0000} : 
                         {3'b000, hwqvqv2vg878jbynag4ryrcx[56:29],4'b0001,22'b0} ;

wire [56:0] im5xxv64qn9u = xm8tp6rdhheq;
wire j3gwgnl_ = fslbafh5[56] ;

wire [56:0] h2e8eht6 = (op5chmv5)? im5xxv64qn9u : rgl7v53v9fe4w;

wire [56:0] nmmz7gswmabdihxn5p  = y0wrqy7l2h51920o898g ;
wire [56:0] po8w3w8z5tnix96ro__n = whoml6jvz_49h7juvthtlt;

wire [56:0] hx5felzbbf = j3gwgnl_ ? po8w3w8z5tnix96ro__n : nmmz7gswmabdihxn5p;

wire [56:0] fded423k;
wire [56:0] h0js8u6p55qu8=bp_c30xz ? 1'b1 : fslbafh5;
assign yh0oeg399pvwaqg13 = (op5chmv5)&(fded423k== {57{1'b0}});

wire [56:0] zsz1wphlt0 = fi4wkjfu_s + lvp4vbfx0yanj2bx;
wire [56:0] afouypklip6  = dxxo5mff9x_pbcd ? zsz1wphlt0 : fi4wkjfu_s ;
wire xpm13cra8w0y         = (afouypklip6== {57{1'b0}});
wire ox3y1gv0vfar4iq        = jlegg9zaqp[56-1] ;
wire sx0shfi3_8zl_pm   = ~ox3y1gv0vfar4iq;
wire rtbvl1ryh8fm2vb0rqc4   = jlegg9zaqp[56] ;


ux607_gnrl_dffl #(57) if1deobm68ju92r( (bp_c30xz|rg10e3avkel), h0js8u6p55qu8,fded423k, gf33atgy, ru_wi);
ux607_gnrl_dffl #(1) i9esawrbkjmokzsz4pw0( bhmxsiib6, j3gwgnl_,dxxo5mff9x_pbcd, gf33atgy, ru_wi);
ux607_gnrl_dffl #(57) l_ljh9nufqq95ylai( bhmxsiib6, fslbafh5,fi4wkjfu_s, gf33atgy, ru_wi);
ux607_gnrl_dffl #(57) st32ct72pogmwjs8j1z( bhmxsiib6, h2e8eht6,lvp4vbfx0yanj2bx, gf33atgy, ru_wi);
ux607_gnrl_dffl #(57) pbl8x5w_9aws( bhmxsiib6, hx5felzbbf,jlegg9zaqp, gf33atgy, ru_wi);
ux607_gnrl_dffl #(1) r4q3o1q490tsgv4x5i( bhmxsiib6, op5chmv5&o2hwq7m3,g3p10kiz99y850a, gf33atgy, ru_wi);
ux607_gnrl_dffl #(1) ly61_zjiqmu9myn9iw( bhmxsiib6, op5chmv5&tpe8tof60d,iapkhff31e8bvi, gf33atgy, ru_wi);
ux607_gnrl_dffl #(1) t06uyncot37pleip27ky13( bhmxsiib6, op5chmv5&m0qhdqaf5,x6zbixrb07sg20, gf33atgy, ru_wi);
ux607_gnrl_dffl #(1) gbfyu85ks4i53bvfeveu4i( vawmftolubc5, g3p10kiz99y850a,mvmgfmewg0eh3, gf33atgy, ru_wi);
ux607_gnrl_dffl #(1) ysbwrd1w3oq87797ewk5( vawmftolubc5, x6zbixrb07sg20,kwwz987lpvix_s, gf33atgy, ru_wi);
ux607_gnrl_dffl #(13) wyfp9lassfzaip_5d4lc( bhmxsiib6, rs_sll4oetbhrkvo,huh3ueqh1jxsvjurg, gf33atgy, ru_wi);
ux607_gnrl_dffl #(6) dnv88j3b7vopxtn( bhmxsiib6, to1yx1mxgbw[5:0],fyhrv__1qga, gf33atgy, ru_wi);
ux607_gnrl_dffl #(1) tmxocrvc5g373iuso7_wu( bhmxsiib6, pg6vffbz3lj1aqrks,xmlpt3as21gtcu65s, gf33atgy, ru_wi);

w8pxut7bux607aof8nd6je #(.onr7l(13)) h7urdk3t58yxu9hbvef(
  .gf33atgy        (gf33atgy),
  .ru_wi    (ru_wi),
  .bp_c30xz (bp_c30xz),
  .ii         ({2'b0,cs118t0ggohu0}),
  .fij51v         (~{2'b0,yruj_3_m8kmx8}),
  .cuzhl9         (q02bklc ? 13'h3FF:13'h7F),
  .oho1e63         ({7'b0,dvmjxjsqko9mdgn}),
  .hl69c         (~{7'b0,a0_2x3l9euvn1ixa6}),
  .mck7r06         (13'd2),
  .tsa1sag7   (rs_sll4oetbhrkvo)
);

w8pxut7bux607aof8nd6je #(.onr7l(13)) vm_zoh5001c70uk2uds(
  .gf33atgy        (gf33atgy),
  .ru_wi    (ru_wi),
  .bp_c30xz (bp_c30xz),
  .ii         (~{2'b0,cs118t0ggohu0}),
  .fij51v         ({2'b0,yruj_3_m8kmx8}),
  .cuzhl9         (~(q02bklc ? 13'h3FF:13'h7F)),
  .oho1e63         (~{7'b0,dvmjxjsqko9mdgn}),
  .hl69c         ({7'b0,a0_2x3l9euvn1ixa6}),
  .mck7r06         (13'd4),
  .tsa1sag7   (to1yx1mxgbw)
);


wire f6dc_rhcaz;
wire [11:0] f85ls0c84jdusxpj0fqqbr1175;
wire [11:0] qwk89od3zqk9ocn6hw6rm42xjc;

wire   aw8h6wznps9fw_d9cm5a7v = rs_sll4oetbhrkvo[12];                     
wire   s8q0bcqtftp3 = (rs_sll4oetbhrkvo == 13'b0);

wire y95w4pry23vsxc33_ex = (to1yx1mxgbw[5:1]>28) & aw8h6wznps9fw_d9cm5a7v;
wire gz30tebme8k22oo53bm5x = (to1yx1mxgbw[5:1]>14) & aw8h6wznps9fw_d9cm5a7v;

wire[4:0] ugixkk95fnte94g= (~op5chmv5) ? 5'd14  
          : (~gz30tebme8k22oo53bm5x) ? (5'd14 + (~({5{aw8h6wznps9fw_d9cm5a7v}} & to1yx1mxgbw[5:1])) + 1'b1)
          : 5'd0;

wire[4:0] iqn0_owvr06= (~op5chmv5) ? 5'd28 
          : (~y95w4pry23vsxc33_ex) ? (5'd28 + (~({5{aw8h6wznps9fw_d9cm5a7v}} & to1yx1mxgbw[5:1])) + 1'b1)
          : 5'd0;

wire [11:0] rvah9en2chetm8w6mf = {1'b0,a4meogg6iciznynf} + {{5{rvezutl8owb63ik2aznm[6]}},rvezutl8owb63ik2aznm};

assign gd2wkhivb2 = nv_meva_f5 ?  iqn0_owvr06 : ugixkk95fnte94g;
assign tpe8tof60d = (rs_sll4oetbhrkvo == 13'b1);
assign m0qhdqaf5 = (~s8q0bcqtftp3) & (~tpe8tof60d) & (~aw8h6wznps9fw_d9cm5a7v);
assign o2hwq7m3 = (s8q0bcqtftp3 | aw8h6wznps9fw_d9cm5a7v);
assign pg6vffbz3lj1aqrks = (to1yx1mxgbw>53) & aw8h6wznps9fw_d9cm5a7v;



wire [56:0] vsmguz1__im81kqzn9y;
wire [56:0] yeazfbb8egum7gjtt3zl9fh;
wire [12:0] jr3tmmwtj06wdrg;
wire [52:0] p9qeu2pjdxh;
wire [3:0] bk7x5cj2zoyv9t;
wire h7x1e7166csgyh1;
wire [56:0] qwwfo8xgne6nu71t45n7n;
wire [52:0] gdowa, apc943j7j, sqtqelcz862j78;
wire h8vwv1, fll_n3vj832wn, km84pb15bchx0g7;

assign {vsmguz1__im81kqzn9y,yeazfbb8egum7gjtt3zl9fh} = {jlegg9zaqp,{(56+1){1'b0}}}>>fyhrv__1qga;


wire [56:0] r0u1kyleu = ({57{g3p10kiz99y850a}} & (xmlpt3as21gtcu65s ? {57{1'b0}} : vsmguz1__im81kqzn9y))
                     | ({57{iapkhff31e8bvi}} & jlegg9zaqp)
                     | ({57{x6zbixrb07sg20}} & (ox3y1gv0vfar4iq ? {jlegg9zaqp[56:0]} : {jlegg9zaqp[56-1:0],1'b0}));

wire [12:0] fpqy39n3k8abm = ({13{g3p10kiz99y850a}} & (13'd1))
                        | ({13{iapkhff31e8bvi}} & huh3ueqh1jxsvjurg)
                        | ({13{x6zbixrb07sg20}} & (huh3ueqh1jxsvjurg + {13{sx0shfi3_8zl_pm}}));

wire [56:0] xk23eae8gc91n9ec = xmlpt3as21gtcu65s ? jlegg9zaqp : yeazfbb8egum7gjtt3zl9fh; 
wire wglm82x5c1mnfcp_q6hkb82  = mvmgfmewg0eh3 & (|qwwfo8xgne6nu71t45n7n);

wire [52:0] zebs5mq2l = rtbvl1ryh8fm2vb0rqc4 ? {jlegg9zaqp[56:56-52]} : {jlegg9zaqp[56-1:56-53]} ;
wire [3:0] vhnbq98y2hnl2zzus = rtbvl1ryh8fm2vb0rqc4 ? {jlegg9zaqp[56-52-1:0]} : {jlegg9zaqp[56-53-1:0],1'b0} ;

wire [52:0] a8uv18 = (jdnbsmmk7_x9) ? r0u1kyleu[56-1:56-53] : zebs5mq2l ;
wire [3:0] a309pces6p0p = (jdnbsmmk7_x9) ? {r0u1kyleu[56-53-1:0],1'b0} : vhnbq98y2hnl2zzus ;


ux607_gnrl_dffl #(12)rdp3qnfwm9721uyw1lw_07o6kts2xid( bhmxsiib6, rvah9en2chetm8w6mf,f85ls0c84jdusxpj0fqqbr1175,          gf33atgy, ru_wi);
ux607_gnrl_dffl #(12)r3rt7z7iodwa5a0tg6qwamcnece( vawmftolubc5, f85ls0c84jdusxpj0fqqbr1175,qwk89od3zqk9ocn6hw6rm42xjc, gf33atgy, ru_wi);
ux607_gnrl_dffl #(13) p8oyg77jkojke9n7i7ucic( vawmftolubc5, fpqy39n3k8abm,jr3tmmwtj06wdrg, gf33atgy, ru_wi);
ux607_gnrl_dffl #(57) aqzjs8syb55azjciefg_u8ah( vawmftolubc5, xk23eae8gc91n9ec,qwwfo8xgne6nu71t45n7n, gf33atgy, ru_wi);
ux607_gnrl_dffl #(53) zvyi3kxip8i3lw( vawmftolubc5, a8uv18,p9qeu2pjdxh, gf33atgy, ru_wi) ;
ux607_gnrl_dffl #(4) ktjb31i_3cipvl_cpjk( vawmftolubc5, a309pces6p0p,bk7x5cj2zoyv9t, gf33atgy, ru_wi) ;
ux607_gnrl_dffl #(1) a85nlh1iwwst4li4xz9q( vawmftolubc5, xpm13cra8w0y,h7x1e7166csgyh1, gf33atgy, ru_wi) ;

wire c8u66cjxyns73yg = p9qeu2pjdxh[0];
wire ho3nmrzws6vtaemz8p = bk7x5cj2zoyv9t[3];
wire l00yueru68d12d4f2 = bk7x5cj2zoyv9t[2];
wire g07b4c8ge45w3atcf = (|bk7x5cj2zoyv9t[1:0]) | (~h7x1e7166csgyh1);

wire t6sznn5l0ldwir_ztjy = p9qeu2pjdxh[29] ;                       
wire b8ghkgch59xnntr8jmel = p9qeu2pjdxh[28] ;                       
wire jy2uvfc7go8xx_q76v = p9qeu2pjdxh[27] ;                       
wire a89wuxey1pwezizw7 = p9qeu2pjdxh[26] | (~h7x1e7166csgyh1);

wire njbfrll57hduz0gcbsz = p9qeu2pjdxh[0] ;
wire yzbrdedseueb6r = bk7x5cj2zoyv9t[3] ;
wire kz8kqw9evz55kpey6 = bk7x5cj2zoyv9t[2] ;
wire fciacunit76jsppip = (|bk7x5cj2zoyv9t[1:0]) | (~h7x1e7166csgyh1);
                                                                             
wire dsxw4njkuwpmci97bw = p9qeu2pjdxh[29] ;                       
wire chv6pqxt9jgtcvubm = p9qeu2pjdxh[28] ;                       
wire ab9xmsvp3lk8k3l = p9qeu2pjdxh[27] ;                       
wire swo1071z6suyo5wv = p9qeu2pjdxh[26] | (~h7x1e7166csgyh1) ;

wire cj608wi42e = ka66jgi ? njbfrll57hduz0gcbsz : c8u66cjxyns73yg ;
wire vnivl57c9sfut = ka66jgi ? yzbrdedseueb6r : ho3nmrzws6vtaemz8p ;
wire pcd9vwjlol = ka66jgi ? kz8kqw9evz55kpey6 : l00yueru68d12d4f2 ;
wire gi4fsbataoo = ka66jgi ? fciacunit76jsppip : g07b4c8ge45w3atcf ;

wire q9l1j1xjo9s200 = ka66jgi ? dsxw4njkuwpmci97bw : t6sznn5l0ldwir_ztjy ;
wire xuysysmjpoddo = ka66jgi ? chv6pqxt9jgtcvubm : b8ghkgch59xnntr8jmel ;
wire xnlli6ptlmwd = ka66jgi ? ab9xmsvp3lk8k3l : jy2uvfc7go8xx_q76v ;
wire x7cvs2r3etdiv1 = ka66jgi ? swo1071z6suyo5wv : a89wuxey1pwezizw7 ;

wire p8j7vc63dn8v = y_zx8qolynd ? cj608wi42e : q9l1j1xjo9s200; 
wire o8eq0fhbx_h = y_zx8qolynd ? vnivl57c9sfut : xuysysmjpoddo; 
wire sm8nhlw = y_zx8qolynd ? pcd9vwjlol : xnlli6ptlmwd; 

wire aebb51i = (y_zx8qolynd ? gi4fsbataoo : x7cvs2r3etdiv1) 
                    | (ka66jgi &
                        (wglm82x5c1mnfcp_q6hkb82 | 
                        ((~y_zx8qolynd) & mvmgfmewg0eh3 & (|{p9qeu2pjdxh[26-1:0],
                        bk7x5cj2zoyv9t[3]})))); 

el7n_zz16sk_ntvue9v fg2z6emqrpgfdyuxg (   
	            .l     (p8j7vc63dn8v),          
                .g     (o8eq0fhbx_h),        
                .r     (sm8nhlw),        
                .s     (aebb51i),             
                .ly53de  (fvz__7_m),        
                .nfj6b    (ljxpmbsqoaz),    
                .f6dc_rhcaz(f6dc_rhcaz) );

assign {km84pb15bchx0g7, sqtqelcz862j78} = y_zx8qolynd ? ({1'b0, p9qeu2pjdxh} + 1'b1) : ({1'b0, p9qeu2pjdxh[52:29], 29'b0} + {1'b0,23'b0, 1'b1, 29'b0});
assign {fll_n3vj832wn, apc943j7j} = y_zx8qolynd ? {1'b0,p9qeu2pjdxh} : {1'b0, p9qeu2pjdxh[52:29], 29'b0} ;
assign gdowa  = f6dc_rhcaz ? sqtqelcz862j78 : apc943j7j;
assign h8vwv1 = f6dc_rhcaz ? km84pb15bchx0g7 : fll_n3vj832wn;

wire [63:0] et2w664wl8r ;
wire [31:0] v12nwpm6b862ua ;
wire i2a4sa38;

assign et2w664wl8r[63] = fvz__7_m;
assign v12nwpm6b862ua[31] = fvz__7_m;

wire oh15w5jmoca3r5;
wire ttrnyu5c0pc5;
wire [11:0] b4mdgpn31fgjrul_1p;
wire [12:0] mht1y4n6zc2aajj;
wire [9:0] uopbiut50sdz;
assign et2w664wl8r[62:52] = ka66jgi ? ({11{~oh15w5jmoca3r5}} & mht1y4n6zc2aajj[10:0]) : { b4mdgpn31fgjrul_1p[11:1]} ;
assign v12nwpm6b862ua[30:23] = ka66jgi ? ({8{~ttrnyu5c0pc5}}  & uopbiut50sdz[7:0]) : { b4mdgpn31fgjrul_1p[8:1]} ;

assign et2w664wl8r[51:0] = ((~kwwz987lpvix_s) | gdowa[52] | h8vwv1) ? {gdowa[51:0]} : {gdowa[50:0], p8j7vc63dn8v} ;
assign v12nwpm6b862ua[22:0] = ((~kwwz987lpvix_s) | gdowa[52] | h8vwv1) ? gdowa[51:29] : gdowa[50:28] ;
wire si234d0f = ((((~kwwz987lpvix_s) | gdowa[52]) ? gdowa[52] : gdowa[51])|h8vwv1);
wire dvouzr = ((((~kwwz987lpvix_s) | gdowa[52]) ? gdowa[52] : gdowa[51])|h8vwv1);
wire sm3rrrhja_p6d6utl7e = (((~kwwz987lpvix_s) | apc943j7j[52]) ? apc943j7j[52] : apc943j7j[51]) ;
wire i7k31a_zvsq9nstij = (((~kwwz987lpvix_s) | apc943j7j[52]) ? apc943j7j[52] : apc943j7j[51]) ;

assign uopbiut50sdz = jr3tmmwtj06wdrg[09:0];
assign mht1y4n6zc2aajj = jr3tmmwtj06wdrg[12:0];

wire [09:0] matiyswm3pmubak_r022adjn = jr3tmmwtj06wdrg[09:0];
wire [12:0] tgkw76xftrgb1f91du6 = jr3tmmwtj06wdrg[12:0];

assign b4mdgpn31fgjrul_1p = h8vwv1 ? (qwk89od3zqk9ocn6hw6rm42xjc + 1'b1 +(y_zx8qolynd ? 12'd1023:12'd127))
                              :(qwk89od3zqk9ocn6hw6rm42xjc +(y_zx8qolynd ? 12'd1023:12'd127));

wire flauo_jzxcn = ((|mht1y4n6zc2aajj[12:11]) | (mht1y4n6zc2aajj==2047));
wire zonduy8o72hw8f = ((|uopbiut50sdz[9:8]) | (uopbiut50sdz==255));

wire ox2rkt49cl = flauo_jzxcn & ka66jgi ;
wire ibzugz1v = zonduy8o72hw8f & ka66jgi ;

wire xwk7fm0 = y_zx8qolynd ? ox2rkt49cl : ibzugz1v ;

assign oh15w5jmoca3r5 = (mht1y4n6zc2aajj==13'b1)&(~si234d0f)&ka66jgi;
assign ttrnyu5c0pc5 = (uopbiut50sdz==10'b1)&(~dvouzr)&ka66jgi;

wire p9bg8yc6 = (tgkw76xftrgb1f91du6==13'b1)&(~sm3rrrhja_p6d6utl7e)&ka66jgi;
wire dlwqm1 = (matiyswm3pmubak_r022adjn==10'b1)&(~i7k31a_zvsq9nstij)&ka66jgi;

assign i2a4sa38 = ((o8eq0fhbx_h | sm8nhlw | aebb51i) & (y_zx8qolynd ? p9bg8yc6 : dlwqm1 ));

wire a_xtsojke05dnao = 1'b0; 
wire gp5nsjv6nris3nx7zm2 = 1'b0; 
wire ixn122itx74ljf0e8dk = y_zx8qolynd ? ox2rkt49cl : ibzugz1v ;
wire fipd_e_m294cc01e54bb = i2a4sa38 ;
wire wb3pal8jhelc__t0 = ((o8eq0fhbx_h | sm8nhlw | aebb51i | ixn122itx74ljf0e8dk)) ;


wire bn60jfu_ewb = 
             ( (xwk7fm0 & (ljxpmbsqoaz == 3'b100))
             | (xwk7fm0 & (ljxpmbsqoaz == 3'b000))
             | (xwk7fm0 & (ljxpmbsqoaz == 3'b11) & (~fvz__7_m))
             | (xwk7fm0 & (ljxpmbsqoaz == 3'b10) &  fvz__7_m))
             & (~ilnqntxsop67);

wire ongdihwv8i = ( ((ljxpmbsqoaz == 3'b10) & xwk7fm0 & (~fvz__7_m))
               | ((ljxpmbsqoaz == 3'b01) & xwk7fm0)
               | ((ljxpmbsqoaz == 3'b11) & xwk7fm0 &  fvz__7_m))
               & (~ilnqntxsop67);

wire dnlvg2ua7g18 = 1'b0;
wire [62:0] q066f9sz1wy28dm = {{11{1'b0}}, {52{1'b0}}};
wire [30:0] zmeqgppv3pjswx = {{8{1'b0}}, {23{1'b0}}};


wire wcose8catghq = (bn60jfu_ewb | ongdihwv8i | dnlvg2ua7g18 | ilnqntxsop67);
wire r_7ptkidm = ~wcose8catghq;



wire [31:0] pc7dgw1nyhsdlr6y = ({32{bn60jfu_ewb   }} & {fvz__7_m, 31'h7F80_0000})
                             | ({32{ongdihwv8i    }} & {fvz__7_m, 31'h7F7F_FFFF})
                             | ({32{dnlvg2ua7g18    }} & {fvz__7_m, zmeqgppv3pjswx} )
                             | ({32{ilnqntxsop67 }} & powr[31:0]);

wire [63:0] n4xfku6k9juladeoa8c7 = ({64{bn60jfu_ewb  }} & {fvz__7_m, 63'h7FF0_0000_0000_0000})
                             | ({64{ongdihwv8i   }} & {fvz__7_m, 63'h7FEF_FFFF_FFFF_FFFF})
                             | ({64{dnlvg2ua7g18   }} & {fvz__7_m, q066f9sz1wy28dm          })
                             | ({64{ilnqntxsop67}} & powr);

wire [31:0] aiv5a9vlee68jk2yz = v12nwpm6b862ua[31:0];
wire [63:0] twyqo8fo2b3rppnpc = et2w664wl8r[63:0];


wire [31:0] f6xnozunpt = ({32{r_7ptkidm}} & aiv5a9vlee68jk2yz) | ({32{wcose8catghq}} & pc7dgw1nyhsdlr6y);
wire [63:0] u8jj29yi9jywk = ({64{r_7ptkidm}} & twyqo8fo2b3rppnpc) | ({64{wcose8catghq}} & n4xfku6k9juladeoa8c7);


wire [63:0] zbggcho1tucaz8fe;
wire [63:0] mca66cdvg_a98;
wire[5:0] ksqmfb7wfr_46ha_9x;

assign zbggcho1tucaz8fe[31:00] = (ilnqntxsop67 | y_zx8qolynd) ? u8jj29yi9jywk[31:0] : f6xnozunpt; 
assign zbggcho1tucaz8fe[63:32] = u8jj29yi9jywk[63:32] ;

wire[5:0] im68j6624nd6dpsy_611n = {1'b0, wb3pal8jhelc__t0, fipd_e_m294cc01e54bb, ixn122itx74ljf0e8dk, gp5nsjv6nris3nx7zm2, a_xtsojke05dnao};
wire[5:0] q1kl83tne5qcxf9cii2 =ilnqntxsop67 ? ey7de2vqxx : im68j6624nd6dpsy_611n;

assign xptd3f_t3cg5 = mca66cdvg_a98[31:00];
assign r4nxuj5xq_p = (~ux0s4l13o) ? 32'hFFFFFFFF : mca66cdvg_a98[63:32];

assign g2gmxy0taet_c61t = ksqmfb7wfr_46ha_9x;

ux607_gnrl_dffl #(64) xjfxz4rlehtsff1kcgrr( c6yo0on_3i, zbggcho1tucaz8fe,mca66cdvg_a98, gf33atgy, ru_wi);
ux607_gnrl_dffl #(6) jzh9lnm168c5qcozbvdph( c6yo0on_3i, q1kl83tne5qcxf9cii2,ksqmfb7wfr_46ha_9x, gf33atgy, ru_wi);

endmodule






module vz0a9sv0gw3w9am21j3ue6qp (
    output eypswghjg4a5o,

    input           hsxngq7neaj187i70n, 
    output          a2kaizumm2cx6tylhsg, 
    output [32-1:0] ww3enujjopw1vz9, 
    output [5-1:0] s1910mdw_o4lix, 
    output [4-1:0] ogfp_yyiz39, 
    output [32-1:0] jk8q8hf4c7enovxal, 

    input [63:0] miesq8xb,
    input [63:0] l5o8oedt,
    input i88m5b2zjh,
    input kmku5oaqfkit5,
    input jaio35_tn,
    input [2:0] ncf9rmc,
    input pg_nt6lde,
    output tbqq6db__lsqi,
    input [4-1:0] vu2b4w8p, 

    input gf33atgy,
    input ru_wi
);

wire [4-1:0] nnvn3q = {{4-4{1'b0}},vu2b4w8p};
wire y7s8lz156ibl;
wire ilnqntxsop67;
wire [63:0] powr;
wire [5:0]  g2gmxy0taet_c61t;
wire [5:0]  ey7de2vqxx;







wire q1hmdngt1v4x5958y;
wire [4-1:0] ju_5ti46ayy7vdw;
assign ogfp_yyiz39 = ju_5ti46ayy7vdw[4-1:0] ;
assign s1910mdw_o4lix = {
    g2gmxy0taet_c61t[0],
    g2gmxy0taet_c61t[1],
    g2gmxy0taet_c61t[2],
    g2gmxy0taet_c61t[3],
    g2gmxy0taet_c61t[4]}; 


wire [4:0] gd2wkhivb2;        
wire yh0oeg399pvwaqg13;
wire mg9we1s5d77ws;
wire bhmxsiib6;
wire vawmftolubc5;
wire c6yo0on_3i;
wire cl_ffrx4sh;
wire bp_c30xz;
wire rg10e3avkel ;

wire [5:0] a0_2x3l9euvn1ixa6;
wire [5:0] dvmjxjsqko9mdgn;
wire [63:0] zc_86cgz6a;
wire [63:0] dqspoelekb5d;
wire m0e2_guluq90ndzyt;

wire q02bklc;
wire nv_meva_f5;
wire lzbquud;
wire y_zx8qolynd;
wire ux0s4l13o;

jgdiavy4q4l1fecbof09xfij9 rd92yzmw5906c8cpt2 ( 
        .xptd3f_t3cg5          (ww3enujjopw1vz9),
        .r4nxuj5xq_p          (jk8q8hf4c7enovxal),
        .g2gmxy0taet_c61t     (g2gmxy0taet_c61t),
        .yh0oeg399pvwaqg13  (yh0oeg399pvwaqg13),
        .ie_pkh83p_8          (zc_86cgz6a[63:32]),
        .r1pjdyql2t19          (dqspoelekb5d[63:32]),
        .e3oq_fn1szj61          (zc_86cgz6a[31:00]),
        .wswzu1c4y6et          (dqspoelekb5d[31:00]),
        .a0_2x3l9euvn1ixa6      (a0_2x3l9euvn1ixa6),
        .dvmjxjsqko9mdgn      (dvmjxjsqko9mdgn),
        .m0e2_guluq90ndzyt  (m0e2_guluq90ndzyt ),
        .tqpavw30         (jaio35_tn),
        .kjauvty_w            (i88m5b2zjh),
        .j5crtzpyh           (kmku5oaqfkit5),
        .rg10e3avkel           (rg10e3avkel),
        .cl_ffrx4sh          (cl_ffrx4sh),
        .bp_c30xz          (bp_c30xz),
        .bhmxsiib6          (bhmxsiib6),
        .vawmftolubc5          (vawmftolubc5),
        .c6yo0on_3i          (c6yo0on_3i),
        .ilnqntxsop67   (ilnqntxsop67),
        .powr         (powr),
        .ey7de2vqxx  (ey7de2vqxx),
        .gd2wkhivb2        (gd2wkhivb2),
        .n5900it0gq9hnv         (ncf9rmc),
        .q02bklc    (q02bklc),
        .nv_meva_f5    (nv_meva_f5),
        .lzbquud    (lzbquud),
        .y_zx8qolynd    (y_zx8qolynd),
        .ux0s4l13o    (ux0s4l13o),
        .gf33atgy           (gf33atgy),
        .ru_wi         (ru_wi)
);

cjellcyv3z8y1t_ad hlob51dykvac9l(
        .miesq8xb                     (miesq8xb ),
        .l5o8oedt                     (l5o8oedt ),
        .ohq4d3f_j                     (64'b0 ),
        .pg_nt6lde                (pg_nt6lde), 
        .i88m5b2zjh                  (i88m5b2zjh),
        .jaio35_tn               (jaio35_tn),
        .vu2b4w8p              (nnvn3q),
        .y7s8lz156ibl  (y7s8lz156ibl),
        .powr           (powr),
        .ey7de2vqxx    (ey7de2vqxx),
        .zc_86cgz6a             (zc_86cgz6a),
        .dqspoelekb5d             (dqspoelekb5d),
        .a0_2x3l9euvn1ixa6        (a0_2x3l9euvn1ixa6),
        .dvmjxjsqko9mdgn        (dvmjxjsqko9mdgn),
        .m0e2_guluq90ndzyt    (m0e2_guluq90ndzyt ),
        .q1hmdngt1v4x5958y(q1hmdngt1v4x5958y),
        .mg9we1s5d77ws          (mg9we1s5d77ws),
        .cl_ffrx4sh            (cl_ffrx4sh),
        .gf33atgy                     (gf33atgy),
        .ru_wi                 (ru_wi)
);

ur945ax08pidlnz7_o24hdlr uk4e2ldc0ahwf(
        .baefqz_y6q1d7            (hsxngq7neaj187i70n),
        .jdo6mn_o05686d2cl           (a2kaizumm2cx6tylhsg),
        .ju_5ti46ayy7vdw               (ju_5ti46ayy7vdw),
        .eypswghjg4a5o             (eypswghjg4a5o),

        .cl_ffrx4sh             (cl_ffrx4sh),
        .bp_c30xz             (bp_c30xz),
        .rg10e3avkel              (rg10e3avkel),
        .bhmxsiib6             (bhmxsiib6),
        .vawmftolubc5             (vawmftolubc5),
        .c6yo0on_3i             (c6yo0on_3i),
        .mg9we1s5d77ws           (mg9we1s5d77ws),
        .am_rltp_3w              (tbqq6db__lsqi),
        .p_rmwvx8z               (nnvn3q),
        .vwd0ug0ks5l                 (pg_nt6lde),
        .uu3yswtakfh              (jaio35_tn),
        .gd2wkhivb2           (gd2wkhivb2),
        .yh0oeg399pvwaqg13     (yh0oeg399pvwaqg13),
        .y7s8lz156ibl   (y7s8lz156ibl),
        .ilnqntxsop67   (ilnqntxsop67),
        .q02bklc    (q02bklc),
        .nv_meva_f5    (nv_meva_f5),
        .lzbquud    (lzbquud),
        .y_zx8qolynd    (y_zx8qolynd),
        .ux0s4l13o    (ux0s4l13o),
        .gf33atgy                      (gf33atgy),
        .ru_wi                  (ru_wi)
);


endmodule

module o_6c7gxntcc9ta0bisv_(
  input [56:0] rydw,
  input [56:0] d4y,
  output ust6kl,
  output p2yjv_h8o ,
  output v2f5pmhic4
);

wire [3:0] wv9;
assign wv9 = rydw[56-1:56-4] + d4y[56-1:56-4] ;
assign ust6kl = ~wv9[3] ;
assign p2yjv_h8o = &wv9[3:0];
assign v2f5pmhic4 = wv9[3] & ~(wv9[2] & wv9[1] & wv9[0]) ;

endmodule








module cjellcyv3z8y1t_ad (
  input [63:0] miesq8xb,
  input [63:0] l5o8oedt,
  input [63:0] ohq4d3f_j,
  input pg_nt6lde,
  input i88m5b2zjh,
  input jaio35_tn,
  input [4-1:0] vu2b4w8p,
  
  output y7s8lz156ibl,
  output [63:0] powr,
  output [5:0] ey7de2vqxx,
  output [63:0] zc_86cgz6a,
  output [63:0] dqspoelekb5d,
  output [5:0] a0_2x3l9euvn1ixa6,
  output [5:0] dvmjxjsqko9mdgn,
  output m0e2_guluq90ndzyt,
  output q1hmdngt1v4x5958y,
  
  input mg9we1s5d77ws,
  input cl_ffrx4sh,
  input gf33atgy,
  input ru_wi
);



wire exiyz1djym8k = i88m5b2zjh & (jaio35_tn ? (miesq8xb[51:0] == 52'b0) : (miesq8xb[22:0] == 23'b0));
wire plon1c5v = jaio35_tn ? (l5o8oedt[51:0] == 52'b0) : (l5o8oedt[22:0] == 23'b0);
wire i48mlnnyzur = i88m5b2zjh & (jaio35_tn ? (miesq8xb[62:52] == 11'h000) : (miesq8xb[30:23] == 8'h00));
wire td1glnmfo2 = jaio35_tn ? (l5o8oedt[62:52] == 11'h000) : (l5o8oedt[30:23] == 8'h00);

wire zpep1bwfqe77i4 = i88m5b2zjh & (jaio35_tn ? (miesq8xb[62:52] == 11'h7FF) : (miesq8xb[30:23] == 8'hFF));
wire zr0n8j2nw5z = jaio35_tn ? (l5o8oedt[62:52] == 11'h7FF) : (l5o8oedt[30:23] == 8'hFF);

wire h6m9q2omm = i88m5b2zjh & (jaio35_tn ? miesq8xb[51] : miesq8xb[22]);
wire yl2yeycmx = zpep1bwfqe77i4 & (~exiyz1djym8k) & (~h6m9q2omm);
wire om1oy2pjja66r = zpep1bwfqe77i4 & (~exiyz1djym8k) & h6m9q2omm;

wire ly5v6vrmdv = jaio35_tn ? l5o8oedt[51] : l5o8oedt[22];
wire w20nt86h9cw9d = zr0n8j2nw5z & (~plon1c5v) & (~ly5v6vrmdv);
wire uuc63syvkcf = zr0n8j2nw5z & (~plon1c5v) & ly5v6vrmdv;

wire dmr_pwxw617e = om1oy2pjja66r | yl2yeycmx;
wire slze1vivbq = uuc63syvkcf | w20nt86h9cw9d;

wire zipbe43g9h7 = zpep1bwfqe77i4 & exiyz1djym8k;
wire dv4hotijmb6g = zr0n8j2nw5z & plon1c5v;

wire b284for6 = i48mlnnyzur & (~exiyz1djym8k);
wire uojp70 = td1glnmfo2 & (~plon1c5v);

wire cpgs9inefc3sa = (i48mlnnyzur & exiyz1djym8k);
wire ugf0mrh7o7c = (td1glnmfo2 & plon1c5v);

wire bkzlmzat = i88m5b2zjh & (jaio35_tn ? miesq8xb[63] : miesq8xb[31]);   
wire qxzlt1eb = jaio35_tn ? l5o8oedt[63] : l5o8oedt[31];


wire mmq8l6gaf9c5kd6or = yl2yeycmx | (om1oy2pjja66r & (~w20nt86h9cw9d));
wire jj87229baeh4z = ((~yl2yeycmx) & w20nt86h9cw9d) | ((~dmr_pwxw617e) & uuc63syvkcf);
wire m1__badzg8bj5 = (zipbe43g9h7 & dv4hotijmb6g) | (cpgs9inefc3sa & ugf0mrh7o7c);

wire t2z8gbhpar6y  = (~dmr_pwxw617e) & (~slze1vivbq) & ((zipbe43g9h7 & (~dv4hotijmb6g)) | ((ugf0mrh7o7c ) &  (~cpgs9inefc3sa)));
wire wslyx6wdh2zscnmk = (~dmr_pwxw617e) & (~slze1vivbq) & (((~zipbe43g9h7) & dv4hotijmb6g) | ((~ugf0mrh7o7c)  & ( cpgs9inefc3sa)));

wire ik1ovu7aet8bjry = qxzlt1eb & ugf0mrh7o7c;
wire z4n1us1p6n_3da1tpth = slze1vivbq;
wire aisf7ki_o37x4xk = qxzlt1eb & (~ugf0mrh7o7c) & (~slze1vivbq);
wire lcfrs3q9qjoj = (~qxzlt1eb) & dv4hotijmb6g;
wire sgv36cvy1bnwx = ugf0mrh7o7c;

wire q4zw_uqzjk96exkjn = i88m5b2zjh & mmq8l6gaf9c5kd6or;
wire bis3cjeu7szfz61gi60gj = i88m5b2zjh & jj87229baeh4z;
wire oe2dqsjscnhx5q2kxc_hb = i88m5b2zjh & m1__badzg8bj5;
wire b7usi4u5ajquale1 = t2z8gbhpar6y & i88m5b2zjh;
wire mphlgmk35t3xh67wfy = wslyx6wdh2zscnmk & i88m5b2zjh;

wire pw7tc77f4uzzmhyp9cm4 = (~i88m5b2zjh) & z4n1us1p6n_3da1tpth;
wire muuhv62bcaq7vzqb4g06z = (~i88m5b2zjh) & aisf7ki_o37x4xk;
wire ad6gjmd_j2lh0kp9o  = lcfrs3q9qjoj  & (~i88m5b2zjh);
wire qr_6dj7opoc_4zsralc84 = sgv36cvy1bnwx & (~i88m5b2zjh);

wire rc6rk1liyqaw = bkzlmzat ^ qxzlt1eb;
wire rh2obkqt47c2v = (i88m5b2zjh & rc6rk1liyqaw & (~oe2dqsjscnhx5q2kxc_hb)) 
              | ((~i88m5b2zjh) & ik1ovu7aet8bjry & (~muuhv62bcaq7vzqb4g06z))  ;
wire f95e667o_1elu = (q4zw_uqzjk96exkjn & bkzlmzat) 
                  | (bis3cjeu7szfz61gi60gj & qxzlt1eb) 
                  | (pw7tc77f4uzzmhyp9cm4 & qxzlt1eb);

wire k104r9vcv3mkys = bis3cjeu7szfz61gi60gj;
wire h528f4qoy1rfu7s4yn = q4zw_uqzjk96exkjn | pw7tc77f4uzzmhyp9cm4; 
wire yrbpeeob2ll34ssu = oe2dqsjscnhx5q2kxc_hb | muuhv62bcaq7vzqb4g06z;

wire b39ic_jw7xqj  = b7usi4u5ajquale1  | ad6gjmd_j2lh0kp9o ;
wire evz1mi2gw18u5d = mphlgmk35t3xh67wfy | qr_6dj7opoc_4zsralc84;

wire [63:0] k28ab74q0b9wb = jaio35_tn ? {miesq8xb[63:52], 1'b1, miesq8xb[50:0]} : {32'b0, miesq8xb[31:23], 1'b1, miesq8xb[21:0]} ;
wire [63:0] f8sy6ibyoem6 = jaio35_tn ? {l5o8oedt[63:52], 1'b1, l5o8oedt[50:0]} : {32'b0, l5o8oedt[31:23], 1'b1, l5o8oedt[21:0]} ;

wire [32-1:0] e5otgqgjkm78gyd = 32'h7FC00000;
wire [64-1:0] k7gcz3dfv8 = 64'h7FF80000_00000000;

wire [31:0] bq2tf7lb2o= ({32{h528f4qoy1rfu7s4yn}} & e5otgqgjkm78gyd)
                  | ({32{k104r9vcv3mkys}} & e5otgqgjkm78gyd)
                  | ({32{yrbpeeob2ll34ssu}} & e5otgqgjkm78gyd)
                  | ({32{b39ic_jw7xqj  }} & {rh2obkqt47c2v, 8'hFF, 23'b0})
                  | ({32{evz1mi2gw18u5d }} & {rh2obkqt47c2v, 8'h00, 23'b0});

wire [63:0] lvgamcgahrm= ({64{h528f4qoy1rfu7s4yn}} & k7gcz3dfv8)
                  | ({64{k104r9vcv3mkys}} & k7gcz3dfv8)
                  | ({64{yrbpeeob2ll34ssu}} & k7gcz3dfv8)
                  | ({64{b39ic_jw7xqj  }} & {rh2obkqt47c2v, 11'h7FF, 52'b0})
                  | ({64{evz1mi2gw18u5d }} & {rh2obkqt47c2v, 11'h000, 52'b0});

assign y7s8lz156ibl = (ugf0mrh7o7c | 
                    (cpgs9inefc3sa & i88m5b2zjh) |
                    dv4hotijmb6g |
                    (zipbe43g9h7 & i88m5b2zjh) |
                    slze1vivbq |
                    (dmr_pwxw617e & i88m5b2zjh) |
                    ((~i88m5b2zjh) & qxzlt1eb));

wire d7zrtfixg4j = (~dmr_pwxw617e) & (~slze1vivbq) & (ugf0mrh7o7c & (~cpgs9inefc3sa) & (~zipbe43g9h7));
wire ycxzcgbh_qi = yl2yeycmx | w20nt86h9cw9d | (zipbe43g9h7 & dv4hotijmb6g) | (cpgs9inefc3sa & ugf0mrh7o7c);
wire wsbraq8wt2jt8vy1q = w20nt86h9cw9d | qxzlt1eb & (~ugf0mrh7o7c) & (~slze1vivbq); 

wire rquiw3t80u1d = d7zrtfixg4j & i88m5b2zjh; 
wire f9lqman5 = (i88m5b2zjh & ycxzcgbh_qi) | ((~i88m5b2zjh) & wsbraq8wt2jt8vy1q); 

wire [5:0] po7otfo5au= {1'b0, 3'b0, rquiw3t80u1d, f9lqman5};


wire [63:0] ab6pksukst = (jaio35_tn) ? lvgamcgahrm : {32'b0, bq2tf7lb2o};

wire [5:0] o2vx0pkre9qn65j5x;
wire [5:0] p8py2x6fkwhrya4vj;

wire [63:0] cw_oxt7ji4e4kc46 = jaio35_tn ? {1'b0,miesq8xb[51:0],11'h0}:{1'b0,miesq8xb[22:0],40'h0};
wire [63:0] lva5491u_hlrhnda = jaio35_tn ? {1'b0,l5o8oedt[51:0],11'h0}:{1'b0,l5o8oedt[22:0],40'h0};

xh5dey_d_oxo365f0d85q3d #(.onr7l(64),.hw3qvr(6)) jgwf_lj0ajz5m (.bjh(cw_oxt7ji4e4kc46), .ht70(o2vx0pkre9qn65j5x));
xh5dey_d_oxo365f0d85q3d #(.onr7l(64),.hw3qvr(6)) j7_ojcrh1awubkk (.bjh(lva5491u_hlrhnda), .ht70(p8py2x6fkwhrya4vj));

wire [63:0] mtww7c_hh26s4p692f =  {miesq8xb[63:32],miesq8xb[31],(b284for6 ? 8'b1:miesq8xb[30:23]), miesq8xb[22:0]} ;
wire [63:0] ilmxwyolncb7udp4 =  {l5o8oedt[63:32],l5o8oedt[31],(uojp70 ? 8'b1:l5o8oedt[30:23]), l5o8oedt[22:0]} ;
wire [63:0] bzqw10cpiymnf3s =  {miesq8xb[63],(b284for6 ? 11'b1:miesq8xb[62:52]), miesq8xb[51:0]} ;
wire [63:0] v7coqk_qc6b66s4aj50 =  {l5o8oedt[63],(uojp70 ? 11'b1:l5o8oedt[62:52]), l5o8oedt[51:0]} ;

wire [63:0] dlugxssmfh7goc = jaio35_tn ? bzqw10cpiymnf3s :mtww7c_hh26s4p692f;
wire [63:0] f7pma6bl69r4 = jaio35_tn ? v7coqk_qc6b66s4aj50 :ilmxwyolncb7udp4;

wire [63:0] vbu3miugy3;
wire [63:0] yebzb3y44t4b;

wire [5:0] mibv81vx47ongia_dpmtvtaz6=o2vx0pkre9qn65j5x;
wire [5:0] kbmzaxhpk5ckj_y319jic5r8x=p8py2x6fkwhrya4vj;
wire [5:0] fphl1_5u8f_qpcvhl6fo;
wire [5:0] m2bq98uxnqwav69pfary6;
wire jir8l7e5c7nm;
wire pyf7pjru1zz;
wire o_h1gf_gxagl;
wire flbjy_dd7ep;

ux607_gnrl_dffl #(64) kehgli1( mg9we1s5d77ws, ab6pksukst, powr, gf33atgy, ru_wi);
ux607_gnrl_dffl #(6) g1lvwcp873sbdbk( mg9we1s5d77ws, po7otfo5au,ey7de2vqxx, gf33atgy, ru_wi);
ux607_gnrl_dffl #(1) iyeqgl1s31gk6ernkpus2qu( mg9we1s5d77ws, (b284for6|uojp70),q1hmdngt1v4x5958y, gf33atgy, ru_wi);
ux607_gnrl_dffl #(64) sng7e8gzmx2b4gt7( cl_ffrx4sh, dlugxssmfh7goc,vbu3miugy3, gf33atgy, ru_wi);
ux607_gnrl_dffl #(64) j10a001ia9dq5( cl_ffrx4sh, f7pma6bl69r4,yebzb3y44t4b, gf33atgy, ru_wi);
ux607_gnrl_dffl #(6) kwmr3_8q08cz_30f2kmd6w7( cl_ffrx4sh, mibv81vx47ongia_dpmtvtaz6,fphl1_5u8f_qpcvhl6fo, gf33atgy, ru_wi);
ux607_gnrl_dffl #(6) bl_4vblb230siiv0qyxfpl2aura( cl_ffrx4sh, kbmzaxhpk5ckj_y319jic5r8x,m2bq98uxnqwav69pfary6, gf33atgy, ru_wi);

ux607_gnrl_dffl #(1) w0bm42k6daje44m8a( cl_ffrx4sh, b284for6,jir8l7e5c7nm, gf33atgy, ru_wi);
ux607_gnrl_dffl #(1) v8agl0tk3hao4o9wb( cl_ffrx4sh, uojp70,pyf7pjru1zz, gf33atgy, ru_wi);

ux607_gnrl_dffl #(1) mj6qspy7ew431hzojp( cl_ffrx4sh, jaio35_tn,o_h1gf_gxagl, gf33atgy, ru_wi);
ux607_gnrl_dffl #(1) k6t3jxcrxi_7kt8oli81( cl_ffrx4sh, i88m5b2zjh,flbjy_dd7ep, gf33atgy, ru_wi);


assign a0_2x3l9euvn1ixa6 = ({6{flbjy_dd7ep & jir8l7e5c7nm}} & fphl1_5u8f_qpcvhl6fo);
assign dvmjxjsqko9mdgn = ({6{pyf7pjru1zz}} & (m2bq98uxnqwav69pfary6));

wire [51:0] znaxifrxzp2mv_ = vbu3miugy3[51:0] << ({6{jir8l7e5c7nm}}&fphl1_5u8f_qpcvhl6fo);

wire [51:0] gmzx2ys6ryuhv02ayms;
wire xdlb48kf9qu38lv_z9yq7xw;

assign {xdlb48kf9qu38lv_z9yq7xw,gmzx2ys6ryuhv02ayms} =
    {1'b0,yebzb3y44t4b[51:0]} << ({6{pyf7pjru1zz}}&m2bq98uxnqwav69pfary6);

wire n3a40hv19aa9pqdlqjd8 = (~m2bq98uxnqwav69pfary6[0]);

wire [51:0] rwf8r3e3xddregnvp7m =gmzx2ys6ryuhv02ayms[51:0];

wire [22:0] d4muc9bqeo9oj1 = znaxifrxzp2mv_[22:0];
wire [22:0] ge185olj9mlnsq = rwf8r3e3xddregnvp7m[22:0]; 

wire [63:0] khk2coia6gz8e4 = {vbu3miugy3[63:32], vbu3miugy3[31], vbu3miugy3[30:23], d4muc9bqeo9oj1[22:0]} ;
wire [63:0] tzza542k8ckdfy8 = {yebzb3y44t4b[63:32], yebzb3y44t4b[31], yebzb3y44t4b[30:23], ge185olj9mlnsq[22:0]} ;
wire [63:0] dq8rdqkacekra6n = {vbu3miugy3[63], vbu3miugy3[62:52], znaxifrxzp2mv_[51:0]} ;
wire [63:0] daird_nrpsu = {yebzb3y44t4b[63], yebzb3y44t4b[62:52], rwf8r3e3xddregnvp7m[51:0]} ;

assign zc_86cgz6a = (o_h1gf_gxagl) ? dq8rdqkacekra6n : khk2coia6gz8e4;
assign dqspoelekb5d = (o_h1gf_gxagl) ? daird_nrpsu : tzza542k8ckdfy8;

wire [10:0] yruj_3_m8kmx8 = o_h1gf_gxagl ? yebzb3y44t4b[62:52] : {3'b0,yebzb3y44t4b[30:23]};
assign m0e2_guluq90ndzyt = pyf7pjru1zz ? n3a40hv19aa9pqdlqjd8 : yruj_3_m8kmx8[0];


endmodule

    








module drpp7_8vqsgvijw(

 
  output  eypswghjg4a5o,

  
  
  
  
  input  cfk6xv54sxw51e,
  output ay4xay0aajxpqki,

  input  [64-1:0] rx7xp4yfzkxxwe,
  input  [64-1:0] yh6637l46fxr,
  input  [48-1:0] fx3oxnmunmg5,
  input  [4-1:0] ylzz2nmn2fx8vx,
  input  [3-1:0] i7mguch8rrz_acmgw,

  
  
  
  output o1ic53wzueq3rdj, 
  input  q5hfrt_ivi2var, 
  output [64-1:0] xw5sonra6wr1qw86is7,
  output [5-1:0] zghahb2tb_ksbg78bg4,
  output [4 -1:0] u3_iseqd_x1swj1y1ikzv,
  output aau8gpkszf2jvnjbmhfpm , 

  input  gf33atgy,
  input  ru_wi
  );

  wire nn8hi7fy9 = fx3oxnmunmg5[13:13];
  wire toc7itgvlx  = fx3oxnmunmg5[11:11   ];
  wire nna5gl9h5lo = fx3oxnmunmg5[12:12  ];
  wire [64-1:0] tcck0j = rx7xp4yfzkxxwe;
  wire [64-1:0] onuou7_ = nna5gl9h5lo ? rx7xp4yfzkxxwe : yh6637l46fxr;

  assign aau8gpkszf2jvnjbmhfpm = 1'b0; 

vz0a9sv0gw3w9am21j3ue6qp sgivryy6dpb7fckcoj8rwcwnu (
    .eypswghjg4a5o           (eypswghjg4a5o),
    .hsxngq7neaj187i70n     (q5hfrt_ivi2var),  
    .a2kaizumm2cx6tylhsg     (o1ic53wzueq3rdj),  
    .ww3enujjopw1vz9        (xw5sonra6wr1qw86is7[31:0]),
    .jk8q8hf4c7enovxal        (xw5sonra6wr1qw86is7[63:32]),
    .s1910mdw_o4lix         (zghahb2tb_ksbg78bg4),
    .ogfp_yyiz39          (u3_iseqd_x1swj1y1ikzv),

    .miesq8xb           (tcck0j),
    .l5o8oedt           (onuou7_),
    .jaio35_tn        (nn8hi7fy9),
    .i88m5b2zjh        (toc7itgvlx),
    .kmku5oaqfkit5       (nna5gl9h5lo),
    .ncf9rmc         (i7mguch8rrz_acmgw),
    .pg_nt6lde      (cfk6xv54sxw51e),
    .tbqq6db__lsqi      (ay4xay0aajxpqki),
    .vu2b4w8p       (ylzz2nmn2fx8vx),

    .gf33atgy           (gf33atgy),
    .ru_wi       (ru_wi) 
);


endmodule

module ikddk6f6fc0_2t0g5wt #(
    parameter onr7l = 106 
)(
  input [onr7l-1:0] frgfco,
  input [onr7l-1:0] ii,
  input [onr7l-1:0] fij51v,
  input [onr7l-1:0] cuzhl9,
  output [onr7l-1:0] c,
  output [onr7l-1:0] s 
);

   wire [onr7l-1:0] i885 = (frgfco & ii) | (ii & fij51v) | (frgfco & fij51v);
   wire [onr7l-1:0] smqrocit = {i885[onr7l-2:0], 1'b0};

   wire [onr7l-1:0] tqxp_8 = smqrocit ^ cuzhl9;
   wire [onr7l-1:0] ddaxu87 = (frgfco ^ ii) ^ fij51v;

   assign s = tqxp_8 ^ ddaxu87;

   wire [onr7l-1:0] hgtxv = (ddaxu87 & cuzhl9) |  (cuzhl9 & smqrocit) | (smqrocit & ddaxu87);

   assign c = {hgtxv[onr7l-2:0], 1'b0};

endmodule

module j3aa8h4yagvjsr416mg #(
  parameter onr7l = 106 
)(
  input [onr7l-1:0] frgfco,
  input [onr7l-1:0] ii,
  input [onr7l-1:0] fij51v,
  output [onr7l-1:0] c,
  output [onr7l-1:0] s 
);

assign s = (frgfco ^ ii) ^ fij51v;

wire [onr7l-1:0] oz7_y5 = (frgfco & ii) | (frgfco & fij51v) | (ii & fij51v);

assign c = {oz7_y5[onr7l-2:0], 1'b0};

endmodule

module el7n_zz16sk_ntvue9v (
  input l,
  input g,
  input r,
  input s,
  input ly53de,
  input [2:0] nfj6b,
  output f6dc_rhcaz 
);

wire c5gschl9oda1a = 1'b0 ;

wire cv9u8eujnn7 = ~ly53de & (g | r | s) ;
wire vqt52loy53 = ly53de & (g | r | s) ;
wire hmkm4bg1ix3fqz  = g & (l | r | s) ;
wire bwwwfquqiwv4m  = g;

assign f6dc_rhcaz = (nfj6b == 3'b000)&hmkm4bg1ix3fqz 
              |(nfj6b == 3'b011)&cv9u8eujnn7 
              |(nfj6b == 3'b010)&vqt52loy53
              |(nfj6b == 3'b001)&1'b0  
              |(nfj6b == 3'b100)&bwwwfquqiwv4m;

endmodule








module iojbcv7tg90u(

 
  output  g9ruu8swf4b_,

  
  
  
  
  input  aa9_kdx_kb35fx,
  output z30wkcif1o8is5w9,

  input  [64-1:0] a4_acuaz1sfb5,
  input  [64-1:0] q3ek793hh,
  input  [48-1:0] z1oylnyp4ryl4v,
  input  [4-1:0] du24en2x_2qkjfw,
  input  [2:0] eyaonb2nm4ox,

  
  
  
  output ycjcjdm1fjmdo_j, 
  input  j0s42ouqf5zv1a, 
  output [64-1:0] bqc9gh1yogik7q5r,
  output [5-1:0] dd4hyq5oe67rhyvoye,
  output [4 -1:0] k4euvut15h32iq7j,
  output b60gak_58icq19sfs_ , 

  input  gf33atgy,
  input  ru_wi
  );

  wire zxo6khy1ic0d4p1  = z1oylnyp4ryl4v[19:19 ];
  wire wzf5u5qgu_9jg2wuf = z1oylnyp4ryl4v[20:20];
  wire pfo9ob4rnnslccuy  = z1oylnyp4ryl4v[21:21 ];
  wire akeh5qohkbjhf = z1oylnyp4ryl4v[22:22];
  wire ca2zy5rakjh1  = z1oylnyp4ryl4v[23:23 ];
  wire mjbj7q63yu0c  = z1oylnyp4ryl4v[24:24 ];
  wire kimruawu3hx2609k  = z1oylnyp4ryl4v[25:25 ];
  wire aow77uvoxp9i = z1oylnyp4ryl4v[26:26];
  wire sahahgr77v6  = z1oylnyp4ryl4v[27:27 ];
  wire rtxu4mywvri6 = z1oylnyp4ryl4v[28:28];
  wire gmtcz_y3rutu5mz  = z1oylnyp4ryl4v[30:30 ];
  wire e540r67hz2u7 = z1oylnyp4ryl4v[31:31];
  wire bpdqvi5i6n95qe7  = z1oylnyp4ryl4v[32:32 ];
  wire a6mdgi0ed1s_kbe = z1oylnyp4ryl4v[33:33];
  wire v4pl9zyada0sp  = z1oylnyp4ryl4v[34:34 ];
  wire rj6dvlwj0iy2tf7o = z1oylnyp4ryl4v[35:35];
  wire rln9tn6f_5c  = z1oylnyp4ryl4v[36:36 ];
  wire ydsyvkyqns88ata = z1oylnyp4ryl4v[37:37];

  wire v659v2hvrtej = zxo6khy1ic0d4p1;
  wire p940nw4duiie64 = wzf5u5qgu_9jg2wuf;
  wire ersv4d_m80ir1 = kimruawu3hx2609k;
  wire lc9pop79cuks = aow77uvoxp9i;
  wire af8gggx2rbk5w = pfo9ob4rnnslccuy;
  wire z9ydb68fp_la3j = akeh5qohkbjhf;
  wire im1jxeoei8g = sahahgr77v6;
  wire c2o9xduz06 = rtxu4mywvri6;
  wire azpnhv65b4= gmtcz_y3rutu5mz;
  wire ji57bityrdt= e540r67hz2u7;
  wire ex14gbip3a= v4pl9zyada0sp;
  wire f_xw6g_ldgz= rj6dvlwj0iy2tf7o;
  wire cix9qipqelc7k= bpdqvi5i6n95qe7;
  wire wpio23m13to3o0= a6mdgi0ed1s_kbe;
  wire u9bwc77pa3= rln9tn6f_5c;
  wire k937n2wbqgq= ydsyvkyqns88ata;
  wire ayc3vpo7   = ca2zy5rakjh1;
  wire goy441jl   = mjbj7q63yu0c;

  wire nn8hi7fy9 = z1oylnyp4ryl4v[29:29];

  wire fp36oxlnph;
  wire mzfgvfleu = 
            v659v2hvrtej 
          | p940nw4duiie64 
          | ersv4d_m80ir1 
          | lc9pop79cuks 
          | af8gggx2rbk5w 
          | z9ydb68fp_la3j 
          | im1jxeoei8g 
          | c2o9xduz06 
          | azpnhv65b4 
          | ji57bityrdt 
          | ex14gbip3a 
          | f_xw6g_ldgz 
          | cix9qipqelc7k 
          | wpio23m13to3o0 
          | u9bwc77pa3 
          | k937n2wbqgq 
          | ayc3vpo7   
          | goy441jl  ;


  wire [64-1:0] nrw_p_xi41_m;
  wire [64-1:0] uzjy58pkyanv;
  wire [48-1:0] ldd0t9ec4ucnlz86;
  wire [4-1:0] jqtb_mr6nt1uro;
  wire [3-1:0] xs0g801ygdou7f9l5i;

  ux607_gnrl_dfflr #(64         )v8bf171imwh8xq   (aa9_kdx_kb35fx, a4_acuaz1sfb5[64-1:0] , nrw_p_xi41_m , gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(64         )e19tf5ll13t_ebyn  (aa9_kdx_kb35fx, q3ek793hh[64-1:0] , uzjy58pkyanv , gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(48)npgohsqmldped4rp  (aa9_kdx_kb35fx, z1oylnyp4ryl4v, ldd0t9ec4ucnlz86, gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(4   )arp3z5w2l21jsi17   (aa9_kdx_kb35fx, du24en2x_2qkjfw, jqtb_mr6nt1uro, gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(3                  )w5g6z591t60kamo  (aa9_kdx_kb35fx, eyaonb2nm4ox, xs0g801ygdou7f9l5i, gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1                  )mn0yxx2od_mb   (aa9_kdx_kb35fx, mzfgvfleu,    fp36oxlnph,      gf33atgy, ru_wi);



  assign k4euvut15h32iq7j = jqtb_mr6nt1uro;

  ux607_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(1)
  ) q2m4di71ne6ce3 (
   .i_vld(aa9_kdx_kb35fx), 
   .i_rdy(z30wkcif1o8is5w9), 
   .i_dat(1'b0),
   .o_vld(ycjcjdm1fjmdo_j), 
   .o_rdy(j0s42ouqf5zv1a), 
   .o_dat(),
 
   .clk  (gf33atgy  ),
   .rst_n(ru_wi)  
  );

  assign g9ruu8swf4b_ = ycjcjdm1fjmdo_j;

  assign b60gak_58icq19sfs_ = 1'b0; 

  wire m7s5rkmh = ldd0t9ec4ucnlz86[29:29];
  wire nlb5566a2kkzrak  = (~m7s5rkmh) & ldd0t9ec4ucnlz86[11:11 ];
  wire t82iq62ywf1u_5 = (~m7s5rkmh) & ldd0t9ec4ucnlz86[12:12];
  wire byqkkp26xdsszd = (~m7s5rkmh) & ldd0t9ec4ucnlz86[13:13];
  wire l6qpfpq3ro_9gr = (~m7s5rkmh) & ldd0t9ec4ucnlz86[16:16];
  wire nxf52k3xp6im5o6p3 = (~m7s5rkmh) & ldd0t9ec4ucnlz86[17:17 ];
  wire gkj8ltdpe4tcqini4h = (~m7s5rkmh) & ldd0t9ec4ucnlz86[14:14 ];
  wire tr03xi8fsjspsc = (~m7s5rkmh) & ldd0t9ec4ucnlz86[18:18 ];
  wire va7j9_tx3li0xd = (~m7s5rkmh) & ldd0t9ec4ucnlz86[15:15 ];
  wire vdmyb8x4qmwi7on2  = m7s5rkmh & ldd0t9ec4ucnlz86[11:11 ];
  wire tfoxw8ia_xdt0 = m7s5rkmh & ldd0t9ec4ucnlz86[12:12];
  wire f128ccj13txxdwpl = m7s5rkmh & ldd0t9ec4ucnlz86[13:13];
  wire u72qi7gmhj37d_h5c = m7s5rkmh & ldd0t9ec4ucnlz86[16:16];

  wire [64-1:0] mbi1a;
  wire [5-1:0] taferz5nhfy1ttu;


  wire [64-1:0] ey8xno0w51z = a4_acuaz1sfb5 & {64{mzfgvfleu}};
  wire cr7bv45kj7l = aa9_kdx_kb35fx & mzfgvfleu;

  swhs3pkf0sfg9ix peq54p36so3aj9x4(
    .gf33atgy   (gf33atgy),
    .ru_wi (ru_wi),
    .cr7bv45kj7l (cr7bv45kj7l),
    .ticq8ng (ey8xno0w51z[63:32]),
    .y4a7pqq0kkz (ey8xno0w51z[31:0]),
    .v659v2hvrtej(v659v2hvrtej),
    .p940nw4duiie64(p940nw4duiie64),
    .af8gggx2rbk5w(af8gggx2rbk5w),
    .z9ydb68fp_la3j(z9ydb68fp_la3j),
    .ersv4d_m80ir1(ersv4d_m80ir1),
    .lc9pop79cuks(lc9pop79cuks),
    .im1jxeoei8g(im1jxeoei8g),
    .c2o9xduz06(c2o9xduz06),
    .ayc3vpo7  (ayc3vpo7  ),
    .goy441jl  (goy441jl  ),
    .azpnhv65b4(azpnhv65b4),
    .ji57bityrdt(ji57bityrdt),
    .cix9qipqelc7k(cix9qipqelc7k),
    .wpio23m13to3o0(wpio23m13to3o0),
    .ex14gbip3a(ex14gbip3a),
    .f_xw6g_ldgz(f_xw6g_ldgz),
    .u9bwc77pa3(u9bwc77pa3),
    .k937n2wbqgq(k937n2wbqgq),
    .vc529nuu(eyaonb2nm4ox),
    .uiwlxd (mbi1a),
    .adnx9wgdt2 (taferz5nhfy1ttu)
  );


  wire [9:0] tcfrqq029;
  wire yla1361h = (l6qpfpq3ro_9gr | u72qi7gmhj37d_h5c);
  wire [64-1:0] bzimv_ki4_0ft9e1 = nrw_p_xi41_m[64-1:0] & {64{yla1361h}};

  r5e39tculmqtcj5 tqa5p274nn_8fx10s(
    .ticq8ng (bzimv_ki4_0ft9e1[63:32]),
    .nn8hi7fy9 (m7s5rkmh),
    .y4a7pqq0kkz (bzimv_ki4_0ft9e1[31:0]),

    .uwkhmy2e_yju     (),
    .k1fnd9t0fsu     (),
    .la186rvvv7gcy   (),
    .kd65qo8qkm0kgmw     (),
    .a7atgbs19h1     (),
    .kzl0hy0qswsidji5   (),
    .boll1pzurodbj     (),
    .kt7mps652so     (),
    .em08qdw         (),
    .fij5gpv         (),

    .tcfrqq029 (tcfrqq029)
);

  wire [64-1:0] t3yzmt9i3dp5w7pnh;
  wire [64-1:0] vkkt61kb_gomf5;
  wire [64-1:0] vymyvujb_fnw9;
    assign t3yzmt9i3dp5w7pnh [32-2:0] = nrw_p_xi41_m[32-2:0];
    assign vkkt61kb_gomf5[32-2:0] = nrw_p_xi41_m[32-2:0];
    assign vymyvujb_fnw9[32-2:0] = nrw_p_xi41_m[32-2:0];
    assign t3yzmt9i3dp5w7pnh [32-1]   = m7s5rkmh ? nrw_p_xi41_m[32-1] : uzjy58pkyanv[32-1];
    assign vkkt61kb_gomf5[32-1]   = m7s5rkmh ? nrw_p_xi41_m[32-1] : (~uzjy58pkyanv[32-1]);
    assign vymyvujb_fnw9[32-1]   = m7s5rkmh ? nrw_p_xi41_m[32-1] : (nrw_p_xi41_m[32-1] ^ uzjy58pkyanv[32-1]);

    assign t3yzmt9i3dp5w7pnh [64-2:32] = m7s5rkmh ? nrw_p_xi41_m[64-2:32] : 31'h7FFF_FFFF;
    assign vkkt61kb_gomf5[64-2:32] = m7s5rkmh ? nrw_p_xi41_m[64-2:32] : 31'h7FFF_FFFF;
    assign vymyvujb_fnw9[64-2:32] = m7s5rkmh ? nrw_p_xi41_m[64-2:32] : 31'h7FFF_FFFF;
    assign t3yzmt9i3dp5w7pnh [64-1]    = m7s5rkmh ? uzjy58pkyanv[64-1]                       : 1'b1;
    assign vkkt61kb_gomf5[64-1]    = m7s5rkmh ? (~uzjy58pkyanv[64-1])                    : 1'b1;
    assign vymyvujb_fnw9[64-1]    = m7s5rkmh ? (nrw_p_xi41_m[64-1] ^ uzjy58pkyanv[64-1]) : 1'b1;


  wire [64-1:0] pqw788qe9_vqac6gylg = 
              ({64{nlb5566a2kkzrak }} & (t3yzmt9i3dp5w7pnh ))
            | ({64{t82iq62ywf1u_5}} & (vkkt61kb_gomf5)) 
            | ({64{byqkkp26xdsszd}} & (vymyvujb_fnw9)) 
            | ({64{vdmyb8x4qmwi7on2 }} & (t3yzmt9i3dp5w7pnh )) 
            | ({64{tfoxw8ia_xdt0}} & (vkkt61kb_gomf5)) 
            | ({64{f128ccj13txxdwpl}} & (vymyvujb_fnw9)); 

  wire p1rgkrlevkumjwua5x = 
              nlb5566a2kkzrak 
            | t82iq62ywf1u_5 
            | byqkkp26xdsszd 
            | vdmyb8x4qmwi7on2  
            | tfoxw8ia_xdt0 
            | f128ccj13txxdwpl; 

  assign bqc9gh1yogik7q5r = 
              ({64{p1rgkrlevkumjwua5x}} & pqw788qe9_vqac6gylg)
            | ({64{nxf52k3xp6im5o6p3}} & {{64-32{1'b1}},nrw_p_xi41_m[31:0]})
            | ({64{gkj8ltdpe4tcqini4h}} & {{64-32{nrw_p_xi41_m[31]}},nrw_p_xi41_m[31:0]}) 
            | ({64{yla1361h}} & {{64-10{1'b0}},tcfrqq029}) 
            | ({64{fp36oxlnph}} & mbi1a[64-1:0])
            | ({64{va7j9_tx3li0xd}} & nrw_p_xi41_m)
            | ({64{tr03xi8fsjspsc}} & nrw_p_xi41_m)
             ;

  assign dd4hyq5oe67rhyvoye = 
              ({5{p1rgkrlevkumjwua5x}} & 5'b0)
            | ({5{nxf52k3xp6im5o6p3}} & 5'b0)
            | ({5{gkj8ltdpe4tcqini4h}} & 5'b0)
            | ({5{tr03xi8fsjspsc}} & 5'b0)
            | ({5{va7j9_tx3li0xd}} & 5'b0)
            | ({5{yla1361h}} & 5'b0) 
            | ({5{fp36oxlnph}} & taferz5nhfy1ttu);


endmodule

module rwxldxdknfy97dlh 
(
  input  [256-1:0] bjh,
  output [8-1:0] ht70 
);

  genvar i;
  wire [256-1:0] i8hem3;
  
  assign i8hem3[256-1]=bjh[256-1];
  
  generate 
  for (i=256-2; i>=0; i=i-1) begin: idcn4vbo1
      assign i8hem3[i] = (|bjh[256-1:i]);
  end
  endgenerate
  
  wire [256-1:0] uhhzbxc = i8hem3 & {1'b1, ~i8hem3[256-1:1]};
  
  assign ht70[0] = 
      |{uhhzbxc[000], uhhzbxc[002], uhhzbxc[004], uhhzbxc[006], uhhzbxc[008],
        uhhzbxc[010], uhhzbxc[012], uhhzbxc[014], uhhzbxc[016], uhhzbxc[018],
        uhhzbxc[020], uhhzbxc[022], uhhzbxc[024], uhhzbxc[026], uhhzbxc[028],
        uhhzbxc[030], uhhzbxc[032], uhhzbxc[034], uhhzbxc[036], uhhzbxc[038],
        uhhzbxc[040], uhhzbxc[042], uhhzbxc[044], uhhzbxc[046], uhhzbxc[048],
        uhhzbxc[050], uhhzbxc[052], uhhzbxc[054], uhhzbxc[056], uhhzbxc[058],
        uhhzbxc[060], uhhzbxc[062], uhhzbxc[064], uhhzbxc[066], uhhzbxc[068],
        uhhzbxc[070], uhhzbxc[072], uhhzbxc[074], uhhzbxc[076], uhhzbxc[078],
        uhhzbxc[080], uhhzbxc[082], uhhzbxc[084], uhhzbxc[086], uhhzbxc[088],
        uhhzbxc[090], uhhzbxc[092], uhhzbxc[094], uhhzbxc[096], uhhzbxc[098],
        uhhzbxc[100], uhhzbxc[102], uhhzbxc[104], uhhzbxc[106], uhhzbxc[108],
        uhhzbxc[110], uhhzbxc[112], uhhzbxc[114], uhhzbxc[116], uhhzbxc[118],
        uhhzbxc[120], uhhzbxc[122], uhhzbxc[124], uhhzbxc[126], uhhzbxc[128],
        uhhzbxc[130], uhhzbxc[132], uhhzbxc[134], uhhzbxc[136], uhhzbxc[138],
        uhhzbxc[140], uhhzbxc[142], uhhzbxc[144], uhhzbxc[146], uhhzbxc[148],
        uhhzbxc[150], uhhzbxc[152], uhhzbxc[154], uhhzbxc[156], uhhzbxc[158],
        uhhzbxc[160], uhhzbxc[162], uhhzbxc[164], uhhzbxc[166], uhhzbxc[168],
        uhhzbxc[170], uhhzbxc[172], uhhzbxc[174], uhhzbxc[176], uhhzbxc[178],
        uhhzbxc[180], uhhzbxc[182], uhhzbxc[184], uhhzbxc[186], uhhzbxc[188],
        uhhzbxc[190], uhhzbxc[192], uhhzbxc[194], uhhzbxc[196], uhhzbxc[198],
        uhhzbxc[200], uhhzbxc[202], uhhzbxc[204], uhhzbxc[206], uhhzbxc[208],
        uhhzbxc[210], uhhzbxc[212], uhhzbxc[214], uhhzbxc[216], uhhzbxc[218],
        uhhzbxc[220], uhhzbxc[222], uhhzbxc[224], uhhzbxc[226], uhhzbxc[228],
        uhhzbxc[230], uhhzbxc[232], uhhzbxc[234], uhhzbxc[236], uhhzbxc[238],
        uhhzbxc[240], uhhzbxc[242], uhhzbxc[244], uhhzbxc[246], uhhzbxc[248],
        uhhzbxc[250], uhhzbxc[252], uhhzbxc[254]};
  
  assign ht70[1] = 
      |{uhhzbxc[000], uhhzbxc[001], uhhzbxc[004], uhhzbxc[005], 
        uhhzbxc[008], uhhzbxc[009], uhhzbxc[012], uhhzbxc[013], 
        uhhzbxc[016], uhhzbxc[017], uhhzbxc[020], uhhzbxc[021], 
        uhhzbxc[024], uhhzbxc[025], uhhzbxc[028], uhhzbxc[029], 
        uhhzbxc[032], uhhzbxc[033], uhhzbxc[036], uhhzbxc[037],
        uhhzbxc[040], uhhzbxc[041], uhhzbxc[044], uhhzbxc[045], 
        uhhzbxc[048], uhhzbxc[049], uhhzbxc[052], uhhzbxc[053], 
        uhhzbxc[056], uhhzbxc[057], uhhzbxc[060], uhhzbxc[061],
        uhhzbxc[064], uhhzbxc[065], uhhzbxc[068], uhhzbxc[069], 
        uhhzbxc[072], uhhzbxc[073], uhhzbxc[076], uhhzbxc[077],
        uhhzbxc[080], uhhzbxc[081], uhhzbxc[084], uhhzbxc[085], 
        uhhzbxc[088], uhhzbxc[089], uhhzbxc[092], uhhzbxc[093], 
        uhhzbxc[096], uhhzbxc[097], uhhzbxc[100], uhhzbxc[101],
        uhhzbxc[104], uhhzbxc[105], uhhzbxc[108], uhhzbxc[109], 
        uhhzbxc[112], uhhzbxc[113], uhhzbxc[116], uhhzbxc[117],
        uhhzbxc[120], uhhzbxc[121], uhhzbxc[124], uhhzbxc[125],
        uhhzbxc[128], uhhzbxc[129], uhhzbxc[132], uhhzbxc[133],
        uhhzbxc[136], uhhzbxc[137], uhhzbxc[140], uhhzbxc[141],
        uhhzbxc[144], uhhzbxc[145], uhhzbxc[148], uhhzbxc[149],
        uhhzbxc[152], uhhzbxc[153], uhhzbxc[156], uhhzbxc[157],
        uhhzbxc[160], uhhzbxc[161], uhhzbxc[164], uhhzbxc[165],
        uhhzbxc[168], uhhzbxc[169], uhhzbxc[172], uhhzbxc[173],
        uhhzbxc[176], uhhzbxc[177], uhhzbxc[180], uhhzbxc[181],
        uhhzbxc[184], uhhzbxc[185], uhhzbxc[188], uhhzbxc[189],
        uhhzbxc[192], uhhzbxc[193], uhhzbxc[196], uhhzbxc[197],
        uhhzbxc[200], uhhzbxc[201], uhhzbxc[204], uhhzbxc[205],
        uhhzbxc[208], uhhzbxc[209], uhhzbxc[212], uhhzbxc[213],
        uhhzbxc[216], uhhzbxc[217], uhhzbxc[220], uhhzbxc[221],
        uhhzbxc[224], uhhzbxc[225], uhhzbxc[228], uhhzbxc[229],
        uhhzbxc[232], uhhzbxc[233], uhhzbxc[236], uhhzbxc[237],
        uhhzbxc[240], uhhzbxc[241], uhhzbxc[244], uhhzbxc[245],
        uhhzbxc[248], uhhzbxc[249], uhhzbxc[252], uhhzbxc[253]};
  
  assign ht70[2] =
      |{uhhzbxc[000], uhhzbxc[001], uhhzbxc[002], uhhzbxc[003], 
        uhhzbxc[008], uhhzbxc[009], uhhzbxc[010], uhhzbxc[011], 
        uhhzbxc[016], uhhzbxc[017], uhhzbxc[018], uhhzbxc[019], 
        uhhzbxc[024], uhhzbxc[025], uhhzbxc[026], uhhzbxc[027], 
        uhhzbxc[032], uhhzbxc[033], uhhzbxc[034], uhhzbxc[035],
        uhhzbxc[040], uhhzbxc[041], uhhzbxc[042], uhhzbxc[043], 
        uhhzbxc[048], uhhzbxc[049], uhhzbxc[050], uhhzbxc[051], 
        uhhzbxc[056], uhhzbxc[057], uhhzbxc[058], uhhzbxc[059],
        uhhzbxc[064], uhhzbxc[065], uhhzbxc[066], uhhzbxc[067], 
        uhhzbxc[072], uhhzbxc[073], uhhzbxc[074], uhhzbxc[075],
        uhhzbxc[080], uhhzbxc[081], uhhzbxc[082], uhhzbxc[083], 
        uhhzbxc[088], uhhzbxc[089], uhhzbxc[090], uhhzbxc[091], 
        uhhzbxc[096], uhhzbxc[097], uhhzbxc[098], uhhzbxc[099],
        uhhzbxc[104], uhhzbxc[105], uhhzbxc[106], uhhzbxc[107], 
        uhhzbxc[112], uhhzbxc[113], uhhzbxc[114], uhhzbxc[115],
        uhhzbxc[120], uhhzbxc[121], uhhzbxc[122], uhhzbxc[123],
        uhhzbxc[128], uhhzbxc[129], uhhzbxc[130], uhhzbxc[131],
        uhhzbxc[136], uhhzbxc[137], uhhzbxc[138], uhhzbxc[139],
        uhhzbxc[144], uhhzbxc[145], uhhzbxc[146], uhhzbxc[147],
        uhhzbxc[152], uhhzbxc[153], uhhzbxc[154], uhhzbxc[155],
        uhhzbxc[160], uhhzbxc[161], uhhzbxc[162], uhhzbxc[163],
        uhhzbxc[168], uhhzbxc[169], uhhzbxc[170], uhhzbxc[171],
        uhhzbxc[176], uhhzbxc[177], uhhzbxc[178], uhhzbxc[179],
        uhhzbxc[184], uhhzbxc[185], uhhzbxc[186], uhhzbxc[187],
        uhhzbxc[192], uhhzbxc[193], uhhzbxc[194], uhhzbxc[195],
        uhhzbxc[200], uhhzbxc[201], uhhzbxc[202], uhhzbxc[203],
        uhhzbxc[208], uhhzbxc[209], uhhzbxc[210], uhhzbxc[211],
        uhhzbxc[216], uhhzbxc[217], uhhzbxc[218], uhhzbxc[219],
        uhhzbxc[224], uhhzbxc[225], uhhzbxc[226], uhhzbxc[227],
        uhhzbxc[232], uhhzbxc[233], uhhzbxc[234], uhhzbxc[235],
        uhhzbxc[240], uhhzbxc[241], uhhzbxc[242], uhhzbxc[243],
        uhhzbxc[248], uhhzbxc[249], uhhzbxc[250], uhhzbxc[251]};
  
  assign ht70[3] =
      |{uhhzbxc[000], uhhzbxc[001], uhhzbxc[002], uhhzbxc[003], uhhzbxc[004], uhhzbxc[005], uhhzbxc[006], uhhzbxc[007], 
        uhhzbxc[016], uhhzbxc[017], uhhzbxc[018], uhhzbxc[019], uhhzbxc[020], uhhzbxc[021], uhhzbxc[022], uhhzbxc[023], 
        uhhzbxc[032], uhhzbxc[033], uhhzbxc[034], uhhzbxc[035], uhhzbxc[036], uhhzbxc[037], uhhzbxc[038], uhhzbxc[039], 
        uhhzbxc[048], uhhzbxc[049], uhhzbxc[050], uhhzbxc[051], uhhzbxc[052], uhhzbxc[053], uhhzbxc[054], uhhzbxc[055],
        uhhzbxc[064], uhhzbxc[065], uhhzbxc[066], uhhzbxc[067], uhhzbxc[068], uhhzbxc[069], uhhzbxc[070], uhhzbxc[071],
        uhhzbxc[080], uhhzbxc[081], uhhzbxc[082], uhhzbxc[083], uhhzbxc[084], uhhzbxc[085], uhhzbxc[086], uhhzbxc[087], 
        uhhzbxc[096], uhhzbxc[097], uhhzbxc[098], uhhzbxc[099], uhhzbxc[100], uhhzbxc[101], uhhzbxc[102], uhhzbxc[103], 
        uhhzbxc[112], uhhzbxc[113], uhhzbxc[114], uhhzbxc[115], uhhzbxc[116], uhhzbxc[117], uhhzbxc[118], uhhzbxc[119],
        uhhzbxc[128], uhhzbxc[129], uhhzbxc[130], uhhzbxc[131], uhhzbxc[132], uhhzbxc[133], uhhzbxc[134], uhhzbxc[135],
        uhhzbxc[144], uhhzbxc[145], uhhzbxc[146], uhhzbxc[147], uhhzbxc[148], uhhzbxc[149], uhhzbxc[150], uhhzbxc[151],
        uhhzbxc[160], uhhzbxc[161], uhhzbxc[162], uhhzbxc[163], uhhzbxc[164], uhhzbxc[165], uhhzbxc[166], uhhzbxc[167],
        uhhzbxc[176], uhhzbxc[177], uhhzbxc[178], uhhzbxc[179], uhhzbxc[180], uhhzbxc[181], uhhzbxc[182], uhhzbxc[183],
        uhhzbxc[192], uhhzbxc[193], uhhzbxc[194], uhhzbxc[195], uhhzbxc[196], uhhzbxc[197], uhhzbxc[198], uhhzbxc[199],
        uhhzbxc[208], uhhzbxc[209], uhhzbxc[210], uhhzbxc[211], uhhzbxc[212], uhhzbxc[213], uhhzbxc[214], uhhzbxc[215],
        uhhzbxc[224], uhhzbxc[225], uhhzbxc[226], uhhzbxc[227], uhhzbxc[228], uhhzbxc[229], uhhzbxc[230], uhhzbxc[231],
        uhhzbxc[240], uhhzbxc[241], uhhzbxc[242], uhhzbxc[243], uhhzbxc[244], uhhzbxc[245], uhhzbxc[246], uhhzbxc[247]};
  
  assign ht70[4] = 
      |{uhhzbxc[000], uhhzbxc[001], uhhzbxc[002], uhhzbxc[003], uhhzbxc[004], uhhzbxc[005], uhhzbxc[006], uhhzbxc[007], uhhzbxc[008], uhhzbxc[009], uhhzbxc[010], uhhzbxc[011], uhhzbxc[012], uhhzbxc[013], uhhzbxc[014], uhhzbxc[015], 
        uhhzbxc[032], uhhzbxc[033], uhhzbxc[034], uhhzbxc[035], uhhzbxc[036], uhhzbxc[037], uhhzbxc[038], uhhzbxc[039], uhhzbxc[040], uhhzbxc[041], uhhzbxc[042], uhhzbxc[043], uhhzbxc[044], uhhzbxc[045], uhhzbxc[046], uhhzbxc[047], 
        uhhzbxc[064], uhhzbxc[065], uhhzbxc[066], uhhzbxc[067], uhhzbxc[068], uhhzbxc[069], uhhzbxc[070], uhhzbxc[071], uhhzbxc[072], uhhzbxc[073], uhhzbxc[074], uhhzbxc[075], uhhzbxc[076], uhhzbxc[077], uhhzbxc[078], uhhzbxc[079],
        uhhzbxc[096], uhhzbxc[097], uhhzbxc[098], uhhzbxc[099], uhhzbxc[100], uhhzbxc[101], uhhzbxc[102], uhhzbxc[103], uhhzbxc[104], uhhzbxc[105], uhhzbxc[106], uhhzbxc[107], uhhzbxc[108], uhhzbxc[109], uhhzbxc[110], uhhzbxc[111],
        uhhzbxc[128], uhhzbxc[129], uhhzbxc[130], uhhzbxc[131], uhhzbxc[132], uhhzbxc[133], uhhzbxc[134], uhhzbxc[135], uhhzbxc[136], uhhzbxc[137], uhhzbxc[138], uhhzbxc[139], uhhzbxc[140], uhhzbxc[141], uhhzbxc[142], uhhzbxc[143],
        uhhzbxc[160], uhhzbxc[161], uhhzbxc[162], uhhzbxc[163], uhhzbxc[164], uhhzbxc[165], uhhzbxc[166], uhhzbxc[167], uhhzbxc[168], uhhzbxc[169], uhhzbxc[170], uhhzbxc[171], uhhzbxc[172], uhhzbxc[173], uhhzbxc[174], uhhzbxc[175],
        uhhzbxc[192], uhhzbxc[193], uhhzbxc[194], uhhzbxc[195], uhhzbxc[196], uhhzbxc[197], uhhzbxc[198], uhhzbxc[199], uhhzbxc[200], uhhzbxc[201], uhhzbxc[202], uhhzbxc[203], uhhzbxc[204], uhhzbxc[205], uhhzbxc[206], uhhzbxc[207],
        uhhzbxc[224], uhhzbxc[225], uhhzbxc[226], uhhzbxc[227], uhhzbxc[228], uhhzbxc[229], uhhzbxc[230], uhhzbxc[231], uhhzbxc[232], uhhzbxc[233], uhhzbxc[234], uhhzbxc[235], uhhzbxc[236], uhhzbxc[237], uhhzbxc[238], uhhzbxc[239]};
  
  assign ht70[5] =
      |{uhhzbxc[000], uhhzbxc[001], uhhzbxc[002], uhhzbxc[003], uhhzbxc[004], uhhzbxc[005], uhhzbxc[006], uhhzbxc[007], uhhzbxc[008], uhhzbxc[009], uhhzbxc[010], uhhzbxc[011], uhhzbxc[012], uhhzbxc[013], uhhzbxc[014], uhhzbxc[015], 
        uhhzbxc[016], uhhzbxc[017], uhhzbxc[018], uhhzbxc[019], uhhzbxc[020], uhhzbxc[021], uhhzbxc[022], uhhzbxc[023], uhhzbxc[024], uhhzbxc[025], uhhzbxc[026], uhhzbxc[027], uhhzbxc[028], uhhzbxc[029], uhhzbxc[030], uhhzbxc[031],
        uhhzbxc[064], uhhzbxc[065], uhhzbxc[066], uhhzbxc[067], uhhzbxc[068], uhhzbxc[069], uhhzbxc[070], uhhzbxc[071], uhhzbxc[072], uhhzbxc[073], uhhzbxc[074], uhhzbxc[075], uhhzbxc[076], uhhzbxc[077], uhhzbxc[078], uhhzbxc[079],
        uhhzbxc[080], uhhzbxc[081], uhhzbxc[082], uhhzbxc[083], uhhzbxc[084], uhhzbxc[085], uhhzbxc[086], uhhzbxc[087], uhhzbxc[088], uhhzbxc[089], uhhzbxc[090], uhhzbxc[091], uhhzbxc[092], uhhzbxc[093], uhhzbxc[094], uhhzbxc[095],
        uhhzbxc[128], uhhzbxc[129], uhhzbxc[130], uhhzbxc[131], uhhzbxc[132], uhhzbxc[133], uhhzbxc[134], uhhzbxc[135], uhhzbxc[136], uhhzbxc[137], uhhzbxc[138], uhhzbxc[139], uhhzbxc[140], uhhzbxc[141], uhhzbxc[142], uhhzbxc[143],
        uhhzbxc[144], uhhzbxc[145], uhhzbxc[146], uhhzbxc[147], uhhzbxc[148], uhhzbxc[149], uhhzbxc[150], uhhzbxc[151], uhhzbxc[152], uhhzbxc[153], uhhzbxc[154], uhhzbxc[155], uhhzbxc[156], uhhzbxc[157], uhhzbxc[158], uhhzbxc[159], 
        uhhzbxc[192], uhhzbxc[193], uhhzbxc[194], uhhzbxc[195], uhhzbxc[196], uhhzbxc[197], uhhzbxc[198], uhhzbxc[199], uhhzbxc[200], uhhzbxc[201], uhhzbxc[202], uhhzbxc[203], uhhzbxc[204], uhhzbxc[205], uhhzbxc[206], uhhzbxc[207],
        uhhzbxc[208], uhhzbxc[209], uhhzbxc[210], uhhzbxc[211], uhhzbxc[212], uhhzbxc[213], uhhzbxc[214], uhhzbxc[215], uhhzbxc[216], uhhzbxc[217], uhhzbxc[218], uhhzbxc[219], uhhzbxc[220], uhhzbxc[221], uhhzbxc[222], uhhzbxc[223]};
  
  assign ht70[6] =
      |{uhhzbxc[000], uhhzbxc[001], uhhzbxc[002], uhhzbxc[003], uhhzbxc[004], uhhzbxc[005], uhhzbxc[006], uhhzbxc[007], uhhzbxc[008], uhhzbxc[009], uhhzbxc[010], uhhzbxc[011], uhhzbxc[012], uhhzbxc[013], uhhzbxc[014], uhhzbxc[015], 
        uhhzbxc[016], uhhzbxc[017], uhhzbxc[018], uhhzbxc[019], uhhzbxc[020], uhhzbxc[021], uhhzbxc[022], uhhzbxc[023], uhhzbxc[024], uhhzbxc[025], uhhzbxc[026], uhhzbxc[027], uhhzbxc[028], uhhzbxc[029], uhhzbxc[030], uhhzbxc[031],
        uhhzbxc[032], uhhzbxc[033], uhhzbxc[034], uhhzbxc[035], uhhzbxc[036], uhhzbxc[037], uhhzbxc[038], uhhzbxc[039], uhhzbxc[040], uhhzbxc[041], uhhzbxc[042], uhhzbxc[043], uhhzbxc[044], uhhzbxc[045], uhhzbxc[046], uhhzbxc[047], 
        uhhzbxc[048], uhhzbxc[049], uhhzbxc[050], uhhzbxc[051], uhhzbxc[052], uhhzbxc[053], uhhzbxc[054], uhhzbxc[055], uhhzbxc[056], uhhzbxc[057], uhhzbxc[058], uhhzbxc[059], uhhzbxc[060], uhhzbxc[061], uhhzbxc[062], uhhzbxc[063],
        uhhzbxc[128], uhhzbxc[129], uhhzbxc[130], uhhzbxc[131], uhhzbxc[132], uhhzbxc[133], uhhzbxc[134], uhhzbxc[135], uhhzbxc[136], uhhzbxc[137], uhhzbxc[138], uhhzbxc[139], uhhzbxc[140], uhhzbxc[141], uhhzbxc[142], uhhzbxc[143],
        uhhzbxc[144], uhhzbxc[145], uhhzbxc[146], uhhzbxc[147], uhhzbxc[148], uhhzbxc[149], uhhzbxc[150], uhhzbxc[151], uhhzbxc[152], uhhzbxc[153], uhhzbxc[154], uhhzbxc[155], uhhzbxc[156], uhhzbxc[157], uhhzbxc[158], uhhzbxc[159],
        uhhzbxc[160], uhhzbxc[161], uhhzbxc[162], uhhzbxc[163], uhhzbxc[164], uhhzbxc[165], uhhzbxc[166], uhhzbxc[167], uhhzbxc[168], uhhzbxc[169], uhhzbxc[170], uhhzbxc[171], uhhzbxc[172], uhhzbxc[173], uhhzbxc[174], uhhzbxc[175],
        uhhzbxc[176], uhhzbxc[177], uhhzbxc[178], uhhzbxc[179], uhhzbxc[180], uhhzbxc[181], uhhzbxc[182], uhhzbxc[183], uhhzbxc[184], uhhzbxc[185], uhhzbxc[186], uhhzbxc[187], uhhzbxc[188], uhhzbxc[189], uhhzbxc[190], uhhzbxc[191]};
  
  assign ht70[7]=
      |{uhhzbxc[000], uhhzbxc[001], uhhzbxc[002], uhhzbxc[003], uhhzbxc[004], uhhzbxc[005], uhhzbxc[006], uhhzbxc[007], uhhzbxc[008], uhhzbxc[009], uhhzbxc[010], uhhzbxc[011], uhhzbxc[012], uhhzbxc[013], uhhzbxc[014], uhhzbxc[015], 
        uhhzbxc[016], uhhzbxc[017], uhhzbxc[018], uhhzbxc[019], uhhzbxc[020], uhhzbxc[021], uhhzbxc[022], uhhzbxc[023], uhhzbxc[024], uhhzbxc[025], uhhzbxc[026], uhhzbxc[027], uhhzbxc[028], uhhzbxc[029], uhhzbxc[030], uhhzbxc[031],
        uhhzbxc[032], uhhzbxc[033], uhhzbxc[034], uhhzbxc[035], uhhzbxc[036], uhhzbxc[037], uhhzbxc[038], uhhzbxc[039], uhhzbxc[040], uhhzbxc[041], uhhzbxc[042], uhhzbxc[043], uhhzbxc[044], uhhzbxc[045], uhhzbxc[046], uhhzbxc[047], 
        uhhzbxc[048], uhhzbxc[049], uhhzbxc[050], uhhzbxc[051], uhhzbxc[052], uhhzbxc[053], uhhzbxc[054], uhhzbxc[055], uhhzbxc[056], uhhzbxc[057], uhhzbxc[058], uhhzbxc[059], uhhzbxc[060], uhhzbxc[061], uhhzbxc[062], uhhzbxc[063],
        uhhzbxc[064], uhhzbxc[065], uhhzbxc[066], uhhzbxc[067], uhhzbxc[068], uhhzbxc[069], uhhzbxc[070], uhhzbxc[071], uhhzbxc[072], uhhzbxc[073], uhhzbxc[074], uhhzbxc[075], uhhzbxc[076], uhhzbxc[077], uhhzbxc[078], uhhzbxc[079],
        uhhzbxc[080], uhhzbxc[081], uhhzbxc[082], uhhzbxc[083], uhhzbxc[084], uhhzbxc[085], uhhzbxc[086], uhhzbxc[087], uhhzbxc[088], uhhzbxc[089], uhhzbxc[090], uhhzbxc[091], uhhzbxc[092], uhhzbxc[093], uhhzbxc[094], uhhzbxc[095],
        uhhzbxc[096], uhhzbxc[097], uhhzbxc[098], uhhzbxc[099], uhhzbxc[100], uhhzbxc[101], uhhzbxc[102], uhhzbxc[103], uhhzbxc[104], uhhzbxc[105], uhhzbxc[106], uhhzbxc[107], uhhzbxc[108], uhhzbxc[109], uhhzbxc[110], uhhzbxc[111],
        uhhzbxc[112], uhhzbxc[113], uhhzbxc[114], uhhzbxc[115], uhhzbxc[116], uhhzbxc[117], uhhzbxc[118], uhhzbxc[119], uhhzbxc[120], uhhzbxc[121], uhhzbxc[122], uhhzbxc[123], uhhzbxc[124], uhhzbxc[125], uhhzbxc[126], uhhzbxc[127]}; 

endmodule

module wjr2um7_i8ekzqst54wvn1f0 #(
    parameter onr7l = 1,
    parameter ap4sz86dvorgz = 0
)(
  input               abwn, 
  input      [onr7l-1:0] q461tw,
  output     [onr7l-1:0] p4dxkq4k,

  input               gf33atgy ,
  input               ru_wi
);

genvar i;
generate 
if(ap4sz86dvorgz==1) begin:budlxvga9h401opfwvo1rx

reg [onr7l-1:0] nkvgr6w73w;

always @(posedge gf33atgy or negedge ru_wi)
begin : nz_z_r5hu30j
  if (ru_wi == 1'b0)
    nkvgr6w73w <= {onr7l{1'b0}};
  else if (abwn == 1'b1)
    nkvgr6w73w <= q461tw;
end

assign p4dxkq4k = nkvgr6w73w;


end
else begin:z9p6qiexnudiymcatx6l
    assign p4dxkq4k = q461tw;
end

endgenerate
endmodule 


















module dv_v4v1au7ht_i2qt(
  input  [5-1:0] w42_wd9um28vh,
  input  [5-1:0] ssjx8h5cj3q4ffem,
  input  [5-1:0] rwby8vkzgm4y4r,
  output [64-1:0] vuv0917fanv19,
  output [64-1:0] j2xzlc7dmxgmtn6kmk,
  output [64-1:0] tkxnzh2vh65vfutt3,

  input  qd7ilyg140avze,
  input  [5-1:0] n9uum984u41is66h2f,
  input  [64-1:0] kf_pg4o0m8fa8,

  input  gc4b3kdcan6do88ta_,
  input  gf33atgy,
  input  ru_wi
  );

  wire [64-1:0] fbu76k [32-1:0];
  wire [32-1:0] leab8mqf;
  

  
  genvar i;
  generate 
  
      for (i=0; i<32; i=i+1) begin:ubs_7gmy192w
  
        
        
        
        
        
        
        
        
        
        
            assign leab8mqf[i] = qd7ilyg140avze & (n9uum984u41is66h2f == i[5-1:0]) ;
            ux607_gnrl_dfflr #(64) ddzbam3h39f (leab8mqf[i], kf_pg4o0m8fa8, fbu76k[i], gf33atgy, ru_wi);
        
  
      end
  endgenerate
  
  assign vuv0917fanv19 = fbu76k[w42_wd9um28vh];
  assign j2xzlc7dmxgmtn6kmk = fbu76k[ssjx8h5cj3q4ffem];
  assign tkxnzh2vh65vfutt3 = fbu76k[rwby8vkzgm4y4r];
  
endmodule



















module s6iu1fy58ac1rlrw4s8v (
    input  [31:0] v2aj2jo,
    input  dwnd9ctj5,

    output [15:0] uiwlxd,
    output [4:0] adnx9wgdt2

);

  
   wire [3-1:0] vc529nuu = 3'b001; 

   wire v0da13u6ykrw = (v2aj2jo[30:23] == 8'hFF);
   wire rg17tsy6wwx = (v2aj2jo[30:23] == 8'h00);
   wire wb75liyzd6vmew7 = (v2aj2jo[22:0] == 23'b0);
   wire bml43dgqbvm = rg17tsy6wwx & (~wb75liyzd6vmew7);
   wire ib3hkx1k0t = v2aj2jo[22];
   wire mgvwdehh1 = (~v0da13u6ykrw) & (~rg17tsy6wwx);
   wire aswm0l3tr55 = v0da13u6ykrw & (~wb75liyzd6vmew7) & (~ib3hkx1k0t);
   wire r41nzg = v0da13u6ykrw & (~wb75liyzd6vmew7) & ib3hkx1k0t;
   wire jqgto = r41nzg | aswm0l3tr55;
   wire ak6syfq = v0da13u6ykrw & wb75liyzd6vmew7;
   wire sy1qjmixh5e = (rg17tsy6wwx & wb75liyzd6vmew7);

   wire [22:0]  lkish79hpt = v2aj2jo[22:0];
   wire [ 7:0]  dbw_bap_jqyl = v2aj2jo[30:23];
   wire         a8rijdb567ulj = v2aj2jo[31];


   wire [22:0]  d86mct = lkish79hpt;
   wire         mp3k_c3d = a8rijdb567ulj;
   wire [ 7:0]  eff76eu5r  = dbw_bap_jqyl;

   wire [23:0]  xf92vp2m3d = {mgvwdehh1, d86mct};                       

   wire zpwosdnwv0 = ak6syfq & (~mp3k_c3d);
   wire h2pw9rtks0i = ak6syfq & mp3k_c3d;

   wire eqi5fiol = sy1qjmixh5e & (~mp3k_c3d);
   wire kc2obnf0fo = sy1qjmixh5e & mp3k_c3d;

   wire [32-1:0] e5otgqgjkm78gyd   = 32'h7FC00000;
   wire [16-1:0] rphhy7og5shc   = 16'h7E00;
   wire [32-1:0] lkpuz8x2a1y5   = 32'h7F800000;
   wire [16-1:0] wztskukp1m94m   = 16'h7C00;
   wire [32-1:0] w4m58zc6vxjqm   = 32'hFF800000;
   wire [16-1:0] os3en__39s   = 16'hFC00;
   wire [32-1:0] ppp30tohtvbsq   = 32'h00000000;
   wire [32-1:0] l2mifwazi5t_   = 32'h80000000;
   wire [16-1:0] c89mpiadrlqqb   = 16'h0000;
   wire [16-1:0] ged2mj90blbvit   = 16'h8000;
   wire [16-1:0] gz6qduuihnykm = 16'h7BFF;
   wire [16-1:0] s1th5gccdkngj = 16'hFBFF;



















   wire [7:0]  mx2koejh0gysa;
   wire [7:0]  uo3bnxjifojicun;
   wire  giyoqem5ltdmbn4ny_1f;
   wire  bxof3bheoo0ndkjymw;
   assign {giyoqem5ltdmbn4ny_1f,mx2koejh0gysa} = {1'b0,dbw_bap_jqyl} + (~(9'd112)) + 1'b1;
   assign {bxof3bheoo0ndkjymw,uo3bnxjifojicun} = 9'd112 + (~{1'b0,dbw_bap_jqyl}) + 1'b1; 
 
   
   wire qj8e_p7rnbges5rxdwo= (&mx2koejh0gysa[4:0]);
   wire rzf556ieod2ogdok0xlq4= ~(|mx2koejh0gysa[4:0]);
   wire nhkrkbqafcs3pe02ip6f = (~giyoqem5ltdmbn4ny_1f) & ((|mx2koejh0gysa[7:5]) | qj8e_p7rnbges5rxdwo); 
   wire b4tobe5ck4dt68fysscsx = giyoqem5ltdmbn4ny_1f & (|uo3bnxjifojicun[7:4]);
 
   wire ao5qzutvei2pnx = (~giyoqem5ltdmbn4ny_1f) & (~(|mx2koejh0gysa[7:5])) & (~qj8e_p7rnbges5rxdwo) & (~rzf556ieod2ogdok0xlq4);
 
   wire lcq6dingl_mwz2876vd4 = (~(nhkrkbqafcs3pe02ip6f | b4tobe5ck4dt68fysscsx | ao5qzutvei2pnx));
   wire kmcrpnpwy7cgu5iycx   = (~giyoqem5ltdmbn4ny_1f) & (mx2koejh0gysa == 8'd0);

   wire jyi_fwis89t7cyz3a;
   wire [10:0] t34p1fwqw_9vwel;
   wire ke78qjh44u_yl9we;
   wire pcng4dtn_do4tx;
   wire [27:0] p_9df234l2l5wj2i04zr;
   wire ghy7mapy6qzp1zk5sjh = |p_9df234l2l5wj2i04zr;

   
   
   
   wire omaxte58qmuedb = 
               ((vc529nuu == 3'b000) & 1'b1) 
              |((vc529nuu == 3'b011) & (~a8rijdb567ulj)) 
              |((vc529nuu == 3'b010) & a8rijdb567ulj)
              |((vc529nuu == 3'b001) & 1'b0)         
              |((vc529nuu == 3'b100) & 1'b1);

   wire txiyqjrxqklqzoc = |xf92vp2m3d;

   wire [40:0] rjuh2vh4d1gfvl = ({xf92vp2m3d[23:0],17'b0} >>  uo3bnxjifojicun[3:0]);

   assign {t34p1fwqw_9vwel, ke78qjh44u_yl9we, pcng4dtn_do4tx, p_9df234l2l5wj2i04zr} =
                       
                 b4tobe5ck4dt68fysscsx ? {11'b0, 1'b0, 1'b0, txiyqjrxqklqzoc, 27'b0 }: 
                       

                 (nhkrkbqafcs3pe02ip6f & (~omaxte58qmuedb)) ? {(~11'b0), 1'b0, 1'b0, 1'b0, 27'b0} :
                       
                 ao5qzutvei2pnx ? {xf92vp2m3d[23:0], 17'b0} :
                       
                       
                 (rjuh2vh4d1gfvl >> 1'b1);

  assign jyi_fwis89t7cyz3a = 1'b0;  
  wire [22:0] uyf04u627pz9335y = t34p1fwqw_9vwel + jyi_fwis89t7cyz3a;   

  wire ewwgdb6evrflrp0 = 1'b0; 

  wire [ 9:0] mwlhwtvo = ewwgdb6evrflrp0 ? 10'b0 : uyf04u627pz9335y[9:0];

  wire [ 4:0] vgibybipl6i = 
                       
                 b4tobe5ck4dt68fysscsx ? 5'b0 :
                       

                 (nhkrkbqafcs3pe02ip6f & (~omaxte58qmuedb)) ? 5'h1E : 
                       
                       
                 ao5qzutvei2pnx ? (ewwgdb6evrflrp0 ? (mx2koejh0gysa[4:0] + 1'b1) : mx2koejh0gysa[4:0]) :
                       
                 5'h0;

  wire pzolaxcukx08n6d88qz88axk8g = 1'b0;  

  wire [15:0] gyn7zbs8py =
  
                     
                 jqgto   ? rphhy7og5shc :
                     
                 zpwosdnwv0 ? wztskukp1m94m :
                 h2pw9rtks0i ? os3en__39s :
                     
                 eqi5fiol ? c89mpiadrlqqb :
                 kc2obnf0fo ? ged2mj90blbvit : {mp3k_c3d,vgibybipl6i[4:0],mwlhwtvo};

   wire qdsazoqaefdqv0vl9ejx11 = (jqgto | zpwosdnwv0 | h2pw9rtks0i | eqi5fiol | kc2obnf0fo);
   
   
   
   
   wire iuyfqp38m0h3ebb2bv = aswm0l3tr55;
   
   wire ecarjrbm5vjgzgez0 = 1'b0;
   
   
   wire d73m4m2luplwqf = (~qdsazoqaefdqv0vl9ejx11) & (b4tobe5ck4dt68fysscsx | lcq6dingl_mwz2876vd4) 
                          & (ke78qjh44u_yl9we | pcng4dtn_do4tx | ghy7mapy6qzp1zk5sjh);
   
        
   wire jf1dnyje2gl6x = (~qdsazoqaefdqv0vl9ejx11) & (nhkrkbqafcs3pe02ip6f | pzolaxcukx08n6d88qz88axk8g);
   
   wire op9apkpdawjzjnkb = (~qdsazoqaefdqv0vl9ejx11) & (ke78qjh44u_yl9we | pcng4dtn_do4tx | ghy7mapy6qzp1zk5sjh | d73m4m2luplwqf | jf1dnyje2gl6x);

   wire [4:0] vwypdfhpqweqgb9yxjk = {op9apkpdawjzjnkb, d73m4m2luplwqf, jf1dnyje2gl6x, ecarjrbm5vjgzgez0, iuyfqp38m0h3ebb2bv};







  assign uiwlxd = {16{dwnd9ctj5}} & gyn7zbs8py;

  wire [4:0] k6mvi11sj = ({5{dwnd9ctj5}} & vwypdfhpqweqgb9yxjk);

  assign adnx9wgdt2 = {k6mvi11sj[0],k6mvi11sj[1],k6mvi11sj[2],k6mvi11sj[3],k6mvi11sj[4]}; 

endmodule























module re1ncz9e2e3zo(















 
  input  [48-1:0] k9lv9ppimt14qx3d7rj,  
  input  [64-1:0] llskuqv0ehm60atlo,
  input  oug11blpzcta8zyu0ya,
  input  zr1pc8tfxyljdj7a8a3eh5,
  input  qg9g70jgx5r5l_wpc7,
  input  o_qquv0pnx4zpz4h3gwxgl3,
  input  j1fek3jzmt5bhhpnhvrmgt,
  input  ds75nafgmrespy002qvcsb8,

  input                           rclkn1q60a3cbgtn67g,
  input [48-1:0] zamt9z8_hsjwlky8aktxv6,  
  input [64-1:0]          ofmr0b7vez483r8wl ,
  input [64-1:0]          zgn_d2n28xfn1zff ,
  input [64-1:0]          ceewyf1unn6p7peejem ,
  input [64-1:0]          oegl6jlhw01xkqeetu5y ,



  input [5-1:0] ehq614orwiy4ww5,
  input [5-1:0] hgg2w2ca4wsixuj,
  input [5-1:0] lgv405vv46,
  output [64-1:0] vwxjizbv8c62_r6sf,
  output [64-1:0] ft8qpl2cvbar7ci,
  output [64-1:0] fi80hkldjwlh4v,





  
  
  input  dkmuhc79d2wm0wubp, 
  input  u2demhkod_er3kf6b, 
  output uz7pt71lvqit85od, 
  input  [4-1:0] v3uvhtx7e5vbtvie,
  input  [3-1:0] l60zv02z95hlayri,
  output l1xzyldaa9dr2q7mla,
  input  [64-1:0] tmqkgmlzi018,
  input  [64-1:0] lx_olubu7t8h,
  input  [64-1:0] dd1p3tnenmm9r,

  
  
  
  output a5z_23_ryr_m29hhia_p      ,
  
 
  input  vejdvgqormu727s,
  input  [64-1:0] ar9ro1ql86jzmq_p,
  input  [5-1:0] qz1gqv6vh5qturw6v1mz,

  output y7rd1k0an54clel_5q6, 
  input  com03bquiktu249yb0, 
  output [64-1:0] tzg0yjgx9bn98i,
  output [4 -1:0] c2mipfm_6z5ef4p3aoz,
  output y3z8rf7c6hvsiux , 
  output [5-1:0] x8_a2j7z3gz3l0tfjqp,

  output xq0mj5mg2_512eu4, 
  input  e11m1298jo38qcwq9er2, 
  output [64-1:0] ec94_mk193di7tj,
  output [4 -1:0] m2sw40fca0wvnmy,
  output ywhfwlbfro2dmuvf ,
  output [5-1:0] nodrapn01yl1vxle30p,

  output ex_g_cnadtiu1r9u,
  input  orzasugx5h5pio22_,
  output [64-1:0] dxwtzud_wfj8jqk0,
  output [4 -1:0] gi8o690aydhqi8,
  output zl1r9cfvuhltjq ,
  output [5-1:0] dn074lh73rzchvrqzm8,

  output [64-1:0] xsn02pxoid_pw25,
  output [64-1:0] llv_dny70d,


  
  
  
  
  input  gc4b3kdcan6do88ta_,

  output j4xe_w_yjq2,
  output aui65oshqn8b5_iz6,
  output jmoafuo8zb_i1t,
  output sa5of37yr6xn0s3e,

  input  o5q5hev,
  input  o_dsdljul,
  input  juyzxopct4k03sl,
  input  qyqw_37_fxv8z,
  input  hyw0m71z3q3rpt1,
  input  fx_h7chccf02z,

  input  ru_wi
  );
  

  

  
  

  dv_v4v1au7ht_i2qt gycolq597t027sop7182(
    .w42_wd9um28vh (ehq614orwiy4ww5 ),
    .ssjx8h5cj3q4ffem (hgg2w2ca4wsixuj ),
    .rwby8vkzgm4y4r (lgv405vv46 ),
    .vuv0917fanv19 (vwxjizbv8c62_r6sf),
    .j2xzlc7dmxgmtn6kmk (ft8qpl2cvbar7ci),
    .tkxnzh2vh65vfutt3 (fi80hkldjwlh4v),
    
    .qd7ilyg140avze (vejdvgqormu727s),
    .n9uum984u41is66h2f (qz1gqv6vh5qturw6v1mz),
    .kf_pg4o0m8fa8 (ar9ro1ql86jzmq_p),
                                 
    .gc4b3kdcan6do88ta_     (gc4b3kdcan6do88ta_),
    .gf33atgy           (fx_h7chccf02z  ),
    .ru_wi         (ru_wi    ) 
  );















  
  
  wire bum_0_4oz7eoli40; 
  wire i53j9zqmffz8y6oqz7t; 
  wire zt7k3255akax0ouek346m;
  wire [64-1:0] vw3plvpp665o9dv9;
  wire [64-1:0] bzyry2czkd6xk6zjhye;
  wire [64-1:0] cp61fga88rjw8r82n3v;
  wire [48-1:0]  je_9freaj3uhcgylh63_;  
  wire [64-1:0] fqbjly2wnzhx63l;
  wire [4-1:0] bzjarqiyu0mfd0z3p;
  wire [3-1:0] v79ay3621ggo4h0d5aaj;


  
  
  wire kf2dpoq324swtgxgs6p; 
  wire l8kc7o3jpu34qr5q7; 
  wire zgtqckuiafu2aw2bjsy;
  wire [64-1:0] sw6wc3aq6kk892q79y32;
  wire [64-1:0] bgldh5yqcsal9_d;
  wire [64-1:0] pflh54d0tzca0r8_;
  wire [48-1:0]  rbuzk7rvhcg5f8qo25j;  
  wire [64-1:0] k1d77g2k6dmwycm9z8;
  wire [4-1:0] tkda6753pw4u9iq3ht;
  wire [3-1:0] win4d4amp0pkd57fchc;

  
  
  wire ywvgb6n56j5hgb2jrff; 
  wire cbk5zw3f620wbbj1dvrxi; 
  wire kisnmwl5fk22ydrmv4;
  wire [64-1:0] jf1prsiac8pb9waq4q;
  wire [64-1:0] utnh02m2bfr89kp;
  wire [64-1:0] nc5jui2ngra88qjivem;
  wire [48-1:0]  pr309tdfjv528m400czp;  
  wire [64-1:0] vchmkej8wq81b86w2qhu;
  wire [4-1:0] i0d65n3vieh6ywu9yts;
  wire [3-1:0] bucityy4pde4rrsrgrrqj;

  
  
  
  
  wire [64-1:0] m9fq2kwme4dt6asdh;
  wire [64-1:0] hebxwc_3illo41ep;
  wire [64-1:0] ak4g1lnf3qvbb;
  
  wire [64-1:0] nxrvop14jkb_1convg;
  

       wire [64-1:0] qpscc8xem = (oug11blpzcta8zyu0ya & o_qquv0pnx4zpz4h3gwxgl3) ? tmqkgmlzi018 : tmqkgmlzi018;
       wire [64-1:0] u3wdadynlf = (zr1pc8tfxyljdj7a8a3eh5 & j1fek3jzmt5bhhpnhvrmgt) ? lx_olubu7t8h : lx_olubu7t8h;
  wire [64-1:0] igvq6tvqkm = dd1p3tnenmm9r;
  assign xsn02pxoid_pw25 = m9fq2kwme4dt6asdh;
  assign llv_dny70d = hebxwc_3illo41ep;

  avxgym1nr_i6e h62uxxnv8vnv1bdx4kt(
    .yq7_jyt__u          (dkmuhc79d2wm0wubp  ),             
    .p1oz3zlyx9z099ko        (u2demhkod_er3kf6b),
    .i7xpott8rcin        (uz7pt71lvqit85od),
    .xfxtnu32e4          (qpscc8xem    ),
    .bzyabkjyg5aufwj          (u3wdadynlf    ),
    .w_vtk6165e          (igvq6tvqkm    ),
    .nog5k2tkaj_         (k9lv9ppimt14qx3d7rj       ),
    .a1nhqrkfzavps          (llskuqv0ehm60atlo        ),
    .p3g2fj0yq04eh         (v3uvhtx7e5vbtvie),
    .k1hmos4y13oq40h        (l60zv02z95hlayri),
    .hh9xkcr7e1fpzxae1ybn     (l1xzyldaa9dr2q7mla),

    .eg8yja9aryvtp8s      (rclkn1q60a3cbgtn67g     ),
    .ti187a_zcpeoww6gv     (ofmr0b7vez483r8wl    ),
    .zpr8r800wvts9w_mx     (zgn_d2n28xfn1zff    ),
    .gv1t0hwgea_5zw0eibk     (ceewyf1unn6p7peejem    ),
    .ccwkp0gpz76bmkrz     (oegl6jlhw01xkqeetu5y    ),
    .k8zoj8eu8lhoa3e82    (zamt9z8_hsjwlky8aktxv6   ),

    .q5h0basu9fqsocd     (a5z_23_ryr_m29hhia_p),
                         
    .bum_0_4oz7eoli40     (bum_0_4oz7eoli40   ),
    .i53j9zqmffz8y6oqz7t   (i53j9zqmffz8y6oqz7t ),
    .zt7k3255akax0ouek346m   (zt7k3255akax0ouek346m ),
    .vw3plvpp665o9dv9     (vw3plvpp665o9dv9   ),
    .bzyry2czkd6xk6zjhye     (bzyry2czkd6xk6zjhye   ),
    .cp61fga88rjw8r82n3v     (cp61fga88rjw8r82n3v   ),
    .je_9freaj3uhcgylh63_    (je_9freaj3uhcgylh63_  ),
    .fqbjly2wnzhx63l     (fqbjly2wnzhx63l   ),
    .bzjarqiyu0mfd0z3p    (bzjarqiyu0mfd0z3p  ),
    .v79ay3621ggo4h0d5aaj   (v79ay3621ggo4h0d5aaj  ),

    .kf2dpoq324swtgxgs6p     (kf2dpoq324swtgxgs6p   ),
    .l8kc7o3jpu34qr5q7   (l8kc7o3jpu34qr5q7 ),
    .zgtqckuiafu2aw2bjsy   (zgtqckuiafu2aw2bjsy ),
    .sw6wc3aq6kk892q79y32     (sw6wc3aq6kk892q79y32   ),
    .bgldh5yqcsal9_d     (bgldh5yqcsal9_d   ),
    .pflh54d0tzca0r8_     (pflh54d0tzca0r8_   ),
    .rbuzk7rvhcg5f8qo25j    (rbuzk7rvhcg5f8qo25j  ),
    .k1d77g2k6dmwycm9z8     (k1d77g2k6dmwycm9z8   ),
    .tkda6753pw4u9iq3ht    (tkda6753pw4u9iq3ht  ),
    .win4d4amp0pkd57fchc   (win4d4amp0pkd57fchc ),

    .ywvgb6n56j5hgb2jrff     (ywvgb6n56j5hgb2jrff   ),
    .cbk5zw3f620wbbj1dvrxi   (cbk5zw3f620wbbj1dvrxi ),
    .kisnmwl5fk22ydrmv4   (kisnmwl5fk22ydrmv4 ),
    .jf1prsiac8pb9waq4q     (jf1prsiac8pb9waq4q   ),
    .utnh02m2bfr89kp     (utnh02m2bfr89kp   ),
    .nc5jui2ngra88qjivem     (nc5jui2ngra88qjivem   ),
    .pr309tdfjv528m400czp    (pr309tdfjv528m400czp  ),
    .vchmkej8wq81b86w2qhu     (vchmkej8wq81b86w2qhu   ),
    .i0d65n3vieh6ywu9yts    (i0d65n3vieh6ywu9yts  ),
    .bucityy4pde4rrsrgrrqj   (bucityy4pde4rrsrgrrqj  ),

    .ddc4jxtzijwcnfg     (), 
    .h_ur90x_3ax0srnyj   (                ),
    .dytkvkta2hudyfw07   (1'b0            ),
    .xuixtwz82z81xfu02cgu     (m9fq2kwme4dt6asdh   ),
    .r1okty2iji67yzm9     (hebxwc_3illo41ep   ),
    .keu9vxu53w1s5zr     (ak4g1lnf3qvbb   ),
    .a0qgx1mu_gmlc7c6t5    (                ),
    .x0083y1q_m2c9h6     (nxrvop14jkb_1convg   ),
    .mdk0j4bk2l0pmkz25px_h (1'b0            ),
    .z94qawv75fwplf5ze90    ( ) 

  );

  wire frfkcvpr3s1e;
  
  wire g9ruu8swf4b_;
  wire eypswghjg4a5o;

  assign aui65oshqn8b5_iz6 = i53j9zqmffz8y6oqz7t
                        | frfkcvpr3s1e;
  assign sa5of37yr6xn0s3e = cbk5zw3f620wbbj1dvrxi
                        | g9ruu8swf4b_;
  assign jmoafuo8zb_i1t = l8kc7o3jpu34qr5q7
                        | eypswghjg4a5o;

  assign j4xe_w_yjq2 = u2demhkod_er3kf6b 
                    | aui65oshqn8b5_iz6
                    | sa5of37yr6xn0s3e
                    | jmoafuo8zb_i1t;

  drpp7_8vqsgvijw ph18q494f360ky6y(
    .eypswghjg4a5o         (eypswghjg4a5o),

    .cfk6xv54sxw51e          (kf2dpoq324swtgxgs6p),
    .ay4xay0aajxpqki        (zgtqckuiafu2aw2bjsy  ),
     
    .rx7xp4yfzkxxwe          (sw6wc3aq6kk892q79y32),
    .yh6637l46fxr          (bgldh5yqcsal9_d),
    .fx3oxnmunmg5         (rbuzk7rvhcg5f8qo25j),
    .ylzz2nmn2fx8vx         (tkda6753pw4u9iq3ht),
    .i7mguch8rrz_acmgw        (win4d4amp0pkd57fchc),

    .o1ic53wzueq3rdj        (xq0mj5mg2_512eu4   ),  
    .q5hfrt_ivi2var        (e11m1298jo38qcwq9er2   ),
    .xw5sonra6wr1qw86is7    (ec94_mk193di7tj    ),
    .zghahb2tb_ksbg78bg4   (nodrapn01yl1vxle30p    ),
    .u3_iseqd_x1swj1y1ikzv    (m2sw40fca0wvnmy    ),
    .aau8gpkszf2jvnjbmhfpm     (ywhfwlbfro2dmuvf     ),

    .gf33atgy           (qyqw_37_fxv8z  ),
    .ru_wi         (ru_wi    ) 
  );

  joupdqm1ityga9jgy gemk0xsjstmby903t(
    .frfkcvpr3s1e        (frfkcvpr3s1e),

    .rj9pxiv3u3_pir          (bum_0_4oz7eoli40),
    .b972jgf18d478vs1        (zt7k3255akax0ouek346m  ),
     
    .gurbf_74_clu          (vw3plvpp665o9dv9),
    .d1egtw92y1cy          (bzyry2czkd6xk6zjhye),
    .h501hw2_6          (cp61fga88rjw8r82n3v),
    .kiw03i3frj1_6         (je_9freaj3uhcgylh63_),
    .lw3kfp2bybej9         (bzjarqiyu0mfd0z3p),
    .ndsh540w8qc1oph        (v79ay3621ggo4h0d5aaj),

    .ct0b7_gmchg9rz        (y7rd1k0an54clel_5q6   ),  
    .xvcpof07ihp69zc        (com03bquiktu249yb0   ),
    .y3a80wegnmcxvkiw09    (tzg0yjgx9bn98i    ),
    .qngaib4rx7i91p4y2vv   (x8_a2j7z3gz3l0tfjqp    ),
    .bqcca4rpw2hdc6m1    (c2mipfm_6z5ef4p3aoz    ),
    .pjmhhc9l2dpz6y954     (y3z8rf7c6hvsiux     ),

    .gf33atgy           (juyzxopct4k03sl  ),
    .ru_wi         (ru_wi    ) 
  );

  iojbcv7tg90u tc3enfhvcly0ol(
    .g9ruu8swf4b_        (g9ruu8swf4b_),

    .aa9_kdx_kb35fx          (ywvgb6n56j5hgb2jrff),
    .z30wkcif1o8is5w9        (kisnmwl5fk22ydrmv4  ),
     
    .a4_acuaz1sfb5          (jf1prsiac8pb9waq4q),
    .q3ek793hh          (utnh02m2bfr89kp),
    .z1oylnyp4ryl4v         (pr309tdfjv528m400czp),
    .du24en2x_2qkjfw         (i0d65n3vieh6ywu9yts),
    .eyaonb2nm4ox        (bucityy4pde4rrsrgrrqj),

    .ycjcjdm1fjmdo_j        (ex_g_cnadtiu1r9u   ),  
    .j0s42ouqf5zv1a        (orzasugx5h5pio22_   ),
    .bqc9gh1yogik7q5r    (dxwtzud_wfj8jqk0    ),
    .dd4hyq5oe67rhyvoye   (dn074lh73rzchvrqzm8   ),
    .k4euvut15h32iq7j    (gi8o690aydhqi8    ),
    .b60gak_58icq19sfs_     (zl1r9cfvuhltjq     ),

    .gf33atgy           (hyw0m71z3q3rpt1  ),
    .ru_wi         (ru_wi    ) 
  );



endmodule                                      





















module p_nv4xk50a2bh9h4mr5fv #(
    parameter o10eaknnnv = 4
    ) (
    input [o10eaknnnv-1:0]           h1zifc6wetrm6wm,
    output [o10eaknnnv*o10eaknnnv-1:0]  oybz4sq2nhg8_26o,

    input gf33atgy,
    input ru_wi
    );


  genvar i,j;
  wire [o10eaknnnv-1:0] yy05l_vivocx9dom  [o10eaknnnv-1:0];
  wire [o10eaknnnv-1:0] qzntd3kydxpo8rx1ydoh [o10eaknnnv-1:0];
  wire [o10eaknnnv-1:0] nwnpreuq3zixor      [o10eaknnnv-1:0];

  generate
    for (i=0;i<o10eaknnnv;i=i+1) begin :aifg64k59ey5b
      for (j=0;j<o10eaknnnv;j=j+1) begin :mwzjcdc_
        if (i < j) begin:ewf64owjec

          assign yy05l_vivocx9dom[i][j] = h1zifc6wetrm6wm[i] || h1zifc6wetrm6wm[j];
          assign qzntd3kydxpo8rx1ydoh[i][j]= h1zifc6wetrm6wm[i] ? 1'b1 :
                                          h1zifc6wetrm6wm[j] ? 1'b0 :
                                                            1'b0 ;
          ux607_gnrl_dfflr #(1) zg3vvxtlq8 (yy05l_vivocx9dom[i][j], qzntd3kydxpo8rx1ydoh[i][j], nwnpreuq3zixor[i][j], gf33atgy, ru_wi);
        end 
        else begin:gf05giycnv394ndz
          assign yy05l_vivocx9dom[i][j] = 1'b0;
          assign qzntd3kydxpo8rx1ydoh[i][j] = 1'b0;
          assign nwnpreuq3zixor[i][j] = 1'b0;
        end
      end
    end
  endgenerate

  generate
    for (i=0;i<o10eaknnnv;i=i+1) begin :znl924vwl86injct
      assign oybz4sq2nhg8_26o[i*o10eaknnnv+:o10eaknnnv] = nwnpreuq3zixor[i][o10eaknnnv-1:0];
    end
  endgenerate 

endmodule



















module ux607_gnrl_pipe_stage # (


  parameter CUT_READY = 0,
  parameter DP = 1,
  parameter DW = 32
) (
  input           i_vld, 
  output          i_rdy, 
  input  [DW-1:0] i_dat,
  output          o_vld, 
  input           o_rdy, 
  output [DW-1:0] o_dat,

  input           clk,
  input           rst_n
);

  genvar i;
  generate 

  if(DP == 0) begin: kum1oxhw1b434q

      assign o_vld = i_vld;
      assign i_rdy = o_rdy;
      assign o_dat = i_dat;

  end
  else begin: r1f9lplxw0lya5z

      wire d35brwhbkm;
      wire xlzi7_mjg;
      wire xayqet0sd;
      wire ycgzbt;
      wire d0x7t39v;


      assign d35brwhbkm = i_vld & i_rdy;

      assign xlzi7_mjg = o_vld & o_rdy;

      assign xayqet0sd = d35brwhbkm | xlzi7_mjg;
      assign d0x7t39v = d35brwhbkm | (~xlzi7_mjg);

      ux607_gnrl_dfflr #(1) hdti_6iaq (xayqet0sd, d0x7t39v, ycgzbt, clk, rst_n);

      assign o_vld = ycgzbt;

      ux607_gnrl_dffl #(DW) tn7qvilprku (d35brwhbkm, i_dat, o_dat, clk, rst_n);

      if(CUT_READY == 1) begin:lvfon_zgkwp229

          assign i_rdy = (~ycgzbt);
      end
      else begin:ulbqsqnmhe2qhizmyx

          assign i_rdy = (~ycgzbt) | xlzi7_mjg;
      end
  end
  endgenerate


endmodule 








module ux607_gnrl_sync # (
  parameter DP = 2,
  parameter DW = 32
) (
  input  [DW-1:0] din_a,
  output [DW-1:0] dout,

  input           rst_n, 
  input           clk 
);

  wire [DW-1:0] hq1mzczr [DP-1:0];

  genvar i;

  generate 
    for(i=0;i<DP;i=i+1) begin:xgpq9q044nj
      if(i==0) begin:xvpcp9wjmb99kn
        ux607_gnrl_dffr #(DW) zjzw8_1bsf2xfe(din_a,         hq1mzczr[0], clk, rst_n);
      end
      else begin:efbb_rw4_pjzu4jx64w
        ux607_gnrl_dffr #(DW) zjzw8_1bsf2xfe(hq1mzczr[i-1], hq1mzczr[i], clk, rst_n);
      end
    end
  endgenerate

  assign dout = hq1mzczr[DP-1];

endmodule







module ux607_gnrl_rrobin # (
    parameter ARBT_NUM = 4
)(
  output[ARBT_NUM-1:0] grt_vec,  
  input [ARBT_NUM-1:0] req_vec,  
  input arbt_ena,   
  input clk,        
  input rst_n
);

wire               f8li874yxsa;
wire               gr86ihf0sej0;
wire               s1wlajyjpsy9;
wire [ARBT_NUM-1:0] irn9wwe3yz;
wire [ARBT_NUM-1:0] g6dxux10;  

wire [ARBT_NUM-1:0] g_nts5e01i7wzs18;
wire [ARBT_NUM-1:0] l1zpeyxktr5yuw6y8skkp;
assign g_nts5e01i7wzs18[0] = req_vec[0];
genvar i;
generate
  for(i = 1; i < ARBT_NUM; i = i+1)
  begin:bs_isce2_
    assign g_nts5e01i7wzs18[i] = |req_vec[i-1:0];
  end
endgenerate

assign l1zpeyxktr5yuw6y8skkp = {g_nts5e01i7wzs18[ARBT_NUM-2:0],1'b0};

wire [ARBT_NUM-1:0] di198vx7h_6jz47mttgzzchlo;
assign di198vx7h_6jz47mttgzzchlo= l1zpeyxktr5yuw6y8skkp & req_vec;


wire lqa78v8dlc61bn1eunnr = ~(|di198vx7h_6jz47mttgzzchlo);

wire rwybdxe8m84q_z8r7j6 = (|req_vec);
wire bhrkh6058njsyuvz9c6ye  = ~lqa78v8dlc61bn1eunnr;
assign f8li874yxsa = rwybdxe8m84q_z8r7j6 & bhrkh6058njsyuvz9c6ye;
assign gr86ihf0sej0  = f8li874yxsa & arbt_ena;
assign irn9wwe3yz = s1wlajyjpsy9 ? {ARBT_NUM{1'b1}} : g6dxux10 << 1;


generate
  if(ARBT_NUM == 2) begin: e9ads2qqsvc68oz3
    assign s1wlajyjpsy9 = ~(g6dxux10[0]);
  end 
  else begin: mg2ol_ht6p__9utpk
    assign s1wlajyjpsy9 = ~(|g6dxux10[ARBT_NUM-2:0]);
  end
endgenerate

ux607_gnrl_dfflrs #(ARBT_NUM) f2pipltedja (gr86ihf0sej0, irn9wwe3yz, g6dxux10, clk, rst_n);



wire [ARBT_NUM-1:0] tk7o1p3c_ihk8nm8e;
wire [ARBT_NUM-1:0] zaekp6ng4fyw32gp;
wire [ARBT_NUM-1:0] abf5c98n61utwudxn4dhy;
wire [ARBT_NUM-1:0] zits6wm1yr;
wire [ARBT_NUM-1:0] gsbztf6ye5g5rw;      
wire [ARBT_NUM-1:0] a3wwuk1z8b2u5etka;
wire [ARBT_NUM-1:0] idsm6llc5u;
wire [ARBT_NUM-1:0] e75s18podfpe;      

wire [ARBT_NUM-1:0] c0_fjr1ekbr;          
wire [ARBT_NUM-1:0] fyawtijy0_mr;          
wire pjd96vtarupx;          
wire d8_oitpk;          
wire iq56_qt5shnc4;          

assign d8_oitpk = (|grt_vec) & (~arbt_ena);          
assign iq56_qt5shnc4 = arbt_ena;          
assign pjd96vtarupx = d8_oitpk | iq56_qt5shnc4;          
assign fyawtijy0_mr = iq56_qt5shnc4 ? {ARBT_NUM{1'b0}} : (~grt_vec);

ux607_gnrl_dfflr #(ARBT_NUM) vazepyge_wr (pjd96vtarupx, fyawtijy0_mr, c0_fjr1ekbr, clk, rst_n);



wire [ARBT_NUM-1:0] qcu69vmnak6r0jm24;          
assign qcu69vmnak6r0jm24 = req_vec & (~c0_fjr1ekbr);          

assign tk7o1p3c_ihk8nm8e = g6dxux10 & qcu69vmnak6r0jm24;
assign zaekp6ng4fyw32gp = (~g6dxux10) & qcu69vmnak6r0jm24;

generate
  for(i = 0; i < ARBT_NUM; i = i+1)
  begin:tbba994dc372zdu4dbjg
    if(i==0) begin: i6ktna73ot
      assign abf5c98n61utwudxn4dhy[0] = tk7o1p3c_ihk8nm8e[0];
      assign a3wwuk1z8b2u5etka[0] = zaekp6ng4fyw32gp[0];
      assign zits6wm1yr[0] = abf5c98n61utwudxn4dhy[0];
      assign idsm6llc5u[0] = a3wwuk1z8b2u5etka[0];
    end
    else begin: raoucdzq_4
      assign abf5c98n61utwudxn4dhy[i] = |tk7o1p3c_ihk8nm8e[i:0];
      assign a3wwuk1z8b2u5etka[i] = |zaekp6ng4fyw32gp[i:0];
      assign zits6wm1yr[i] = (~abf5c98n61utwudxn4dhy[i-1]) & abf5c98n61utwudxn4dhy[i];
      assign idsm6llc5u[i] = (~a3wwuk1z8b2u5etka[i-1]) & a3wwuk1z8b2u5etka[i];
    end
  end
endgenerate

assign gsbztf6ye5g5rw = zits6wm1yr;
assign e75s18podfpe = idsm6llc5u;

wire helu0kms = |(g6dxux10 & qcu69vmnak6r0jm24);

assign grt_vec = helu0kms ?  gsbztf6ye5g5rw : e75s18podfpe;

endmodule








module ux607_gnrl_cdc_rx
# (
  parameter DW = 32,
  parameter SYNC_DP = 2
) (






  input  i_vld_a, 
  output i_rdy, 
  input  [DW-1:0] i_dat,


  output o_vld, 
  input  o_rdy, 
  output [DW-1:0] o_dat,

  input  clk,
  input  rst_n 
);

wire z12rq5w2beus9e;

ux607_gnrl_sync #(.DP(SYNC_DP), .DW(1)) c2kpioqhczag (
     .clk   (clk),
     .rst_n (rst_n),
     .din_a (i_vld_a),
     .dout  (z12rq5w2beus9e)
    );

wire kbd70p3fy4lm1kv;
ux607_gnrl_dffr #(1) a4s_1yp4ykjuqeo(z12rq5w2beus9e, kbd70p3fy4lm1kv, clk, rst_n);
wire n7y6pqu2ztlgek8ilm = (~z12rq5w2beus9e) & kbd70p3fy4lm1kv;

wire ibm81_gpcaa;
wire yo_gmsn;



wire d3l8fkcc7r3k = ibm81_gpcaa & z12rq5w2beus9e & (~yo_gmsn);
wire d838764py = n7y6pqu2ztlgek8ilm;
wire s1tkq4o_fpxmau = d3l8fkcc7r3k |   d838764py;
wire x2hmpfi0j9 = d3l8fkcc7r3k | (~d838764py);
ux607_gnrl_dfflr #(1) dyluac1_hk_3(s1tkq4o_fpxmau, x2hmpfi0j9, yo_gmsn, clk, rst_n);
assign i_rdy = yo_gmsn;


wire pppcao07cf2;
wire [DW-1:0] p5d9udwxfrj6;



wire hwg_mzj91ik3 = d3l8fkcc7r3k;
ux607_gnrl_dfflr #(DW) mbvgfav9scrcwpjy(hwg_mzj91ik3, i_dat, p5d9udwxfrj6, clk, rst_n);


wire crj8ju_avbpyfzw = hwg_mzj91ik3;

wire d94r1t3t4611r_d = o_vld & o_rdy;
wire j2icql4g_flg = crj8ju_avbpyfzw | d94r1t3t4611r_d;
wire enthl38h0f7j47 = crj8ju_avbpyfzw | (~d94r1t3t4611r_d);
ux607_gnrl_dfflr #(1) b_l4hs2nvep0t9g(j2icql4g_flg, enthl38h0f7j47, pppcao07cf2, clk, rst_n);

assign ibm81_gpcaa = (~pppcao07cf2);

assign o_vld = pppcao07cf2;
assign o_dat = p5d9udwxfrj6;

endmodule 











module ux607_gnrl_cdc_tx
# (
  parameter DW = 32,
  parameter SYNC_DP = 2
) (


  input  i_vld, 
  output i_rdy, 
  input  [DW-1:0] i_dat,







  output o_vld, 
  input  o_rdy_a, 
  output [DW-1:0] o_dat,

  input  clk,
  input  rst_n 
);

wire kzr1g_mdx_0;


ux607_gnrl_sync #(
    .DP(SYNC_DP), 
    .DW(1)
) xz7fyd05mq8yc9n (
         .clk   (clk),
         .rst_n (rst_n),
         .din_a (o_rdy_a),
         .dout  (kzr1g_mdx_0)
        );

wire ycgzbt;
wire [DW-1:0] c37pfa;


wire d35brwhbkm = i_vld & i_rdy;

wire xlzi7_mjg = o_vld & kzr1g_mdx_0;
wire xayqet0sd = d35brwhbkm | xlzi7_mjg;
wire d0x7t39v = d35brwhbkm | (~xlzi7_mjg);
ux607_gnrl_dfflr #(1) hdti_6iaq(xayqet0sd, d0x7t39v, ycgzbt, clk, rst_n);

ux607_gnrl_dfflr #(DW) tn7qvilprku(d35brwhbkm, i_dat, c37pfa, clk, rst_n);


wire rqq8wcvzx53dhnw;
ux607_gnrl_dffr #(1) g0cjr_eg_hnon2li(kzr1g_mdx_0, rqq8wcvzx53dhnw, clk, rst_n);
wire ij66ap_p1pq9g3n = (~kzr1g_mdx_0) & rqq8wcvzx53dhnw;


wire wdrid04qp0u;

wire wmnujevga2 = d35brwhbkm;

wire t17hjolm9l = ij66ap_p1pq9g3n;
wire bn10iistuty6 = wmnujevga2 | t17hjolm9l;
wire iobyipyut = wmnujevga2 | (~t17hjolm9l);
ux607_gnrl_dfflr #(1) xlw1j6ei2_0ob5_x8(bn10iistuty6, iobyipyut, wdrid04qp0u, clk, rst_n);


assign o_vld = ycgzbt;

assign o_dat = c37pfa;


assign i_rdy = (~wdrid04qp0u) | t17hjolm9l;

endmodule 








module ux607_gnrl_bypbuf # (
  parameter DP = 8,
  parameter DW = 32
) (
  input           i_vld,
  output          i_rdy,
  input  [DW-1:0] i_dat,

  output          o_vld,
  input           o_rdy,
  output [DW-1:0] o_dat,

  input           clk,
  input           rst_n
);


  wire          zvyiwdpyvt;
  wire          o0ozobxf1oc2t5;
  wire [DW-1:0] jf92hqkj0cxz;

  wire          mgjqsgpiza1dr;
  wire          qos62pcur8;
  wire [DW-1:0] jae1i1kz83d2c;

  ux607_gnrl_fifo # (
       .DP(DP),
       .DW(DW),
       .CUT_READY(1) 
  ) tk61pi32v0g9or0o3v(
    .i_vld   (zvyiwdpyvt),
    .i_rdy   (o0ozobxf1oc2t5),
    .i_dat   (jf92hqkj0cxz),
    .o_vld   (mgjqsgpiza1dr),
    .o_rdy   (qos62pcur8),
    .o_dat   (jae1i1kz83d2c),
    .clk     (clk  ),
    .rst_n   (rst_n)
  );




  assign i_rdy = o0ozobxf1oc2t5;



  wire fzf_yfd = i_vld & o_rdy & (~mgjqsgpiza1dr);


  assign qos62pcur8 = o_rdy;


  assign o_vld = mgjqsgpiza1dr | i_vld;


  assign o_dat = mgjqsgpiza1dr ? jae1i1kz83d2c : i_dat;

  assign jf92hqkj0cxz  = i_dat; 


  assign zvyiwdpyvt = i_vld & (~fzf_yfd);


endmodule 










module hs5vxvpng41zt1s2gdyu6psryf # (
  parameter mhdlk = 8,
  parameter onr7l = 32
) (
  input           fz8gtuc,

  input           bw6ftrau0,
  output          eef2g8,
  input  [onr7l-1:0] qbjvs30wtb,

  output          wqljp,
  input           h9378,
  output [onr7l-1:0] dqgck5s,

  input           gf33atgy,
  input           ru_wi
);


  wire          zvyiwdpyvt;
  wire          o0ozobxf1oc2t5;
  wire [onr7l-1:0] jf92hqkj0cxz;

  wire          mgjqsgpiza1dr;
  wire          qos62pcur8;
  wire [onr7l-1:0] jae1i1kz83d2c;

  vq28fpkbg0dxljs8bf0k # (
       .hejad2_b4dywimoxw5(1),
       .evi4vkasjp742kf4(1),
       .mhdlk(mhdlk),
       .onr7l(onr7l)
  ) wz_vb6ba3vsy0log02u7(
    .geml8twgru(fz8gtuc),
    .td5hjljc_(fz8gtuc),
    .bw6ftrau0   (zvyiwdpyvt),
    .eef2g8   (o0ozobxf1oc2t5),
    .qbjvs30wtb   (jf92hqkj0cxz),
    .wqljp   (mgjqsgpiza1dr),
    .h9378   (qos62pcur8),
    .dqgck5s   (jae1i1kz83d2c),
    .i0lklnhw28rc7dj(),
    .gf33atgy     (gf33atgy  ),
    .ru_wi   (ru_wi)
  );




  assign eef2g8 = o0ozobxf1oc2t5;



  wire fzf_yfd = bw6ftrau0 & h9378 & (~mgjqsgpiza1dr);


  assign qos62pcur8 = h9378;


  assign wqljp = mgjqsgpiza1dr | bw6ftrau0;


  assign dqgck5s = mgjqsgpiza1dr ? jae1i1kz83d2c : qbjvs30wtb;

  assign jf92hqkj0cxz  = qbjvs30wtb; 


  assign zvyiwdpyvt = bw6ftrau0 & (~fzf_yfd);


endmodule 










module ux607_gnrl_fifo # (







  parameter CUT_READY = 0,
  parameter MSKO = 0,
  parameter DP   = 8,
  parameter DW   = 32
) (

  input           i_vld, 
  output          i_rdy, 
  input  [DW-1:0] i_dat,
  output          o_vld, 
  input           o_rdy, 
  output [DW-1:0] o_dat,

  input           clk,
  input           rst_n
);

genvar i;
generate 

  if(DP == 0) begin: o3wv6_2_uu

     assign o_vld = i_vld;
     assign i_rdy = o_rdy;
     assign o_dat = i_dat;

  end
  else begin: ggp3zuzuwf9w87z


    wire [DW-1:0] w2z87rfaf8 [DP-1:0];
    wire [DP-1:0] k8cq9veedzws;


    wire kxaplzy = i_vld & i_rdy;
    wire fumg8 = o_vld & o_rdy;



    wire [DP-1:0] tzr9_pu0gkgq459gy; 
    wire [DP-1:0] dz1thuu43r;
    wire [DP-1:0] kv5lv5mhl4m9_kh; 
    wire [DP-1:0] wxlsjrqo2a;

    if(DP == 1) begin:g9_p9c0apem00fcj_
      assign tzr9_pu0gkgq459gy = 1'b1; 
    end
    else begin:k05cliuyoxplv354gkh
      assign tzr9_pu0gkgq459gy = 
          dz1thuu43r[DP-1] ? {{DP-1{1'b0}}, 1'b1} :
                          (dz1thuu43r << 1);
    end

    if(DP == 1) begin:kzd56tqvj_6_wu
      assign kv5lv5mhl4m9_kh = 1'b1; 
    end
    else begin:vm1yxa6ea3yg5lu56c_jbw
      assign kv5lv5mhl4m9_kh =
          wxlsjrqo2a[DP-1] ? {{DP-1{1'b0}}, 1'b1} :
                          (wxlsjrqo2a << 1);
    end

    ux607_gnrl_dfflrs #(1)    qnwogo1l036nyvzk_i  (fumg8, tzr9_pu0gkgq459gy[0]     , dz1thuu43r[0]     , clk, rst_n);
    ux607_gnrl_dfflrs #(1)    mn4pzjreki9yvykae  (kxaplzy, kv5lv5mhl4m9_kh[0]     , wxlsjrqo2a[0]     , clk, rst_n);
    if(DP > 1) begin:rujquo369cvzmr5
    ux607_gnrl_dfflr  #(DP-1) fipb6zpafcl9yge96au  (fumg8, tzr9_pu0gkgq459gy[DP-1:1], dz1thuu43r[DP-1:1], clk, rst_n);
    ux607_gnrl_dfflr  #(DP-1) hh9891_eoeau0wkyll5  (kxaplzy, kv5lv5mhl4m9_kh[DP-1:1], wxlsjrqo2a[DP-1:1], clk, rst_n);
    end



    wire [DP:0] uipdtjs;
    wire [DP:0] acm0zbhvam;
    wire [DP:0] oi40qurrxr; 
    wire [DP:0] n89fv;

    wire jlo7_b_z = (fumg8 ^ kxaplzy );
    assign oi40qurrxr = kxaplzy ? {n89fv[DP-1:0], 1'b1} : (n89fv >> 1);  

    ux607_gnrl_dfflrs #(1)  svv3sz17bdpp     (jlo7_b_z, oi40qurrxr[0]     , n89fv[0]     ,     clk, rst_n);
    ux607_gnrl_dfflr  #(DP) j3hui4o9q5lg     (jlo7_b_z, oi40qurrxr[DP:1], n89fv[DP:1],     clk, rst_n);

    assign uipdtjs = {1'b0,n89fv[DP:1]};
    assign acm0zbhvam = {1'b0,n89fv[DP:1]};

    if(DP == 1) begin:tv7hfw9czbztt19
        if(CUT_READY == 1) begin:lvfon_zgkwp229

          assign i_rdy = (~uipdtjs[DP-1]);
        end
        else begin:ulbqsqnmhe2qhizmyx

          assign i_rdy = (~uipdtjs[DP-1]) | fumg8;
        end
    end
    else begin : ums8cgjwy0afp93
      assign i_rdy = (~uipdtjs[DP-1]);
    end



    for (i=0; i<DP; i=i+1) begin:m_wwntxzhohqg5
      assign k8cq9veedzws[i] = kxaplzy & wxlsjrqo2a[i];

      ux607_gnrl_dfflr  #(DW) anynep9ymzbmqsgf (k8cq9veedzws[i], i_dat, w2z87rfaf8[i], clk, rst_n);
    end


    integer j;
    reg [DW-1:0] ui9y38d1t;
    always @*
    begin : e82692n5bc4eh
      ui9y38d1t = {DW{1'b0}};
      for(j=0; j<DP; j=j+1) begin
        ui9y38d1t = ui9y38d1t | ({DW{dz1thuu43r[j]}} & w2z87rfaf8[j]);
      end
    end

    if(MSKO == 1) begin:nxdryocmrcvmkh54cu_9

        assign o_dat = {DW{o_vld}} & ui9y38d1t;
    end
    else begin:lkweycxyox5vpftvd1yym7

        assign o_dat = ui9y38d1t;
    end


    assign o_vld = (acm0zbhvam[0]);

  end
endgenerate

endmodule 










module vq28fpkbg0dxljs8bf0k # (
  parameter hejad2_b4dywimoxw5 = 0,
  parameter evi4vkasjp742kf4 = 0,
  parameter mhdlk   = 8,
  parameter onr7l   = 32
) (

  input           geml8twgru,

  input           bw6ftrau0, 
  output          eef2g8, 
  input  [onr7l-1:0] qbjvs30wtb,


  input           td5hjljc_,

  output          wqljp, 
  input           h9378, 
  output [onr7l-1:0] dqgck5s,

  output          i0lklnhw28rc7dj,

  input           gf33atgy,
  input           ru_wi
);


genvar i;
generate 

  if(mhdlk == 0) begin: o3wv6_2_uu

     assign wqljp = bw6ftrau0;
     assign eef2g8 = h9378;
     assign dqgck5s = qbjvs30wtb;
     assign i0lklnhw28rc7dj =  1'b0;

  end
  else begin: ggp3zuzuwf9w87z



    wire [onr7l-1:0] w2z87rfaf8 [mhdlk-1:0];
    wire [mhdlk-1:0] k8cq9veedzws;


    wire kxaplzy = bw6ftrau0 & eef2g8 & geml8twgru;
    wire fumg8 = wqljp & h9378 & td5hjljc_;



    wire [mhdlk-1:0] tzr9_pu0gkgq459gy; 
    wire [mhdlk-1:0] dz1thuu43r;
    wire [mhdlk-1:0] kv5lv5mhl4m9_kh; 
    wire [mhdlk-1:0] wxlsjrqo2a;

      if (mhdlk == 1) begin:nunbyyrd2bei03kp
          assign tzr9_pu0gkgq459gy = 1'b1;
          assign kv5lv5mhl4m9_kh = 1'b1;
      end 
      else begin:jh8ttlqf8d3zs1fvgewi
          assign tzr9_pu0gkgq459gy = 
            dz1thuu43r[mhdlk-1] ? {{mhdlk-1{1'b0}}, 1'b1} :
                            (dz1thuu43r << 1);
          assign kv5lv5mhl4m9_kh =
            wxlsjrqo2a[mhdlk-1] ? {{mhdlk-1{1'b0}}, 1'b1} :
                            (wxlsjrqo2a << 1);
      end


    ux607_gnrl_dfflrs #(1)    qnwogo1l036nyvzk_i  (fumg8, tzr9_pu0gkgq459gy[0]     , dz1thuu43r[0]     , gf33atgy, ru_wi);
    ux607_gnrl_dfflrs #(1)    mn4pzjreki9yvykae  (kxaplzy, kv5lv5mhl4m9_kh[0]     , wxlsjrqo2a[0]     , gf33atgy, ru_wi);
      if(mhdlk>1) begin:rujquo369cvzmr5
         ux607_gnrl_dfflr  #(mhdlk-1) fipb6zpafcl9yge96au  (fumg8, tzr9_pu0gkgq459gy[mhdlk-1:1], dz1thuu43r[mhdlk-1:1], gf33atgy, ru_wi);
         ux607_gnrl_dfflr  #(mhdlk-1) hh9891_eoeau0wkyll5  (kxaplzy, kv5lv5mhl4m9_kh[mhdlk-1:1], wxlsjrqo2a[mhdlk-1:1], gf33atgy, ru_wi);
      end



    wire [mhdlk:0] uipdtjs;
    wire [mhdlk:0] acm0zbhvam;
    wire [mhdlk:0] oi40qurrxr; 
    wire [mhdlk:0] n89fv;

    wire jlo7_b_z = (fumg8 ^ kxaplzy );
    assign oi40qurrxr = kxaplzy ? {n89fv[mhdlk-1:0], 1'b1} : (n89fv >> 1);  

    ux607_gnrl_dfflrs #(1)  svv3sz17bdpp     (jlo7_b_z, oi40qurrxr[0]     , n89fv[0]     ,     gf33atgy, ru_wi);
    ux607_gnrl_dfflr  #(mhdlk) j3hui4o9q5lg     (jlo7_b_z, oi40qurrxr[mhdlk:1], n89fv[mhdlk:1],     gf33atgy, ru_wi);

    assign uipdtjs = {1'b0,n89fv[mhdlk:1]};
    assign acm0zbhvam = {1'b0,n89fv[mhdlk:1]};

  wire cds3152c6iisjx;
  if (!hejad2_b4dywimoxw5) begin : ztfii8187qhhtkw9
    assign eef2g8 = (~uipdtjs[mhdlk-1]);
    assign cds3152c6iisjx = 1'b0;
  end
  else begin
    wire l_ehdje55iwjqc6;
    wire h8p9a9dnu1urx2;
    wire yo_gmsn;
    wire gz9qt0181m7xl;
    wire aahd54_6alaloln04qn;
    wire ztc38ot3jhq5etl5ef67a;
    wire w3tf_jr90pvogxsu72u8ap;
    wire mnlyuiaq_evcghkx5bhfxy;
    wire h0a65gmxxcpara5pf;
    assign gz9qt0181m7xl = jlo7_b_z; 
    assign aahd54_6alaloln04qn = (gz9qt0181m7xl && !geml8twgru);
    assign ztc38ot3jhq5etl5ef67a = (h0a65gmxxcpara5pf && geml8twgru);
    assign w3tf_jr90pvogxsu72u8ap = aahd54_6alaloln04qn || ztc38ot3jhq5etl5ef67a;
    assign mnlyuiaq_evcghkx5bhfxy = aahd54_6alaloln04qn;
    ux607_gnrl_dfflr  #(1) jm5hpo5kmcdpk736me9zfs1sa    (w3tf_jr90pvogxsu72u8ap, mnlyuiaq_evcghkx5bhfxy, h0a65gmxxcpara5pf,     gf33atgy, ru_wi);

    assign l_ehdje55iwjqc6 = geml8twgru && (gz9qt0181m7xl || h0a65gmxxcpara5pf);
    assign h8p9a9dnu1urx2 = (jlo7_b_z) ? (~oi40qurrxr[mhdlk]) : (~uipdtjs[mhdlk-1]);
    ux607_gnrl_dfflrs  #(1) zqxw503ze_semtw81i4    (l_ehdje55iwjqc6, h8p9a9dnu1urx2, yo_gmsn,     gf33atgy, ru_wi);
    assign eef2g8 = yo_gmsn;
    assign cds3152c6iisjx = h0a65gmxxcpara5pf;
  end


    for (i=0; i<mhdlk; i=i+1) begin:m_wwntxzhohqg5
      assign k8cq9veedzws[i] = kxaplzy & wxlsjrqo2a[i];

      ux607_gnrl_dfflr  #(onr7l) anynep9ymzbmqsgf (k8cq9veedzws[i], qbjvs30wtb, w2z87rfaf8[i], gf33atgy, ru_wi);
    end


    integer j;
    reg [onr7l-1:0] ui9y38d1t;
    always @*
    begin : e82692n5bc4eh
      ui9y38d1t = {onr7l{1'b0}};
      for(j=0; j<mhdlk; j=j+1) begin
        ui9y38d1t = ui9y38d1t | ({onr7l{dz1thuu43r[j]}} & w2z87rfaf8[j]);
      end
    end


    assign dqgck5s = ui9y38d1t & {onr7l{wqljp}};

  wire olrdw6s_d_1bnbf9j;
  if (!evi4vkasjp742kf4) begin : vgavgfjzf293iy5b

    assign wqljp = (acm0zbhvam[0]);
    assign olrdw6s_d_1bnbf9j = 1'b0;
  end
  else begin : jv69teibe7a4   
    wire fnompgcuoys3av;
    wire cqjuz__0d5wryt;
    wire mxqwnph;
    wire l2kwhv43umaib;
    wire y9phf0tdehb0aev83ri;
    wire tr_pczcm87014ah6h9;
    wire w5tjv7yt39rnigu_u_l;
    wire lmanup378q1qzwldb5;
    wire kun4jk6p0x4b2bao34n;
    assign l2kwhv43umaib = jlo7_b_z;
    assign y9phf0tdehb0aev83ri = (l2kwhv43umaib   && !td5hjljc_);
    assign tr_pczcm87014ah6h9 = (kun4jk6p0x4b2bao34n &&  td5hjljc_);
    assign w5tjv7yt39rnigu_u_l = y9phf0tdehb0aev83ri || tr_pczcm87014ah6h9;
    assign lmanup378q1qzwldb5 = y9phf0tdehb0aev83ri;
    ux607_gnrl_dfflr  #(1) bgspwk95kxsppsiarqazq7sm    (w5tjv7yt39rnigu_u_l, lmanup378q1qzwldb5, kun4jk6p0x4b2bao34n,     gf33atgy, ru_wi);

    assign fnompgcuoys3av = td5hjljc_ && (l2kwhv43umaib || kun4jk6p0x4b2bao34n);
    assign cqjuz__0d5wryt = (jlo7_b_z) ? (oi40qurrxr[1]) : (acm0zbhvam[0]);
    ux607_gnrl_dfflr  #(1) mkv2_cnjr4yvhbizcx    (fnompgcuoys3av, cqjuz__0d5wryt, mxqwnph,     gf33atgy, ru_wi);
    assign wqljp = mxqwnph;

    assign olrdw6s_d_1bnbf9j = kun4jk6p0x4b2bao34n;

  end

  assign i0lklnhw28rc7dj =  bw6ftrau0 || cds3152c6iisjx || wqljp || olrdw6s_d_1bnbf9j;

  end
endgenerate

endmodule 








module togf4n__xsiylxzli0xu5ty3 # (
    parameter mhdlk = 4,
    parameter onr7l = 32
)(
    input  u22pp,
    input  irka0,


    input  [onr7l-1:0] qbjvs30wtb,
    output [onr7l-1:0] dqgck5s,

    input  gf33atgy,
    input  ru_wi
);

  wire [onr7l-1:0] olf4xmxku9u9k8 [mhdlk-1:0];
  wire [mhdlk-1:0] cryhplg9_24tqw;



  wire [mhdlk-1:0] uipdtjs;
  wire [mhdlk-1:0] acm0zbhvam;
  wire [mhdlk-1:0] oi40qurrxr; 
  wire [mhdlk-1:0] n89fv;

  wire jlo7_b_z = (irka0 ^ u22pp);
  assign oi40qurrxr =     irka0 ? 
                   (n89fv[0] ? {1'b1,{mhdlk-1{1'b0}}} : (n89fv >> 1)) :
                (n89fv[mhdlk-1] ? {{mhdlk-1{1'b0}},1'b1} : (n89fv << 1))
                             ;  

  ux607_gnrl_dfflrs #(1)    svv3sz17bdpp(jlo7_b_z, oi40qurrxr[0]     , n89fv[0]     , gf33atgy, ru_wi);
  ux607_gnrl_dfflr  #(mhdlk-1) o0mc8mg4cq9iqbw(jlo7_b_z, oi40qurrxr[mhdlk-1:1], n89fv[mhdlk-1:1], gf33atgy, ru_wi);


  assign uipdtjs = n89fv; 
  assign acm0zbhvam = (n89fv == {{mhdlk-1{1'b0}},1'b1}) ? {1'b1, {mhdlk-1{1'b0}}}
                                                : (n89fv >> 1); 

  genvar i;
  generate 

    for (i=0; i<mhdlk; i=i+1) begin:eyoclcjcy41
      assign cryhplg9_24tqw[i] = u22pp & uipdtjs[i];      
      ux607_gnrl_dfflr  #(onr7l) s3y1py6je3tms (cryhplg9_24tqw[i], qbjvs30wtb, olf4xmxku9u9k8[i], gf33atgy, ru_wi);
    end
  endgenerate


  integer j;
  reg [onr7l-1:0] ui9y38d1t;
  always @*
  begin : e82692n5bc4eh
    ui9y38d1t = {onr7l{1'b0}};
    for(j=0; j<mhdlk; j=j+1) begin
      ui9y38d1t = ui9y38d1t | ({onr7l{acm0zbhvam[j]}} & olf4xmxku9u9k8[j]);
    end
  end

  assign dqgck5s = ui9y38d1t;

endmodule










module m4ye826sgj3blndc # (
  parameter mhdlk   = 8,
  parameter onr7l   = 32
) (

  input           u22pp, 
  input  [onr7l-1:0] qbjvs30wtb,
  input           irka0, 
  output [onr7l-1:0] dqgck5s,

  input           gf33atgy,
  input           ru_wi
);




  wire [onr7l-1:0] olf4xmxku9u9k8 [mhdlk-1:0];
  wire [mhdlk-1:0] cryhplg9_24tqw;



  wire [mhdlk:0] uipdtjs;
  wire [mhdlk:0] acm0zbhvam;
  wire [mhdlk:0] oi40qurrxr; 
  wire [mhdlk:0] n89fv;

  wire jlo7_b_z = (irka0 ^ u22pp );
  assign oi40qurrxr = u22pp ? (n89fv << 1) : (n89fv >> 1);  

  ux607_gnrl_dfflrs #(1)  svv3sz17bdpp(jlo7_b_z, oi40qurrxr[0]   , n89fv[0]   , gf33atgy, ru_wi);
  ux607_gnrl_dfflr  #(mhdlk) o0mc8mg4cq9iqbw(jlo7_b_z, oi40qurrxr[mhdlk:1], n89fv[mhdlk:1], gf33atgy, ru_wi);


  assign uipdtjs = n89fv; 
  assign acm0zbhvam = (n89fv >> 1); 

  genvar i;
  generate 

    for (i=0; i<mhdlk; i=i+1) begin:eyoclcjcy41
      assign cryhplg9_24tqw[i] = u22pp & uipdtjs[i];      
      ux607_gnrl_dffl  #(onr7l) otz17hdw3zq3ny (cryhplg9_24tqw[i], qbjvs30wtb, olf4xmxku9u9k8[i], gf33atgy, ru_wi);
    end
  endgenerate


  integer j;
  reg [onr7l-1:0] ui9y38d1t;
  always @*
  begin : e82692n5bc4eh
    ui9y38d1t = {onr7l{1'b0}};
    for(j=0; j<mhdlk; j=j+1) begin
      ui9y38d1t = ui9y38d1t | ({onr7l{acm0zbhvam[j]}} & olf4xmxku9u9k8[j]);
    end
  end

  assign dqgck5s = ui9y38d1t;


endmodule 






















































module ux607_gnrl_0dffl # (
  parameter DW = 32
) (

  input               lden, 
  input      [DW-1:0] dnxt,
  output     [DW-1:0] qout,

  input               clk 
);

assign qout = dnxt;

endmodule






































module ux607_gnrl_dfflrs # (
  parameter DW = 32
) (

  input               lden, 
  input      [DW-1:0] dnxt,
  output     [DW-1:0] qout,

  input               clk,
  input               rst_n
);

reg [DW-1:0] qout_r;

always @(posedge clk or negedge rst_n)
begin : DFFLRS_PROC
  if (rst_n == 1'b0)
    qout_r <= {DW{1'b1}};
  else if (lden == 1'b1)
    qout_r <= dnxt;
end

assign qout = qout_r;



endmodule








module ux607_gnrl_dfflr # (
  parameter DW = 32
) (

  input               lden, 
  input      [DW-1:0] dnxt,
  output     [DW-1:0] qout,

  input               clk,
  input               rst_n
);

reg [DW-1:0] qout_r;

always @(posedge clk or negedge rst_n)
begin : DFFLR_PROC
  if (rst_n == 1'b0)
    qout_r <= {DW{1'b0}};
  else if (lden == 1'b1)
    qout_r <= dnxt;
end

assign qout = qout_r;



endmodule







module ux607_gnrl_dffl # (
  parameter DW = 32
) (

  input               lden, 
  input      [DW-1:0] dnxt,
  output     [DW-1:0] qout,

  input               clk,
  input               rst_n
);

reg [DW-1:0] qout_r;

always @(posedge clk or negedge rst_n)
begin : DFFLR_PROC
  if (rst_n == 1'b0)
    qout_r <= {DW{1'b0}};
  else if (lden == 1'b1)
    qout_r <= dnxt;
end







assign qout = qout_r;



endmodule








module ux607_gnrl_dffrs # (
  parameter DW = 32
) (

  input      [DW-1:0] dnxt,
  output     [DW-1:0] qout,

  input               clk,
  input               rst_n
);

reg [DW-1:0] qout_r;

always @(posedge clk or negedge rst_n)
begin : DFFRS_PROC
  if (rst_n == 1'b0)
    qout_r <= {DW{1'b1}};
  else                  
    qout_r <= dnxt;
end

assign qout = qout_r;

endmodule








module ux607_gnrl_dffr # (
  parameter DW = 32
) (

  input      [DW-1:0] dnxt,
  output     [DW-1:0] qout,

  input               clk,
  input               rst_n
);

reg [DW-1:0] qout_r;

always @(posedge clk or negedge rst_n)
begin : DFFR_PROC
  if (rst_n == 1'b0)
    qout_r <= {DW{1'b0}};
  else                  
    qout_r <= dnxt;
end

assign qout = qout_r;

endmodule











































































module dnxaqv6inphtvqkx85l8 # (
  parameter nm_fj = 32,
  parameter onr7l = 32,
  parameter h1b = 4,
  parameter o7hawonznex2 = 0,
  parameter cibz = 4,
  parameter s3xvyho = 1
) (
  input                         g4k11xiitgz962r,
  output                        nxfnmkeh2_oxuinwhs,
  input [nm_fj-1:0]                kez7oy1hkm0x_mba, 
  input                         czm7bw78q_ctanruda, 

  input                         r_zpoqtmqxzq_tli1, 

  input                         lqpb44qv17cgsfo8x,
  input                         kn1a55n2gcpb5fq,
  input                         yfqn924tp_05c,
  input                         qozylwb2v0y4igv8, 
  input [onr7l-1:0]                d6w6ulxl95ras8b4jl,
  input [h1b-1:0]                hdfxyj_9lnc9x9ls099,
  input [2:0]                   p6apzeecwtoem_e2x87,
  input [1:0]                   xmas5gu2txl3r66b1f,
  input                         ephj95nxeaa_zq,
  input                         mrpmr1jpfod77q,
  input [1:0]                   om7id6y4jtcq4,
  input [s3xvyho-1:0]             jq3nag_rg7k24ivb,
  input                         fl34njp9k3y4ar0ni,

  input                         wh6iy6zpdqsnv2y,
  output                        bd6yatp5cqq,
  output [cibz-1:0]             fl1qsvyu,
  output [nm_fj-1:0]               b9889wezsu,
  output [7:0]                  an__mxugc4,
  output [2:0]                  poj6g8vw9e,
  output [1:0]                  dafaivw3ze9g3hi,
  output [1:0]                  q2c0d6fxz_1bw,
  output [3:0]                  wblesminvapwua,
  output [2:0]                  v3cim36gj8g,
  output [3:0]                  ss22f8fuy2uhr,
  output [3:0]                  hoaoalj5pcdnpnm0,
  output [s3xvyho-1:0]            rh8f1e3jgg3xi,

  input                         su81e8dxdzng9d,

  input                         gf33atgy,
  input                         ru_wi
  );

  localparam lz4sj516 = cibz+nm_fj+8+3+2+2+4+3+4+4+s3xvyho;

  wire              jjzyws5k2y;
  wire [cibz-1:0]   oxg_62rd;
  wire [nm_fj-1:0]     t81yn8tjj3w9;
  wire [7:0]        vs54w5c2ooj;
  wire [2:0]        uzx7w674;
  wire [1:0]        dumrm6jjys;
  wire [1:0]        zb6d1sdg8;
  wire [3:0]        xrownimt0;
  wire [2:0]        bswkrhnbw48;
  wire [3:0]        ktm0lkro5_o;
  wire [3:0]        ehwfq189_ihl;
  wire [s3xvyho-1:0]  b1flhed5odia;

  wire [lz4sj516-1:0] df5moo3d13q4u;
  wire [lz4sj516-1:0] g4w1yi_zyhgm3ge;
  wire q53bqe63zmc;
  wire v4_z18v6rk;
  wire foqp7o_7fw4;
  wire oqz8s2vautyzl;

  wire gsah_6u4uzun7es;
  wire kdpm897dm7ouma;
  wire lsujd2xqfcpvjp;
  wire n7uomqy4ff238cfij1q;
  wire erg1ck3i657tivpvo;

  assign lsujd2xqfcpvjp = n7uomqy4ff238cfij1q || erg1ck3i657tivpvo;

  assign gsah_6u4uzun7es = wh6iy6zpdqsnv2y;


  generate
    if (o7hawonznex2 == 0) begin :t2uoqogn_6otbq02avby
  assign kdpm897dm7ouma   = 1'b0;
  assign n7uomqy4ff238cfij1q = 1'b0;
  assign erg1ck3i657tivpvo = 1'b0;
    end
    else begin :ib9gmgog8cyk6zc7qyxc8
  assign n7uomqy4ff238cfij1q = nxfnmkeh2_oxuinwhs && g4k11xiitgz962r && xmas5gu2txl3r66b1f[0];
  assign erg1ck3i657tivpvo = kdpm897dm7ouma && nxfnmkeh2_oxuinwhs && g4k11xiitgz962r && xmas5gu2txl3r66b1f[1];
  ux607_gnrl_dfflr #(1) gt_e9bu3kwaow1wwznyl (lsujd2xqfcpvjp, n7uomqy4ff238cfij1q, kdpm897dm7ouma, gf33atgy, ru_wi);
    end
  endgenerate

  assign nxfnmkeh2_oxuinwhs = v4_z18v6rk | kdpm897dm7ouma;

  assign jjzyws5k2y = g4k11xiitgz962r & (~kdpm897dm7ouma);

  assign oxg_62rd     = {cibz{1'b0}};
  assign t81yn8tjj3w9   = kez7oy1hkm0x_mba;
  generate
    if (onr7l == 32) begin :ni_mx7tf3elt
  assign vs54w5c2ooj = (p6apzeecwtoem_e2x87 == 3'b0) ? 8'b0 : 8'b00000111;
    end
    else begin :vm69kdoyqgi12
  assign vs54w5c2ooj = (p6apzeecwtoem_e2x87 == 3'b0) ? 8'b0 : 8'b00000011;
    end
  endgenerate

  assign uzx7w674    = {1'b0,om7id6y4jtcq4};
  assign dumrm6jjys   = p6apzeecwtoem_e2x87[1:0];
  assign zb6d1sdg8    = {ephj95nxeaa_zq,mrpmr1jpfod77q}; 
  assign xrownimt0   =  kn1a55n2gcpb5fq ? 4'b0000 :
                        yfqn924tp_05c     ? 4'b0010 : 4'b1111;

  assign bswkrhnbw48[0] = czm7bw78q_ctanruda | r_zpoqtmqxzq_tli1;



  assign bswkrhnbw48[1] = 1'b0; 
  assign bswkrhnbw48[2] = fl34njp9k3y4ar0ni;
  assign ktm0lkro5_o     = 4'b0;
  assign ehwfq189_ihl  = 4'b0;
  assign b1flhed5odia    = jq3nag_rg7k24ivb;

  assign df5moo3d13q4u = 
                      {
                        oxg_62rd,
                        t81yn8tjj3w9,
                        vs54w5c2ooj,
                        uzx7w674,
                        dumrm6jjys,
                        zb6d1sdg8,
                        xrownimt0,
                        bswkrhnbw48,
                        ktm0lkro5_o,
                        ehwfq189_ihl,
                        b1flhed5odia 
                      };
  assign {
           fl1qsvyu,
           b9889wezsu,
           an__mxugc4,
           poj6g8vw9e,
           dafaivw3ze9g3hi,
           q2c0d6fxz_1bw,
           wblesminvapwua,
           v3cim36gj8g,
           ss22f8fuy2uhr,
           hoaoalj5pcdnpnm0,
           rh8f1e3jgg3xi 
         } = g4w1yi_zyhgm3ge;
  assign bd6yatp5cqq = foqp7o_7fw4;

  assign q53bqe63zmc = jjzyws5k2y;

  assign oqz8s2vautyzl = gsah_6u4uzun7es;

  vq28fpkbg0dxljs8bf0k # (
        .hejad2_b4dywimoxw5 (0),
        .evi4vkasjp742kf4 (1),
        .mhdlk  (2),
        .onr7l  (lz4sj516)
  ) aprrbyg85wsud_3ri_ (
        .geml8twgru(1'b1),
        .bw6ftrau0(q53bqe63zmc),
        .eef2g8(v4_z18v6rk),
        .qbjvs30wtb(df5moo3d13q4u),

        .td5hjljc_(su81e8dxdzng9d),
        .wqljp(foqp7o_7fw4),
        .h9378(oqz8s2vautyzl),  
        .dqgck5s(g4w1yi_zyhgm3ge),  

        .i0lklnhw28rc7dj(),
        .gf33atgy  (gf33atgy),
        .ru_wi(ru_wi)
  );

endmodule








module serhetfxiy9lcu5155j03mqqa # (
  parameter nm_fj = 32,
  parameter onr7l = 32,
  parameter h1b = 4,
  parameter o7hawonznex2 = 0,
  parameter cibz = 4,
  parameter s3xvyho = 1
) (
  input                         v5brbv_o0cwz8ltkbnv,
  output                        h6vhmpdy12279cq0xb6,
  input [nm_fj-1:0]                zh16cx29t0l33, 
  input                         f14hyggy6ln5pyn, 

  input                         a_bzkj6xlfrxcts, 

  input                         rbd2kwb5sl2qjjspc_3,
  input                         xij68avnrqqthb23rwq9,
  input                         trqijdd7kcw97e,
  input                         kg6c6siv37bjp1, 
  input [onr7l-1:0]                ka4nz5iwhho4_t,
  input [h1b-1:0]                fzedypimn06pveo8,
  input [2:0]                   gsh3nost5unqiaqgo,
  input [1:0]                   ld9htofs52b7nj,
  input                         tzhgbyplxl9mi,
  input                         f22pg5kqjpfmk83h2e,
  input [1:0]                   iwvo07en81_3rvne,
  input [s3xvyho-1:0]             hi_0bv4ttpvt3lv,

  input                         roral7fym4h3_,
  output                        b_gwvq35iq0_yvk,
  output [cibz-1:0]             lqm2hm0cjm5zt,
  output [nm_fj-1:0]               f3n3tpjs44e0_,
  output [7:0]                  dmc59hxf352z,
  output [2:0]                  a63l3og_8qak5jy,
  output [1:0]                  m0wp58qmji79,
  output [1:0]                  c8qmnfk1vqai,
  output [3:0]                  pbov8g9yizcwr,
  output [2:0]                  t8qjehupeajtzjr,
  output [3:0]                  hhp1rh0x0jn,
  output [3:0]                  w9yptl69xj6p,
  output [s3xvyho-1:0]            yvcpy_gyehs4lji, 

  input                         kted7ph0krq,
  output                        a93i3d2hji,
  output [cibz-1:0]             of5p5cb8p4,
  output [onr7l-1:0]               g1bi1xzuv64,
  output [h1b-1:0]               gj6p5b5ik3r9p,
  output                        m1fmaas4oww6,

  input                         su81e8dxdzng9d,

  input                         gf33atgy,
  input                         ru_wi
  );

  localparam z_zas5vxa9tm6 = cibz+nm_fj+8+3+2+2+4+3+4+4+s3xvyho;
  localparam vbin99rg = cibz+onr7l+h1b+1;

  wire veevjhsee4m1xr;
  wire ylzs7afax46fexip;
  wire kdpm897dm7ouma;
  wire lsujd2xqfcpvjp;
  wire n7uomqy4ff238cfij1q;
  wire erg1ck3i657tivpvo;






  wire [z_zas5vxa9tm6-1:0] gov0_o3355d7n;
  wire [z_zas5vxa9tm6-1:0] hqlf5lb77a_5_ljzv;
  wire [vbin99rg-1:0] rtjg74o29s8vna;
  wire [vbin99rg-1:0] cekagfs42vmj;
  wire swl1m6fogsw6ozr;
  wire qsuolgu9fsxyy6p;
  wire xqw4n7_2r8xe;
  wire fuupnrnlzj9d;
  wire dp9oloqrkupwlc2m;
  wire wa1no6q55zwv3wdz;
  wire o7clr1w1aiy6g;
  wire iia1yvb0gyr00;

  wire                voiq2spycj_;
  wire                odpkxjfem7a;
  wire [cibz-1:0]     ascpf2;
  wire [nm_fj-1:0]       ii_lw9ywmoc;
  wire [7:0]          ns_iou4i4pr;
  wire [2:0]          yrwy90nlljfg3;
  wire [1:0]          yfm2n751el84;
  wire [1:0]          blffjrtqe;
  wire [3:0]          izcefcjcun;
  wire [2:0]          s_iwmvhkrn;
  wire [3:0]          rgaxv89;
  wire [3:0]          d92rp7q081s4qxk;
  wire [s3xvyho-1:0]    htp29e1v4nj1; 

  wire                c4yb_u8p;
  wire                ht9pk4ei10i96;
  wire [cibz-1:0]     d8ffhz;
  wire [onr7l-1:0]       d89w_0uizmen;
  wire [h1b-1:0]       bzjc7dm;
  wire                abfk9hyf2;

  assign veevjhsee4m1xr = roral7fym4h3_ ;
  assign ylzs7afax46fexip  = kted7ph0krq  ;

  assign gov0_o3355d7n = 
                      {
                        ascpf2,
                        ii_lw9ywmoc,
                        ns_iou4i4pr,
                        yrwy90nlljfg3,
                        yfm2n751el84,
                        blffjrtqe,
                        izcefcjcun,
                        s_iwmvhkrn,
                        rgaxv89,
                        d92rp7q081s4qxk,
                        htp29e1v4nj1  
                      };
  assign swl1m6fogsw6ozr = odpkxjfem7a;
  assign voiq2spycj_ = qsuolgu9fsxyy6p; 
  assign {
          lqm2hm0cjm5zt,
          f3n3tpjs44e0_,
          dmc59hxf352z,
          a63l3og_8qak5jy,
          m0wp58qmji79,
          c8qmnfk1vqai,
          pbov8g9yizcwr,
          t8qjehupeajtzjr,
          hhp1rh0x0jn,
          w9yptl69xj6p,
          yvcpy_gyehs4lji  
         } = hqlf5lb77a_5_ljzv;
  assign b_gwvq35iq0_yvk = xqw4n7_2r8xe;
  assign fuupnrnlzj9d = veevjhsee4m1xr;

  assign rtjg74o29s8vna = 
                      {
                       d8ffhz,
                       d89w_0uizmen,
                       bzjc7dm,
                       abfk9hyf2
                      };
  assign dp9oloqrkupwlc2m = ht9pk4ei10i96;
  assign c4yb_u8p    = wa1no6q55zwv3wdz; 
  assign {
          of5p5cb8p4,
          g1bi1xzuv64,
          gj6p5b5ik3r9p,
          m1fmaas4oww6
         } = cekagfs42vmj;

  assign a93i3d2hji  = o7clr1w1aiy6g;
  assign iia1yvb0gyr00 = ylzs7afax46fexip;

  vq28fpkbg0dxljs8bf0k # (
        .hejad2_b4dywimoxw5 (0),
        .evi4vkasjp742kf4 (1),
        .mhdlk  (2),
        .onr7l  (z_zas5vxa9tm6)
  ) mv67njo098wtgffd (
        .geml8twgru(1'b1),
        .bw6ftrau0(swl1m6fogsw6ozr),
        .eef2g8(qsuolgu9fsxyy6p),
        .qbjvs30wtb(gov0_o3355d7n),

        .td5hjljc_(su81e8dxdzng9d),
        .wqljp(xqw4n7_2r8xe),
        .h9378(fuupnrnlzj9d),  
        .dqgck5s(hqlf5lb77a_5_ljzv),  

        .i0lklnhw28rc7dj(),
        .gf33atgy  (gf33atgy),
        .ru_wi(ru_wi)
  );

  vq28fpkbg0dxljs8bf0k # (
        .hejad2_b4dywimoxw5 (0),
        .evi4vkasjp742kf4 (1),
        .mhdlk  (2),
        .onr7l  (vbin99rg)
  ) jfz87di8otj6 (
        .geml8twgru(1'b1),
        .bw6ftrau0(dp9oloqrkupwlc2m),
        .eef2g8(wa1no6q55zwv3wdz),
        .qbjvs30wtb(rtjg74o29s8vna),

        .td5hjljc_(su81e8dxdzng9d),
        .wqljp(o7clr1w1aiy6g),
        .h9378(iia1yvb0gyr00),  
        .dqgck5s(cekagfs42vmj),  

        .i0lklnhw28rc7dj(),
        .gf33atgy  (gf33atgy),
        .ru_wi(ru_wi)
  );

  assign lsujd2xqfcpvjp = n7uomqy4ff238cfij1q || erg1ck3i657tivpvo;


  generate
    if (o7hawonznex2 == 0) begin :t2uoqogn_6otbq02avby
  assign kdpm897dm7ouma   = 1'b0;
  assign n7uomqy4ff238cfij1q = 1'b0;
  assign erg1ck3i657tivpvo = 1'b0;
    end
    else begin :ib9gmgog8cyk6zc7qyxc8
  assign n7uomqy4ff238cfij1q = h6vhmpdy12279cq0xb6 && v5brbv_o0cwz8ltkbnv && ld9htofs52b7nj[0];
  assign erg1ck3i657tivpvo = kdpm897dm7ouma && h6vhmpdy12279cq0xb6 && v5brbv_o0cwz8ltkbnv && ld9htofs52b7nj[1];
  ux607_gnrl_dfflr #(1) gt_e9bu3kwaow1wwznyl (lsujd2xqfcpvjp, n7uomqy4ff238cfij1q, kdpm897dm7ouma, gf33atgy, ru_wi);
    end
  endgenerate

  assign h6vhmpdy12279cq0xb6 =   (voiq2spycj_ || kdpm897dm7ouma) && (c4yb_u8p);
  assign odpkxjfem7a = v5brbv_o0cwz8ltkbnv && (!kdpm897dm7ouma) && c4yb_u8p;
  assign ht9pk4ei10i96  = v5brbv_o0cwz8ltkbnv && (voiq2spycj_ || kdpm897dm7ouma);

  assign ascpf2     = {cibz{1'b0}};
  assign ii_lw9ywmoc   = zh16cx29t0l33;
  generate
    if (onr7l == 32) begin :vhk2cd6mozpn7
  assign ns_iou4i4pr = (gsh3nost5unqiaqgo == 3'b0) ? 8'b0 : 8'b00000111;
    end
    else begin :aaqzj21gbcv
  assign ns_iou4i4pr = (gsh3nost5unqiaqgo == 3'b0) ? 8'b0 : 8'b00000011;
    end
  endgenerate

  assign yrwy90nlljfg3    = {1'b0,iwvo07en81_3rvne};
  assign yfm2n751el84   = gsh3nost5unqiaqgo[1:0];
  assign blffjrtqe    = {tzhgbyplxl9mi,f22pg5kqjpfmk83h2e}; 
  assign izcefcjcun   =  xij68avnrqqthb23rwq9 ? 4'b0000 :
                        trqijdd7kcw97e     ? 4'b0010 : 4'b1111;

  assign s_iwmvhkrn[0] = f14hyggy6ln5pyn | a_bzkj6xlfrxcts;



  assign s_iwmvhkrn[1] = 1'b0; 
  assign s_iwmvhkrn[2] = 1'b0;
  assign rgaxv89     = 4'b0;
  assign d92rp7q081s4qxk  = 4'b0;
  assign htp29e1v4nj1    = hi_0bv4ttpvt3lv;

  assign d8ffhz       = {cibz{1'b0}};
  assign d89w_0uizmen     = ka4nz5iwhho4_t;
  assign bzjc7dm     = fzedypimn06pveo8;   
  assign abfk9hyf2    = ((ld9htofs52b7nj == 2'b00) && !kdpm897dm7ouma) || ld9htofs52b7nj[1];
endmodule








module ux607_gnrl_icb2axi_r # (
  parameter AW = 32,
  parameter DW = 32,
  parameter MW = 4,
  parameter ALLOW_BURST = 0,
  parameter ID_W = 4
) (
  output                         icb_rrsp_valid,
  input                          icb_rrsp_ready,
  output [DW-1:0]                icb_rrsp_rdata,
  output                         icb_rrsp_err,
  output                         icb_rrsp_excl_ok,
  output                         icb_rrsp_rlast,

  output                         axi_rready,
  input                          axi_rvalid,
  input [ID_W-1:0]               axi_rid,
  input [DW-1:0]                 axi_rdata,
  input [1:0]                    axi_rresp,
  input                          axi_rlast,

  input                         axi_bus_clk_en,



  input                         clk,
  input                         rst_n
  );

  localparam lz4sj516 = ID_W+DW+2+1;
  wire                          ximmd6ve7;
  wire [ID_W-1:0]               nm3kvsg;
  wire [DW-1:0]                 f6uxao0sgpg;
  wire [1:0]                    jq10segu8__;
  wire                          nov_dsjah;

  wire [lz4sj516-1:0] df5moo3d13q4u;
  wire [lz4sj516-1:0] g4w1yi_zyhgm3ge;
  wire q53bqe63zmc;
  wire v4_z18v6rk;
  wire foqp7o_7fw4;
  wire oqz8s2vautyzl;

  assign df5moo3d13q4u = 
                      {
                        axi_rid,
                        axi_rdata,
                        axi_rresp,
                        axi_rlast 
                      };
  assign {
          nm3kvsg,
          f6uxao0sgpg,
          jq10segu8__,
          nov_dsjah 
         } = g4w1yi_zyhgm3ge;

  assign ximmd6ve7 = foqp7o_7fw4;

  assign q53bqe63zmc = axi_rvalid ;
  assign axi_rready = v4_z18v6rk;

  assign oqz8s2vautyzl = icb_rrsp_ready;

  vq28fpkbg0dxljs8bf0k # (
        .hejad2_b4dywimoxw5 (1),
        .evi4vkasjp742kf4 (0),
        .mhdlk  (2),
        .onr7l  (lz4sj516)
  ) q35nsujqlr5e2ql (
        .geml8twgru(axi_bus_clk_en),
        .bw6ftrau0(q53bqe63zmc),
        .eef2g8(v4_z18v6rk),
        .qbjvs30wtb(df5moo3d13q4u),

        .td5hjljc_(1'b1),
        .wqljp(foqp7o_7fw4),
        .h9378(oqz8s2vautyzl),  
        .dqgck5s(g4w1yi_zyhgm3ge),  

        .i0lklnhw28rc7dj(),
        .gf33atgy  (clk),
        .ru_wi(rst_n)
  );

  assign icb_rrsp_valid   = ximmd6ve7;

  assign icb_rrsp_err     = jq10segu8__[1] ; 
  assign icb_rrsp_excl_ok = (jq10segu8__ == 2'b01);
  assign icb_rrsp_rdata   = f6uxao0sgpg;
  assign icb_rrsp_rlast   = nov_dsjah;
endmodule








module ux607_gnrl_icb2axi_b # (
  parameter AW = 32,
  parameter DW = 32,
  parameter MW = 4,
  parameter ALLOW_BURST = 0,
  parameter ID_W = 4
) (
  output                         icb_wrsp_valid,
  input                          icb_wrsp_ready,
  output                         icb_wrsp_err,
  output                         icb_wrsp_excl_ok,
  output                         icb_wrsp_last,

  output                         axi_bready,
  input                          axi_bvalid,
  input [ID_W-1:0]               axi_bid,
  input [1:0]                    axi_bresp,

  input                         axi_bus_clk_en,

  input                         wrsp_burst, 
  input                         wrsp_excl,  

  input                         clk,
  input                         rst_n
  );

  localparam lz4sj516 = ID_W+2+1;
  wire                          zbto07id9kb;
  wire [ID_W-1:0]               i_fsr;
  wire [1:0]                    d2ip29ji1;
  wire                          i1ovoiv;

  wire [lz4sj516-1:0] df5moo3d13q4u;
  wire [lz4sj516-1:0] g4w1yi_zyhgm3ge;
  wire q53bqe63zmc;
  wire v4_z18v6rk;
  wire foqp7o_7fw4;
  wire oqz8s2vautyzl;

  wire       afkj5yhhtctg6s;
  wire [2:0] g85wmlhjsfg_;
  wire [2:0] qv6grfmv4g0b663;
  wire       d767w05jxusx0gx6;

  assign df5moo3d13q4u = 
                      {
                        axi_bid,
                        axi_bresp,
                        wrsp_burst
                      };
  assign {
          i_fsr,
          d2ip29ji1,
          i1ovoiv
         } = g4w1yi_zyhgm3ge;

  assign zbto07id9kb = foqp7o_7fw4;

  assign q53bqe63zmc = axi_bvalid ;
  assign axi_bready = v4_z18v6rk;

  assign oqz8s2vautyzl = icb_wrsp_ready && (!i1ovoiv || afkj5yhhtctg6s);

  vq28fpkbg0dxljs8bf0k # (
        .hejad2_b4dywimoxw5 (1),
        .evi4vkasjp742kf4 (0),
        .mhdlk  (2),
        .onr7l  (lz4sj516)
  ) q037u7vw0lyuh8 (
        .geml8twgru(axi_bus_clk_en),
        .bw6ftrau0(q53bqe63zmc),
        .eef2g8(v4_z18v6rk),
        .qbjvs30wtb(df5moo3d13q4u),

        .td5hjljc_(1'b1),
        .wqljp(foqp7o_7fw4),
        .h9378(oqz8s2vautyzl),  
        .dqgck5s(g4w1yi_zyhgm3ge),  

        .i0lklnhw28rc7dj(),
        .gf33atgy  (clk),
        .ru_wi(rst_n)
  );

  generate
    if (ALLOW_BURST == 0) begin :bd14fahfursl
  assign afkj5yhhtctg6s =1'b0;
  assign g85wmlhjsfg_ = 3'b0;
  assign qv6grfmv4g0b663 = 3'b0;
  assign d767w05jxusx0gx6 = 1'b0;
    end
    else begin :j_7fmjdgwqmy5
  assign qv6grfmv4g0b663 = afkj5yhhtctg6s ? 3'b0 : (g85wmlhjsfg_ + 3'b1);
  assign afkj5yhhtctg6s = ((DW==32) && (g85wmlhjsfg_==3'b111)) || ((DW==64) && (g85wmlhjsfg_==3'b011));
  assign d767w05jxusx0gx6 = i1ovoiv && icb_wrsp_valid && icb_wrsp_ready;
  ux607_gnrl_dfflr #(3) azqo5a_gl8snymahf0 (d767w05jxusx0gx6, qv6grfmv4g0b663, g85wmlhjsfg_, clk, rst_n);
    end
  endgenerate

  assign icb_wrsp_valid   = zbto07id9kb;
  assign icb_wrsp_err     = d2ip29ji1[1] || ((d2ip29ji1 == 2'b01) && !wrsp_excl);
  assign icb_wrsp_excl_ok = wrsp_excl && (d2ip29ji1 == 2'b01);
  assign icb_wrsp_last    = afkj5yhhtctg6s;
endmodule



module w17x4i82vejgdgfxy6 # (
  parameter nm_fj = 32,
  parameter onr7l = 32,
  parameter h1b = 4,
  parameter o7hawonznex2 = 0,
  parameter cibz = 4,
  parameter s3xvyho = 1
  ) (

  input                         wh6iy6zpdqsnv2y,
  output                        bd6yatp5cqq,
  output [cibz-1:0]             fl1qsvyu,
  output [nm_fj-1:0]               b9889wezsu,
  output [7:0]                  an__mxugc4,
  output [2:0]                  poj6g8vw9e,
  output [1:0]                  dafaivw3ze9g3hi,
  output [1:0]                  q2c0d6fxz_1bw,
  output [3:0]                  wblesminvapwua,
  output [2:0]                  v3cim36gj8g,
  output [3:0]                  ss22f8fuy2uhr,
  output [3:0]                  hoaoalj5pcdnpnm0,
  output [s3xvyho-1:0]            rh8f1e3jgg3xi,

  output                        hjstsi51gm,
  input                         onpqhy0s69,
  input [cibz-1:0]              aw7xjbi,
  input [onr7l-1:0]                z0cc2y_uzoh_,
  input [1:0]                   y8tc_vywu82ugn,
  input                         o2h9d51o6m6,

  input                         su81e8dxdzng9d,

  input                         b0o3_z1qhzguxuvx03v93gz,
  output                        tslw7f9ona4tph8dm0nt,
  input [nm_fj-1:0]                y2wr5gyopdnthewqrxe7, 
  input                         zlz5s0ait6hwykg4b, 
  input [onr7l-1:0]                v2se1vid1uml27uvf2t4yli,
  input [h1b-1:0]                g8ttk2wz9kvwdwkzp5kwp,
  input [2:0]                   h4a4okoossdfjraixe2sl,
  input [1:0]                   tnppka2a6z82_mietistn,
  input                         tsjfjoan2dw95g05__g5q,
  input                         hy9p1vxnb29wsf43qczd,
  input [1:0]                   zefzgdtbg9u39vfb3,
  input                         hnnr5of3orcsqxyfb86ma,

  input                         jl91z78pj9nm0rbl3t7www6,

  input                         wjtoelq31c7h13gu_yhskwl,
  input                         x_6hf7jugp8hwgu0j10t1,
  input                         t6f_omqkgrkzy903,
  input                         obdyu6w0wqx4b3g8t,

  output                        yk58l7ldat5ahcp4j1i,
  input                         e8h0j_anz7mzuobmbwzv8g,
  output                        uebzayybqiyy1cicc  ,
  output                        afb8snj62vkl7pacmyj3,
  output [onr7l-1:0]               zuv8v13fabr90783u1lc0,

  input                         gf33atgy,
  input                         ru_wi
  );

  wire s6rovfnjby0xp0yy19abab_;

























  dnxaqv6inphtvqkx85l8 # (
            .nm_fj (nm_fj),
            .onr7l (onr7l),
            .h1b (h1b),
            .o7hawonznex2(o7hawonznex2),
            .cibz (cibz),
            .s3xvyho (s3xvyho)
) d6q08tysboaij8mmzpz9t(
            .g4k11xiitgz962r (b0o3_z1qhzguxuvx03v93gz),
            .nxfnmkeh2_oxuinwhs (tslw7f9ona4tph8dm0nt),
            .kez7oy1hkm0x_mba (y2wr5gyopdnthewqrxe7), 
            .czm7bw78q_ctanruda (hnnr5of3orcsqxyfb86ma), 

            .r_zpoqtmqxzq_tli1 (jl91z78pj9nm0rbl3t7www6), 

            .lqpb44qv17cgsfo8x (wjtoelq31c7h13gu_yhskwl),
            .kn1a55n2gcpb5fq (x_6hf7jugp8hwgu0j10t1),
            .yfqn924tp_05c (t6f_omqkgrkzy903),
            .qozylwb2v0y4igv8 (zlz5s0ait6hwykg4b), 
            .d6w6ulxl95ras8b4jl (v2se1vid1uml27uvf2t4yli),
            .hdfxyj_9lnc9x9ls099 (g8ttk2wz9kvwdwkzp5kwp),
            .p6apzeecwtoem_e2x87 (h4a4okoossdfjraixe2sl),
            .xmas5gu2txl3r66b1f (tnppka2a6z82_mietistn),
            .ephj95nxeaa_zq (tsjfjoan2dw95g05__g5q),
            .mrpmr1jpfod77q (hy9p1vxnb29wsf43qczd),
            .om7id6y4jtcq4 (zefzgdtbg9u39vfb3),
            .jq3nag_rg7k24ivb ({s3xvyho{1'b0}}),
            .fl34njp9k3y4ar0ni (obdyu6w0wqx4b3g8t),

            .wh6iy6zpdqsnv2y (wh6iy6zpdqsnv2y),
            .bd6yatp5cqq (bd6yatp5cqq),
            .fl1qsvyu (fl1qsvyu),
            .b9889wezsu (b9889wezsu),
            .an__mxugc4 (an__mxugc4),
            .poj6g8vw9e (poj6g8vw9e),
            .dafaivw3ze9g3hi (dafaivw3ze9g3hi),
            .q2c0d6fxz_1bw (q2c0d6fxz_1bw),
            .wblesminvapwua (wblesminvapwua),
            .v3cim36gj8g (v3cim36gj8g),
            .ss22f8fuy2uhr (ss22f8fuy2uhr),
            .hoaoalj5pcdnpnm0 (hoaoalj5pcdnpnm0),
            .rh8f1e3jgg3xi (rh8f1e3jgg3xi),

            .su81e8dxdzng9d (su81e8dxdzng9d),

            .gf33atgy (gf33atgy),
            .ru_wi (ru_wi)
  );

  ux607_gnrl_icb2axi_r # (
            .AW (nm_fj),
            .DW (onr7l),
            .MW (h1b),
            .ALLOW_BURST(o7hawonznex2),
            .ID_W (cibz) 
  ) mgts9zfavjfv(
            .icb_rrsp_valid (yk58l7ldat5ahcp4j1i),
            .icb_rrsp_ready (e8h0j_anz7mzuobmbwzv8g),
            .icb_rrsp_rdata (zuv8v13fabr90783u1lc0),
            .icb_rrsp_err (uebzayybqiyy1cicc),
            .icb_rrsp_rlast  (s6rovfnjby0xp0yy19abab_),
            .icb_rrsp_excl_ok (afb8snj62vkl7pacmyj3),

            .axi_rready (hjstsi51gm),
            .axi_rvalid (onpqhy0s69),
            .axi_rid (aw7xjbi),
            .axi_rdata (z0cc2y_uzoh_),
            .axi_rresp (y8tc_vywu82ugn),
            .axi_rlast (o2h9d51o6m6),

            .axi_bus_clk_en (su81e8dxdzng9d),



            .clk (gf33atgy),
            .rst_n (ru_wi)
  );
endmodule




module o0kamfqxkze9obdxf3 #(
  parameter nm_fj = 32,
  parameter onr7l = 32,
  parameter h1b = 4,
  parameter o7hawonznex2 = 0,
  parameter n9z24gbmpt_t =4,
  parameter cibz = 4,
  parameter s3xvyho = 1
) (

  input                         roral7fym4h3_,
  output                        b_gwvq35iq0_yvk,
  output [cibz-1:0]             lqm2hm0cjm5zt,
  output [nm_fj-1:0]               f3n3tpjs44e0_,
  output [7:0]                  dmc59hxf352z,
  output [2:0]                  a63l3og_8qak5jy,
  output [1:0]                  m0wp58qmji79,
  output [1:0]                  c8qmnfk1vqai,
  output [3:0]                  pbov8g9yizcwr,
  output [2:0]                  t8qjehupeajtzjr,
  output [3:0]                  hhp1rh0x0jn,
  output [3:0]                  w9yptl69xj6p,
  output [s3xvyho-1:0]            yvcpy_gyehs4lji, 

  input                         kted7ph0krq,
  output                        a93i3d2hji,
  output [cibz-1:0]             of5p5cb8p4,
  output [onr7l-1:0]               g1bi1xzuv64,
  output [h1b-1:0]               gj6p5b5ik3r9p,
  output                        m1fmaas4oww6,

  output                         nneek3ep5xykwl,
  input                          g8khua4l0y77zjp,
  input [cibz-1:0]                wmlp1a2b,
  input [1:0]                    weop50xb_avne,

  input                         su81e8dxdzng9d,

  input                         vzikn9_n0lvrdaomdo5ys,
  output                        n1_vj412ga534kpmgnc7,
  input [nm_fj-1:0]                ksjpl34uepyev0_db5ejr,
  input                         xzlaan0xyx3f5eo20zoo, 
  input [onr7l-1:0]                ww86vetlr_66ts64yhf00,
  input [h1b-1:0]                w76w2dx5nq4zgy_xsa5,
  input [2:0]                   l4eydle02q0gt8sp79xmpj,
  input [1:0]                   u5iq9uuj_lmerh15q8z,
  input                         emsvw7kp7xfm9g5s5y,
  input                         w99a9y3nh8ju8d3ns6jr,
  input [1:0]                   t7rgyydfts3enyenh,
  input                         iwmw44ethjx3dsud0egh,

  input                         l2hjyz8uo5ft9i_3d_,

  input                         ji71tydckvigh3o__p24_m,
  input                         cugxuq_z5o_cojyelhop2,
  input                         ypof75b4bl9g4e_an,

  output                        sg96uazxf6dpizg7vad,
  input                         qe9rerwzfqnxm49kvj69u,
  output                        ba1jgqojkjt_p5wrx1x,
  output                        jgvpcfglnc5lptyi2ca5hkmuv,

  input                         gf33atgy,
  input                         ru_wi
  );



  wire slggcmvgdj;
  wire homm_w8zq;
  wire r8aazdlqr6;
  wire cpspx16gnkw9rv;
  wire zfph1n2fv95oalqawi;
  wire yuwam57krt02tnm8;
  generate
  wire edjq61okne5m2wnwpj4in9;
  assign zfph1n2fv95oalqawi   = b_gwvq35iq0_yvk && roral7fym4h3_;
if (o7hawonznex2 == 1) begin :gq_djhm1ocjq7gp25rij
  assign r8aazdlqr6       = (dmc59hxf352z != 0);
end
else begin :gqoo4lhnmi6vu0cr0
  assign r8aazdlqr6       = 1'b0;
end
endgenerate
  assign cpspx16gnkw9rv        = c8qmnfk1vqai[0];
  assign yuwam57krt02tnm8 = g8khua4l0y77zjp && nneek3ep5xykwl;
  vq28fpkbg0dxljs8bf0k # (
        .hejad2_b4dywimoxw5 (1),
        .evi4vkasjp742kf4 (1),
        .mhdlk  (n9z24gbmpt_t),
        .onr7l  (2)
  ) ha_de4p5a0a9xfv9 (

        .geml8twgru(su81e8dxdzng9d),
        .bw6ftrau0(zfph1n2fv95oalqawi),
        .eef2g8(),
        .qbjvs30wtb({r8aazdlqr6,cpspx16gnkw9rv}),

        .td5hjljc_(su81e8dxdzng9d),
        .wqljp(),
        .h9378(yuwam57krt02tnm8),  
        .dqgck5s({slggcmvgdj,homm_w8zq}),  

        .i0lklnhw28rc7dj(),
        .gf33atgy  (gf33atgy),
        .ru_wi(ru_wi)
  );

  serhetfxiy9lcu5155j03mqqa # (
            .nm_fj (nm_fj),
            .onr7l (onr7l),
            .h1b (h1b),
            .o7hawonznex2(o7hawonznex2),
            .cibz (cibz),
            .s3xvyho (s3xvyho)
) yq2i083ywp2ki_6x82 (
            .v5brbv_o0cwz8ltkbnv (vzikn9_n0lvrdaomdo5ys),
            .h6vhmpdy12279cq0xb6 (n1_vj412ga534kpmgnc7),
            .zh16cx29t0l33 (ksjpl34uepyev0_db5ejr), 
            .f14hyggy6ln5pyn (iwmw44ethjx3dsud0egh), 

            .a_bzkj6xlfrxcts (l2hjyz8uo5ft9i_3d_), 

            .rbd2kwb5sl2qjjspc_3 (ji71tydckvigh3o__p24_m),
            .xij68avnrqqthb23rwq9 (cugxuq_z5o_cojyelhop2),
            .trqijdd7kcw97e (ypof75b4bl9g4e_an),
            .kg6c6siv37bjp1 (xzlaan0xyx3f5eo20zoo), 
            .ka4nz5iwhho4_t (ww86vetlr_66ts64yhf00),
            .fzedypimn06pveo8 (w76w2dx5nq4zgy_xsa5),
            .gsh3nost5unqiaqgo (l4eydle02q0gt8sp79xmpj),
            .ld9htofs52b7nj (u5iq9uuj_lmerh15q8z),
            .tzhgbyplxl9mi (emsvw7kp7xfm9g5s5y),
            .f22pg5kqjpfmk83h2e (w99a9y3nh8ju8d3ns6jr),
            .iwvo07en81_3rvne (t7rgyydfts3enyenh),
            .hi_0bv4ttpvt3lv ({s3xvyho{1'b0}}),

            .roral7fym4h3_ (roral7fym4h3_),
            .b_gwvq35iq0_yvk (b_gwvq35iq0_yvk),
            .lqm2hm0cjm5zt (lqm2hm0cjm5zt),
            .f3n3tpjs44e0_ (f3n3tpjs44e0_),
            .dmc59hxf352z (dmc59hxf352z),
            .a63l3og_8qak5jy (a63l3og_8qak5jy),
            .m0wp58qmji79 (m0wp58qmji79),
            .c8qmnfk1vqai (c8qmnfk1vqai),
            .pbov8g9yizcwr (pbov8g9yizcwr),
            .t8qjehupeajtzjr (t8qjehupeajtzjr),
            .hhp1rh0x0jn (hhp1rh0x0jn),
            .w9yptl69xj6p (w9yptl69xj6p),
            .yvcpy_gyehs4lji (yvcpy_gyehs4lji), 

            .kted7ph0krq (kted7ph0krq),
            .a93i3d2hji (a93i3d2hji),
            .of5p5cb8p4 (of5p5cb8p4),
            .g1bi1xzuv64 (g1bi1xzuv64),
            .gj6p5b5ik3r9p (gj6p5b5ik3r9p),
            .m1fmaas4oww6 (m1fmaas4oww6),

            .su81e8dxdzng9d (su81e8dxdzng9d),

            .gf33atgy (gf33atgy),
            .ru_wi (ru_wi)
  );


  ux607_gnrl_icb2axi_b # (
            .AW (nm_fj),
            .DW (onr7l),
            .MW (h1b),
            .ALLOW_BURST(o7hawonznex2),
            .ID_W (cibz)
) ar26orka1ajeggs8o0dz9(
            .icb_wrsp_valid (sg96uazxf6dpizg7vad),
            .icb_wrsp_ready (qe9rerwzfqnxm49kvj69u),
            .icb_wrsp_err (ba1jgqojkjt_p5wrx1x),
            .icb_wrsp_excl_ok (jgvpcfglnc5lptyi2ca5hkmuv),
            .icb_wrsp_last (edjq61okne5m2wnwpj4in9),

            .axi_bready (nneek3ep5xykwl),
            .axi_bvalid (g8khua4l0y77zjp),
            .axi_bid (wmlp1a2b),
            .axi_bresp (weop50xb_avne),

            .axi_bus_clk_en (su81e8dxdzng9d),

            .wrsp_burst (slggcmvgdj),
            .wrsp_excl  (homm_w8zq),

            .clk (gf33atgy),
            .rst_n (ru_wi)
  );

endmodule




























module ux607_gnrl_icb_arbt # (
  parameter AW = 32,
  parameter DW = 64,
  parameter USR_W = 1,
  parameter ARBT_SCHEME = 3,


  parameter FIFO_OUTS_NUM = 1,
  parameter FIFO_CUT_READY = 0,

  parameter ARBT_NUM = 4,
  parameter ALLOW_0CYCL_RSP = 1,
  parameter ALLOW_BURST = 0,
  parameter ARBT_PTR_W = 2
) (
  output             arbt_active, 

  output             o_icb_cmd_valid, 
  input              o_icb_cmd_ready, 
  output             o_icb_cmd_read, 
  output [AW-1:0]    o_icb_cmd_addr, 
  output [DW-1:0]    o_icb_cmd_wdata, 
  output [(DW/8-1):0]  o_icb_cmd_wmask,
  output [3-1:0]     o_icb_cmd_burst, 
  output [2-1:0]     o_icb_cmd_beat, 
  output             o_icb_cmd_lock,
  output             o_icb_cmd_excl,
  output [1:0]       o_icb_cmd_size,
  output [USR_W-1:0] o_icb_cmd_usr,

  input              o_icb_rsp_valid, 
  output             o_icb_rsp_ready, 
  input              o_icb_rsp_err,
  input              o_icb_rsp_excl_ok,
  input  [DW-1:0]    o_icb_rsp_rdata, 
  input  [USR_W-1:0] o_icb_rsp_usr, 

  input  [ARBT_NUM*1-1:0]     i_bus_icb_cmd_sel_vec, 

  output [ARBT_NUM*1-1:0]     i_bus_icb_cmd_ready, 
  input  [ARBT_NUM*1-1:0]     i_bus_icb_cmd_valid, 
  input  [ARBT_NUM*1-1:0]     i_bus_icb_cmd_read, 
  input  [ARBT_NUM*AW-1:0]    i_bus_icb_cmd_addr, 
  input  [ARBT_NUM*DW-1:0]    i_bus_icb_cmd_wdata, 
  input  [(ARBT_NUM*DW/8-1):0]  i_bus_icb_cmd_wmask,
  input  [ARBT_NUM*3-1:0]     i_bus_icb_cmd_burst,
  input  [ARBT_NUM*2-1:0]     i_bus_icb_cmd_beat ,
  input  [ARBT_NUM*1-1:0]     i_bus_icb_cmd_lock ,
  input  [ARBT_NUM*1-1:0]     i_bus_icb_cmd_excl ,
  input  [ARBT_NUM*2-1:0]     i_bus_icb_cmd_size ,
  input  [ARBT_NUM*USR_W-1:0] i_bus_icb_cmd_usr  ,

  output [ARBT_NUM*1-1:0]     i_bus_icb_rsp_valid, 
  input  [ARBT_NUM*1-1:0]     i_bus_icb_rsp_ready, 
  output [ARBT_NUM*1-1:0]     i_bus_icb_rsp_err,
  output [ARBT_NUM*1-1:0]     i_bus_icb_rsp_excl_ok,
  output [ARBT_NUM*DW-1:0]    i_bus_icb_rsp_rdata, 
  output [ARBT_NUM*USR_W-1:0] i_bus_icb_rsp_usr, 

  input  clk,  
  input  rst_n
  );

  wire             klkflmsyyf5w7ar; 
  wire             wy36iirxspfw56864; 
  wire             lkjqs6kiuyj;
  wire             u245it8jnyhc3eqcy0;
  wire [DW-1:0]    h7f6k_ims_9p3; 
  wire [USR_W-1:0] iwxu78sftoab_xrp; 

  localparam mp26klefy4v2f = (2+DW+USR_W);
  wire [mp26klefy4v2f-1:0] i2pk7kg6dmy2u8yk = {
                                 o_icb_rsp_err,
                                 o_icb_rsp_excl_ok,
                                 o_icb_rsp_rdata, 
                                 o_icb_rsp_usr};

  wire [mp26klefy4v2f-1:0] pq28r_0p1z8tuc;

  assign {
                                 lkjqs6kiuyj,
                                 u245it8jnyhc3eqcy0,
                                 h7f6k_ims_9p3, 
                                 iwxu78sftoab_xrp} = pq28r_0p1z8tuc;


      assign pq28r_0p1z8tuc = i2pk7kg6dmy2u8yk;
      assign klkflmsyyf5w7ar = o_icb_rsp_valid;
      assign o_icb_rsp_ready = wy36iirxspfw56864;























  wire pjisa4vlo9u0rtnt1whf8;       

  wire [ARBT_NUM-1:0] rhyh7gw3h9wjpo6  ;
  wire [ARBT_NUM-1:0] uq7evk9_yg0c4  ;

genvar i;
generate 
  if(ARBT_NUM == 1) begin:za7a9z3h51xloema0dtt
    assign i_bus_icb_cmd_ready = o_icb_cmd_ready    ;
    assign o_icb_cmd_valid     = i_bus_icb_cmd_valid;
    assign o_icb_cmd_read      = i_bus_icb_cmd_read ;
    assign o_icb_cmd_addr      = i_bus_icb_cmd_addr ;
    assign o_icb_cmd_wdata     = i_bus_icb_cmd_wdata;
    assign o_icb_cmd_wmask     = i_bus_icb_cmd_wmask;
    assign o_icb_cmd_burst     = i_bus_icb_cmd_burst;
    assign o_icb_cmd_beat      = i_bus_icb_cmd_beat ;
    assign o_icb_cmd_lock      = i_bus_icb_cmd_lock ;
    assign o_icb_cmd_excl      = i_bus_icb_cmd_excl ;
    assign o_icb_cmd_size      = i_bus_icb_cmd_size ;
    assign o_icb_cmd_usr       = i_bus_icb_cmd_usr  ;

    assign wy36iirxspfw56864     = i_bus_icb_rsp_ready;
    assign i_bus_icb_rsp_valid = klkflmsyyf5w7ar    ;
    assign i_bus_icb_rsp_err   = lkjqs6kiuyj      ;
    assign i_bus_icb_rsp_excl_ok   = u245it8jnyhc3eqcy0      ;
    assign i_bus_icb_rsp_rdata = h7f6k_ims_9p3    ;
    assign i_bus_icb_rsp_usr   = iwxu78sftoab_xrp      ;

    assign pjisa4vlo9u0rtnt1whf8    = 1'b1;       
    assign rhyh7gw3h9wjpo6 = {ARBT_NUM{1'b0}};
    assign uq7evk9_yg0c4 = {ARBT_NUM{1'b0}};


  end
  else begin:phbyjwvv0j85tlg5vbp

    integer j;

    wire [ARBT_NUM-1:0] cdw1279sjt44_h5gwj339; 
    wire [ARBT_NUM-1:0] p_adc2c56l5xmyiu95kx; 
    wire uofey29hpm21uqkvovbgv_z9e; 
    wire v_2seni8d29s8i4ukr8gt7; 

    wire            ogvavqa7ta836s [ARBT_NUM-1:0]; 
    wire [AW-1:0]   aw0a19a967dn7n0x25w [ARBT_NUM-1:0]; 
    wire [DW-1:0]   sc169gxpr38lpe8[ARBT_NUM-1:0]; 
    wire [(DW/8-1):0] hg1g2yh6yktfe_btdst7[ARBT_NUM-1:0];
    wire [3-1:0]    j4d0rl87t28yrb94i[ARBT_NUM-1:0];
    wire [2-1:0]    k994rox28a17feu [ARBT_NUM-1:0];
    wire            h6hn_gz20krea1 [ARBT_NUM-1:0];
    wire            l089k6vccrfphrtw [ARBT_NUM-1:0];
    wire [2-1:0]    leieaos4fnc5s_81kr [ARBT_NUM-1:0];
    wire [USR_W-1:0]qku53_e41ce0r6rtb  [ARBT_NUM-1:0];

    reg            tu8l_ltlfps3u9e_fv; 
    reg [AW-1:0]   iq9sbyfkr_z42610cta72; 
    reg [DW-1:0]   c7lfsuhab9c8cc73eu3wlt; 
    reg [(DW/8-1):0] mc0m0fq5t3t_0r85d3tu3v2;
    reg [3-1:0]    dxi8twzovrwsqcashzc;
    reg [2-1:0]    xu7o989_k6nc4_yscybd3 ;
    reg            or5ecyb2qdd1ock96q ;
    reg            xhwk2yv2cbngrg9jv6_8pf ;
    reg [2-1:0]    r82v2cg5erf3p2krcdkob ;
    reg [USR_W-1:0]pzjm78nzkhijsjsw6ke  ;

    wire o18xphirvb6rzzl33v; 
    wire qju93nlsmz4hbbz1py5;

    wire djmbzt1843lpcet2xr1d1b;
    wire gp0lafw7tngumfeqku5;
    wire m3ho2mulswsyi6r_r;


    wire jxqrb_9po4b1mxj0al90g;
    wire kbtixer0amhrz2dzvhe;
    wire wr80zcrpu3t413geuk;
    wire nhqlx69jse016ld9w87kjm7;
    wire [ARBT_PTR_W-1:0] ibsurazp9nyl3c3a;
    wire [ARBT_PTR_W-1:0] uogk6x1xf6j9v5w;

    wire ns807okp2nn628yu3u;       
    reg [ARBT_PTR_W-1:0] pczv8skzdtc77h4q;

    wire [ARBT_NUM*1-1:0] qpjg40ms0yzkuyocirhhna8; 
    wire [ARBT_NUM*1-1:0] cgxxwbtde0xaow76pjmil3d; 
    wire [ARBT_NUM*1-1:0] xz28dmfytkmyl1xh36qwa8y8awx97; 

    wire j701sr4kuq;

    wire [ARBT_PTR_W-1:0] t9x9lzcn9i6ak8ykzjqj;

    wire [ARBT_NUM-1:0] hmtgswn3qp6guri3ot;
    wire [ARBT_NUM-1:0] ir5hj_acy6t62jhapc;
    wire [ARBT_NUM-1:0] v21p5eaumf7vz6mz9nb;
    wire [ARBT_NUM-1:0] zduo__k11ouiyz7kj4v;

    if(ALLOW_BURST == 0) begin: ehhzd0qjs0u75yfk5gxqj
      assign uq7evk9_yg0c4   = {ARBT_NUM{1'b0}};
      assign hmtgswn3qp6guri3ot = {ARBT_NUM{1'b0}};
      assign ir5hj_acy6t62jhapc = {ARBT_NUM{1'b0}};
      assign v21p5eaumf7vz6mz9nb = {ARBT_NUM{1'b0}};
      assign zduo__k11ouiyz7kj4v = {ARBT_NUM{1'b0}};

    end

    assign cgxxwbtde0xaow76pjmil3d   = (~uq7evk9_yg0c4) & (~rhyh7gw3h9wjpo6) & i_bus_icb_cmd_valid; 
    assign i_bus_icb_cmd_ready       = (~uq7evk9_yg0c4) & (~rhyh7gw3h9wjpo6) & qpjg40ms0yzkuyocirhhna8; 
    assign xz28dmfytkmyl1xh36qwa8y8awx97 = (~uq7evk9_yg0c4) & (~rhyh7gw3h9wjpo6) & i_bus_icb_cmd_sel_vec; 

    assign o_icb_cmd_valid = uofey29hpm21uqkvovbgv_z9e & (~ns807okp2nn628yu3u);
    assign v_2seni8d29s8i4ukr8gt7 = o_icb_cmd_ready & (~ns807okp2nn628yu3u); 


    for(i = 0; i < ARBT_NUM; i = i+1)
    begin:s9dy2pie07n9wcw_a
      assign ogvavqa7ta836s [i] = i_bus_icb_cmd_read [(i+1)*1     -1 : i*1     ];
      assign aw0a19a967dn7n0x25w [i] = i_bus_icb_cmd_addr [(i+1)*AW    -1 : i*AW    ];
      assign sc169gxpr38lpe8[i] = i_bus_icb_cmd_wdata[(i+1)*DW    -1 : i*DW    ];
      assign hg1g2yh6yktfe_btdst7[i] = i_bus_icb_cmd_wmask[(i+1)*(DW/8)-1 : i*(DW/8)];
      assign j4d0rl87t28yrb94i[i] = i_bus_icb_cmd_burst[(i+1)*3     -1 : i*3     ];
      assign k994rox28a17feu [i] = i_bus_icb_cmd_beat [(i+1)*2     -1 : i*2     ];
      assign h6hn_gz20krea1 [i] = i_bus_icb_cmd_lock [(i+1)*1     -1 : i*1     ];
      assign l089k6vccrfphrtw [i] = i_bus_icb_cmd_excl [(i+1)*1     -1 : i*1     ];
      assign leieaos4fnc5s_81kr [i] = i_bus_icb_cmd_size [(i+1)*2     -1 : i*2     ];
      assign qku53_e41ce0r6rtb  [i] = i_bus_icb_cmd_usr  [(i+1)*USR_W -1 : i*USR_W ];

      assign qpjg40ms0yzkuyocirhhna8[i] = cdw1279sjt44_h5gwj339[i] & v_2seni8d29s8i4ukr8gt7;
      assign i_bus_icb_rsp_valid[i] = qju93nlsmz4hbbz1py5 & (t9x9lzcn9i6ak8ykzjqj == i[ARBT_PTR_W-1:0]); 
    end

    assign j701sr4kuq = o_icb_cmd_valid & o_icb_cmd_ready; 

      wire [ARBT_NUM-1:0] ukf9ivzomgw2zcelt;
      wire [ARBT_NUM-1:0] c5cxxwjakgolj2vze;
      wire [ARBT_NUM-1:0] z2me5m7f6tuw4om;
      wire [ARBT_NUM-1:0] ny9mi_hrx7ij0abt;

      for(i = 0; i < ARBT_NUM; i = i+1) begin:b1jl0upfsk5s1eqmpd


        assign ukf9ivzomgw2zcelt[i] = (p_adc2c56l5xmyiu95kx[i] == 1'b0) & o_icb_cmd_lock & j701sr4kuq;

        assign c5cxxwjakgolj2vze[i] = rhyh7gw3h9wjpo6[i] & ((~o_icb_cmd_lock) & j701sr4kuq);
        assign z2me5m7f6tuw4om[i] = ukf9ivzomgw2zcelt[i] |   c5cxxwjakgolj2vze[i];
        assign ny9mi_hrx7ij0abt[i] = ukf9ivzomgw2zcelt[i] & (~c5cxxwjakgolj2vze[i]);

        ux607_gnrl_dfflr #(1) msyixhqcrbqhloy3t (z2me5m7f6tuw4om[i], ny9mi_hrx7ij0abt[i], rhyh7gw3h9wjpo6[i], clk, rst_n);

      end

    if(ALLOW_BURST == 1) begin: i6oayc_fe7m_j
      for(i = 0; i < ARBT_NUM; i = i+1)
      begin:rj4jt0i34jw1gr_ypv



        assign hmtgswn3qp6guri3ot[i] = (p_adc2c56l5xmyiu95kx[i] == 1'b0) & o_icb_cmd_beat[0] & j701sr4kuq;

        assign ir5hj_acy6t62jhapc[i] = uq7evk9_yg0c4[i] & o_icb_cmd_beat[1] & j701sr4kuq;
        assign v21p5eaumf7vz6mz9nb[i] = hmtgswn3qp6guri3ot[i] |   ir5hj_acy6t62jhapc[i];
        assign zduo__k11ouiyz7kj4v[i] = hmtgswn3qp6guri3ot[i] & (~ir5hj_acy6t62jhapc[i]);

        ux607_gnrl_dfflr #(1) p3n1o95nu5xqfa212ma8y (v21p5eaumf7vz6mz9nb[i], zduo__k11ouiyz7kj4v[i], uq7evk9_yg0c4[i], clk, rst_n);

      end
    end

    if(ARBT_SCHEME == 0) begin:f3869788c0h2pov2un

      for(i = 0; i < ARBT_NUM; i = i+1)
      begin:shr0zu2xtqr9_iq9psn

        if(i==0) begin: xvpcp9wjmb99kn
          assign cdw1279sjt44_h5gwj339[i] =  1'b1;
          assign p_adc2c56l5xmyiu95kx[i] = cdw1279sjt44_h5gwj339[i] & cgxxwbtde0xaow76pjmil3d[i];
        end
        else begin:efbb_rw4_pjzu4jx64w
          assign cdw1279sjt44_h5gwj339[i] =  ~(|cgxxwbtde0xaow76pjmil3d[i-1:0]);
          assign p_adc2c56l5xmyiu95kx[i] = cdw1279sjt44_h5gwj339[i] & cgxxwbtde0xaow76pjmil3d[i];
        end

      end

      assign uofey29hpm21uqkvovbgv_z9e = |cgxxwbtde0xaow76pjmil3d; 

    end

   if(ARBT_SCHEME == 1) begin:grac_7xmxn_m1uvhz0l


     ux607_gnrl_rrobin # (
         .ARBT_NUM(ARBT_NUM)
     )jag2p96lla6f8m7d2t(
       .grt_vec  (cdw1279sjt44_h5gwj339),  
       .req_vec  (cgxxwbtde0xaow76pjmil3d),  
       .arbt_ena (j701sr4kuq),   
       .clk      (clk),
       .rst_n    (rst_n)
     );
     assign p_adc2c56l5xmyiu95kx = cdw1279sjt44_h5gwj339;
     assign uofey29hpm21uqkvovbgv_z9e = |cgxxwbtde0xaow76pjmil3d; 

   end

   if(ARBT_SCHEME == 2) begin:h6fhjx3o8hh6ea

     assign cdw1279sjt44_h5gwj339 = xz28dmfytkmyl1xh36qwa8y8awx97;
     assign p_adc2c56l5xmyiu95kx = cdw1279sjt44_h5gwj339;

     assign uofey29hpm21uqkvovbgv_z9e = |(cgxxwbtde0xaow76pjmil3d & xz28dmfytkmyl1xh36qwa8y8awx97); 
   end

   if(ARBT_SCHEME == 3) begin:rd4ugvmmjocd1j7ozmahqckjf

      for(i = 0; i < ARBT_NUM; i = i+1)
      begin:shr0zu2xtqr9_iq9psn

        if(i==0) begin: xvpcp9wjmb99kn
          assign cdw1279sjt44_h5gwj339[i] =  1'b1;
          assign p_adc2c56l5xmyiu95kx[i] = cdw1279sjt44_h5gwj339[i] & xz28dmfytkmyl1xh36qwa8y8awx97[i];
        end
        else if(i==(ARBT_NUM-1)) begin: ufc5qp4_5o2
          assign cdw1279sjt44_h5gwj339[i] =  ~(|xz28dmfytkmyl1xh36qwa8y8awx97[i-1:0]);
          assign p_adc2c56l5xmyiu95kx[i] = cdw1279sjt44_h5gwj339[i];
        end
        else begin:efbb_rw4_pjzu4jx64w
          assign cdw1279sjt44_h5gwj339[i] =  ~(|xz28dmfytkmyl1xh36qwa8y8awx97[i-1:0]);
          assign p_adc2c56l5xmyiu95kx[i] = cdw1279sjt44_h5gwj339[i] & xz28dmfytkmyl1xh36qwa8y8awx97[i];
        end

      end


      assign uofey29hpm21uqkvovbgv_z9e = |(cgxxwbtde0xaow76pjmil3d & p_adc2c56l5xmyiu95kx); 
    end



   if(ARBT_SCHEME == 4) begin:rp_ug1jk_ggt2pqjp5

      wire ywxj0neeoc3l_4ab = |ukf9ivzomgw2zcelt;


      ux607_gnrl_rbin4 # (
          .ARBT_NUM(ARBT_NUM)
      )io7_7vg_jqrqis89uj(
        .grt_vec  (cdw1279sjt44_h5gwj339),  
        .req_vec  (xz28dmfytkmyl1xh36qwa8y8awx97),  
        .arbt_ena (j701sr4kuq & (~ywxj0neeoc3l_4ab)),   
        .clk      (clk),
        .rst_n    (rst_n)
      );
      assign p_adc2c56l5xmyiu95kx = cdw1279sjt44_h5gwj339 & xz28dmfytkmyl1xh36qwa8y8awx97;

      assign uofey29hpm21uqkvovbgv_z9e = |(cgxxwbtde0xaow76pjmil3d & p_adc2c56l5xmyiu95kx); 
   end


    always @ (*) begin : lh82_td_rnhybm4y5zqrzzru2jbcd
      tu8l_ltlfps3u9e_fv  = {1   {1'b0}};
      iq9sbyfkr_z42610cta72  = {AW  {1'b0}};
      c7lfsuhab9c8cc73eu3wlt = {DW  {1'b0}};
      mc0m0fq5t3t_0r85d3tu3v2 = {DW/8{1'b0}};
      dxi8twzovrwsqcashzc = {3   {1'b0}};
      xu7o989_k6nc4_yscybd3  = {2   {1'b0}};
      or5ecyb2qdd1ock96q  = {1   {1'b0}};
      xhwk2yv2cbngrg9jv6_8pf  = {1   {1'b0}};
      r82v2cg5erf3p2krcdkob  = {2   {1'b0}};
      pzjm78nzkhijsjsw6ke   = {USR_W{1'b0}};
      for(j = 0; j < ARBT_NUM; j = j+1) begin
        tu8l_ltlfps3u9e_fv  = tu8l_ltlfps3u9e_fv  | ({1    {p_adc2c56l5xmyiu95kx[j]}} & ogvavqa7ta836s [j]);
        iq9sbyfkr_z42610cta72  = iq9sbyfkr_z42610cta72  | ({AW   {p_adc2c56l5xmyiu95kx[j]}} & aw0a19a967dn7n0x25w [j]);
        c7lfsuhab9c8cc73eu3wlt = c7lfsuhab9c8cc73eu3wlt | ({DW   {p_adc2c56l5xmyiu95kx[j]}} & sc169gxpr38lpe8[j]);
        mc0m0fq5t3t_0r85d3tu3v2 = mc0m0fq5t3t_0r85d3tu3v2 | ({DW/8 {p_adc2c56l5xmyiu95kx[j]}} & hg1g2yh6yktfe_btdst7[j]);
        dxi8twzovrwsqcashzc = dxi8twzovrwsqcashzc | ({3    {p_adc2c56l5xmyiu95kx[j]}} & j4d0rl87t28yrb94i[j]);
        xu7o989_k6nc4_yscybd3  = xu7o989_k6nc4_yscybd3  | ({2    {p_adc2c56l5xmyiu95kx[j]}} & k994rox28a17feu [j]);
        or5ecyb2qdd1ock96q  = or5ecyb2qdd1ock96q  | ({1    {p_adc2c56l5xmyiu95kx[j]}} & h6hn_gz20krea1 [j]);
        xhwk2yv2cbngrg9jv6_8pf  = xhwk2yv2cbngrg9jv6_8pf  | ({1    {p_adc2c56l5xmyiu95kx[j]}} & l089k6vccrfphrtw [j]);
        r82v2cg5erf3p2krcdkob  = r82v2cg5erf3p2krcdkob  | ({2    {p_adc2c56l5xmyiu95kx[j]}} & leieaos4fnc5s_81kr [j]);
        pzjm78nzkhijsjsw6ke   = pzjm78nzkhijsjsw6ke   | ({USR_W{p_adc2c56l5xmyiu95kx[j]}} & qku53_e41ce0r6rtb  [j]);
      end
    end

    always @ (*) begin : uad8nlh5i4rzz6q361jlqx
      pczv8skzdtc77h4q = {ARBT_PTR_W{1'b0}};
      for(j = 0; j < ARBT_NUM; j = j+1) begin
        pczv8skzdtc77h4q = pczv8skzdtc77h4q | ({ARBT_PTR_W{p_adc2c56l5xmyiu95kx[j]}} & $unsigned(j[ARBT_PTR_W-1:0]));
      end
    end

    assign gp0lafw7tngumfeqku5 = o_icb_cmd_valid & o_icb_cmd_ready;
    assign m3ho2mulswsyi6r_r = klkflmsyyf5w7ar & wy36iirxspfw56864;


    if(ALLOW_0CYCL_RSP == 1) begin: ywf24098_gi8bfyn2w
        assign djmbzt1843lpcet2xr1d1b = pjisa4vlo9u0rtnt1whf8 & gp0lafw7tngumfeqku5 & m3ho2mulswsyi6r_r;
        assign t9x9lzcn9i6ak8ykzjqj = pjisa4vlo9u0rtnt1whf8 ? uogk6x1xf6j9v5w : ibsurazp9nyl3c3a;

        assign qju93nlsmz4hbbz1py5 = klkflmsyyf5w7ar;
        assign wy36iirxspfw56864     = o18xphirvb6rzzl33v;
    end
    else begin: ss_g5sktytsbln200rqk
        assign djmbzt1843lpcet2xr1d1b   = 1'b0;
        assign t9x9lzcn9i6ak8ykzjqj   = ibsurazp9nyl3c3a;
        assign qju93nlsmz4hbbz1py5 = (~pjisa4vlo9u0rtnt1whf8) & klkflmsyyf5w7ar;
        assign wy36iirxspfw56864     = (~pjisa4vlo9u0rtnt1whf8) & o18xphirvb6rzzl33v;
    end

    assign jxqrb_9po4b1mxj0al90g = gp0lafw7tngumfeqku5 & (~djmbzt1843lpcet2xr1d1b);
    assign ns807okp2nn628yu3u    = (~wr80zcrpu3t413geuk);
    assign nhqlx69jse016ld9w87kjm7 = m3ho2mulswsyi6r_r & (~djmbzt1843lpcet2xr1d1b);
    assign pjisa4vlo9u0rtnt1whf8   = (~kbtixer0amhrz2dzvhe);

    assign uogk6x1xf6j9v5w   = pczv8skzdtc77h4q;

    if(FIFO_OUTS_NUM == 1) begin:cxgfpc10
      ux607_gnrl_pipe_stage # (
        .CUT_READY (FIFO_CUT_READY),
        .DP  (1),
        .DW  (ARBT_PTR_W)
      ) ahkryar1lc8lsjv5v1c_6ce6 (
        .i_vld(jxqrb_9po4b1mxj0al90g),
        .i_rdy(wr80zcrpu3t413geuk),
        .i_dat(uogk6x1xf6j9v5w ),
        .o_vld(kbtixer0amhrz2dzvhe),
        .o_rdy(nhqlx69jse016ld9w87kjm7),  
        .o_dat(ibsurazp9nyl3c3a ),  
        .clk  (clk),
        .rst_n(rst_n)
      );

    end
    else begin: rujquo369cvzmr5
      ux607_gnrl_fifo # (
        .CUT_READY (FIFO_CUT_READY),
        .MSKO      (0),
        .DP  (FIFO_OUTS_NUM),
        .DW  (ARBT_PTR_W)
      ) ahkryar1lc8lsjv5v1c_6ce6 (
        .i_vld(jxqrb_9po4b1mxj0al90g),
        .i_rdy(wr80zcrpu3t413geuk),
        .i_dat(uogk6x1xf6j9v5w ),
        .o_vld(kbtixer0amhrz2dzvhe),
        .o_rdy(nhqlx69jse016ld9w87kjm7),  
        .o_dat(ibsurazp9nyl3c3a ),  

        .clk  (clk),
        .rst_n(rst_n)
      );
    end

    assign o_icb_cmd_read  = tu8l_ltlfps3u9e_fv ; 
    assign o_icb_cmd_addr  = iq9sbyfkr_z42610cta72 ; 
    assign o_icb_cmd_wdata = c7lfsuhab9c8cc73eu3wlt; 
    assign o_icb_cmd_wmask = mc0m0fq5t3t_0r85d3tu3v2;
    assign o_icb_cmd_burst = dxi8twzovrwsqcashzc;
    assign o_icb_cmd_beat  = xu7o989_k6nc4_yscybd3 ;
    assign o_icb_cmd_lock  = or5ecyb2qdd1ock96q ;
    assign o_icb_cmd_excl  = xhwk2yv2cbngrg9jv6_8pf ;
    assign o_icb_cmd_size  = r82v2cg5erf3p2krcdkob ;
    assign o_icb_cmd_usr   = pzjm78nzkhijsjsw6ke  ;

    assign o18xphirvb6rzzl33v = i_bus_icb_rsp_ready[t9x9lzcn9i6ak8ykzjqj]; 



    assign i_bus_icb_rsp_err     = {ARBT_NUM{lkjqs6kiuyj  }};  
    assign i_bus_icb_rsp_excl_ok = {ARBT_NUM{u245it8jnyhc3eqcy0}};  
    assign i_bus_icb_rsp_rdata   = {ARBT_NUM{h7f6k_ims_9p3}}; 
    assign i_bus_icb_rsp_usr     = {ARBT_NUM{iwxu78sftoab_xrp}}; 
  end
  endgenerate 

  assign arbt_active = (|i_bus_icb_cmd_valid) | (~pjisa4vlo9u0rtnt1whf8) | klkflmsyyf5w7ar  
                     | (|uq7evk9_yg0c4) | (|rhyh7gw3h9wjpo6);

endmodule








module ux607_gnrl_icb_buffer # (
  parameter CMD_MSKO = 0,
  parameter OUTS_CNT_W = 1,
  parameter AW = 32,
  parameter DW = 32,
  parameter CMD_CUT_READY = 0,
  parameter RSP_CUT_READY = 0,
  parameter CMD_DP = 0,
  parameter RSP_DP = 0,

  parameter RSP_ALWAYS_READY = 0,
  parameter USR_W = 1
) (
  input              bus_clk_en,

  output             icb_buffer_active,

  input              i_icb_cmd_valid, 
  output             i_icb_cmd_ready, 
  input              i_icb_cmd_read, 
  input  [AW-1:0]    i_icb_cmd_addr, 
  input  [DW-1:0]    i_icb_cmd_wdata, 
  input  [(DW/8-1):0]  i_icb_cmd_wmask,
  input              i_icb_cmd_lock,
  input              i_icb_cmd_excl,
  input  [1:0]       i_icb_cmd_size,
  input  [2:0]       i_icb_cmd_burst,
  input  [1:0]       i_icb_cmd_beat,
  input  [USR_W-1:0] i_icb_cmd_usr,

  output             i_icb_rsp_valid, 
  input              i_icb_rsp_ready, 
  output             i_icb_rsp_err,
  output             i_icb_rsp_excl_ok,
  output [DW-1:0]    i_icb_rsp_rdata, 
  output [USR_W-1:0] i_icb_rsp_usr,

  output             o_icb_cmd_valid, 
  input              o_icb_cmd_ready, 
  output             o_icb_cmd_read, 
  output [AW-1:0]    o_icb_cmd_addr, 
  output [DW-1:0]    o_icb_cmd_wdata, 
  output [(DW/8-1):0]  o_icb_cmd_wmask,
  output             o_icb_cmd_lock,
  output             o_icb_cmd_excl,
  output [1:0]       o_icb_cmd_size,
  output [2:0]       o_icb_cmd_burst,
  output [1:0]       o_icb_cmd_beat,
  output [USR_W-1:0] o_icb_cmd_usr,

  input              o_icb_rsp_valid, 
  output             o_icb_rsp_ready, 
  input              o_icb_rsp_err,
  input              o_icb_rsp_excl_ok,
  input  [DW-1:0]    o_icb_rsp_rdata, 
  input  [USR_W-1:0] o_icb_rsp_usr,

  input  clk,  
  input  rst_n
  );

  localparam f16zrowg1s1f5 = (1+AW+DW+(DW/8)+1+1+3+2+2+USR_W);

  wire [f16zrowg1s1f5-1:0] vwuqk746df8rzf = {
                                 i_icb_cmd_read, 
                                 i_icb_cmd_addr, 
                                 i_icb_cmd_wdata, 
                                 i_icb_cmd_wmask,
                                 i_icb_cmd_lock,
                                 i_icb_cmd_excl,
                                 i_icb_cmd_size,
                                 i_icb_cmd_burst,
                                 i_icb_cmd_beat,
                                 i_icb_cmd_usr};

  wire [f16zrowg1s1f5-1:0] f1lo32g6mtt5xv;

  assign {
                                 o_icb_cmd_read, 
                                 o_icb_cmd_addr, 
                                 o_icb_cmd_wdata, 
                                 o_icb_cmd_wmask,
                                 o_icb_cmd_lock,
                                 o_icb_cmd_excl,
                                 o_icb_cmd_size,
                                 o_icb_cmd_burst,
                                 o_icb_cmd_beat,
                                 o_icb_cmd_usr} = f1lo32g6mtt5xv;

  wire g2tqgfxuk3a_ininxip0; 
  wire oesnimkjbwlow8m2tt7jix; 

  wire eawl4k3d3kw4r0ijlw8y9; 
  wire r_ka1cs6ztb7tu2j; 
  assign eawl4k3d3kw4r0ijlw8y9 = bus_clk_en & i_icb_cmd_valid; 
  assign i_icb_cmd_ready  = bus_clk_en & r_ka1cs6ztb7tu2j; 

  ux607_gnrl_fifo # (
    .CUT_READY (CMD_CUT_READY),
    .MSKO      (CMD_MSKO),
    .DP  (CMD_DP),
    .DW  (f16zrowg1s1f5)
  ) sonxop729j1hw_fvx7ar4zi (
    .i_vld(eawl4k3d3kw4r0ijlw8y9),
    .i_rdy(r_ka1cs6ztb7tu2j),
    .i_dat(vwuqk746df8rzf ),
    .o_vld(g2tqgfxuk3a_ininxip0),
    .o_rdy(oesnimkjbwlow8m2tt7jix),  
    .o_dat(f1lo32g6mtt5xv ),  

    .clk  (clk),
    .rst_n(rst_n)
  );

  wire xivnbyfcz0ixh;

  generate 
    if(RSP_ALWAYS_READY == 1) begin: loll76014dqv_bk0654z9_jk
      assign o_icb_cmd_valid     = xivnbyfcz0ixh & g2tqgfxuk3a_ininxip0; 
      assign oesnimkjbwlow8m2tt7jix = xivnbyfcz0ixh & o_icb_cmd_ready; 
    end
    else begin: llgd5y_nnmt70jc425enmt
      assign o_icb_cmd_valid     = g2tqgfxuk3a_ininxip0; 
      assign oesnimkjbwlow8m2tt7jix = o_icb_cmd_ready; 
    end
  endgenerate



  localparam mp26klefy4v2f = (2+DW+USR_W);
  wire [mp26klefy4v2f-1:0] i2pk7kg6dmy2u8yk = {
                                 o_icb_rsp_err,
                                 o_icb_rsp_excl_ok,
                                 o_icb_rsp_rdata, 
                                 o_icb_rsp_usr};

  wire [mp26klefy4v2f-1:0] pq28r_0p1z8tuc;

  assign {
                                 i_icb_rsp_err,
                                 i_icb_rsp_excl_ok,
                                 i_icb_rsp_rdata, 
                                 i_icb_rsp_usr} = pq28r_0p1z8tuc;



      ux607_gnrl_fifo # (
        .CUT_READY (RSP_CUT_READY),
        .MSKO      (0),
        .DP  (RSP_DP),
        .DW  (mp26klefy4v2f)
      ) csn98uaoatfnyzyk5x_ksl_ (
        .i_vld(o_icb_rsp_valid),
        .i_rdy(o_icb_rsp_ready),
        .i_dat(i2pk7kg6dmy2u8yk ),
        .o_vld(i_icb_rsp_valid),
        .o_rdy(i_icb_rsp_ready),  
        .o_dat(pq28r_0p1z8tuc ),  

        .clk  (clk),
        .rst_n(rst_n)
      );



























  wire kouhyfs99s2xt8qfr = i_icb_cmd_valid & i_icb_cmd_ready & bus_clk_en;
  wire yk4t8yu2epj8 = i_icb_rsp_valid & i_icb_rsp_ready & bus_clk_en;

  wire r8axmur45uwwts_z = kouhyfs99s2xt8qfr ^ yk4t8yu2epj8;

  wire [OUTS_CNT_W-1:0] ta6v7ss882s4;
  wire [OUTS_CNT_W-1:0] w71i8osb89s79fy = kouhyfs99s2xt8qfr ? (ta6v7ss882s4 + 1'b1) : (ta6v7ss882s4 - 1'b1);
  ux607_gnrl_dfflr #(OUTS_CNT_W) hh67nplqgwfr382l5y7 (r8axmur45uwwts_z, w71i8osb89s79fy, ta6v7ss882s4, clk, rst_n);

  assign icb_buffer_active = 

      i_icb_cmd_valid | (~(ta6v7ss882s4 == {OUTS_CNT_W{1'b0}}));

  wire ac9xzowkbfofvivbgld = o_icb_cmd_valid & o_icb_cmd_ready & bus_clk_en;
  wire d52ga4eujifacqz3fm = i_icb_rsp_valid & i_icb_rsp_ready & bus_clk_en;

  wire gxnrnqvawiublwaex = ac9xzowkbfofvivbgld ^ d52ga4eujifacqz3fm;

  wire [OUTS_CNT_W-1:0] xocrolyqnx55w9_l;
  wire [OUTS_CNT_W-1:0] rap64cg93y4vrhfxj = ac9xzowkbfofvivbgld ? (xocrolyqnx55w9_l + 1'b1) : (xocrolyqnx55w9_l - 1'b1);
  ux607_gnrl_dfflr #(OUTS_CNT_W) dzj2_y_jf3ro_xh1g489 (gxnrnqvawiublwaex, rap64cg93y4vrhfxj, xocrolyqnx55w9_l, clk, rst_n);

  wire [OUTS_CNT_W-1:0] wdg0cf05gpk_lf = gxnrnqvawiublwaex ? rap64cg93y4vrhfxj : xocrolyqnx55w9_l;

  assign xivnbyfcz0ixh = ~(xocrolyqnx55w9_l   == RSP_DP[OUTS_CNT_W-1:0]);


endmodule








module gg8y0ynhq316osuxxk11w2j04po # (
  parameter hejad2_b4dywimoxw5 = 0,
  parameter evi4vkasjp742kf4 = 0, 
  parameter b_qpb_ch = 0,
  parameter ys68i6_dw7b2m2 = 1,
  parameter nm_fj = 32,
  parameter onr7l = 32,
  parameter q8s6zigflsp6aqc4dx = 0,
  parameter m4i6t98hqvrs_enkod = 0,
  parameter xrvos0msri0 = 2,
  parameter b8vod12 = 2,

  parameter w1ztl72rp0snpfsmgyhg = 0,
  parameter s3xvyho = 1
) (
  input              aqamddt_moiuy,
  input              rlwva_uzdseg,

  output             zmzpuim70lsljt2ccu2c1,

  input              v9ov1b3vn5k4ctkb, 
  output             ub9pjiu4juf6nuqoq2w6, 
  input              ogvavqa7ta836s, 
  input  [nm_fj-1:0]    aw0a19a967dn7n0x25w, 
  input  [onr7l-1:0]    sc169gxpr38lpe8, 
  input  [(onr7l/8-1):0]  hg1g2yh6yktfe_btdst7,
  input              h6hn_gz20krea1,
  input              l089k6vccrfphrtw,
  input  [1:0]       leieaos4fnc5s_81kr,
  input  [2:0]       j4d0rl87t28yrb94i,
  input  [1:0]       k994rox28a17feu,
  input  [s3xvyho-1:0] qku53_e41ce0r6rtb,

  output             dy9ll1o6t6ytby71hf4, 
  input              ow4hbh48f0mt6le4o, 
  output             uzwj715coelxmfqs,
  output             sihcnyg6z96riwnnw_np,
  output [onr7l-1:0]    dek0xt7q6guk2vf6, 
  output [s3xvyho-1:0] efi4ga746crcrx,

  output             me2s8h5yw65ail5, 
  input              dtyl4o87hqhm03wj57, 
  output             xiyx61_yd314uojrls, 
  output [nm_fj-1:0]    k68zoq6vpu0olvs99f, 
  output [onr7l-1:0]    m63rlc2ixlaphiq, 
  output [(onr7l/8-1):0]  drdtbfa60cpn5ihc,
  output             da5mm7z1qer9hx385ck,
  output             tg7q7ezs0lgu3bv36l4,
  output [1:0]       hycxa49k327vm1ncjh,
  output [2:0]       rnrkzgtukyiil52jqbp7,
  output [1:0]       wta_51f6oa6zy5t,
  output [s3xvyho-1:0] vzw7nivk4j2idd,

  input              mg6xxata423v5aaikz4v, 
  output             yuew3x5jdkrr87g, 
  input              nkx3bwv604xt1,
  input              db9kwedxc8ekbwcenl8s9,
  input  [onr7l-1:0]    lbvrc0jeu6t70bw, 
  input  [s3xvyho-1:0] wxjl9xtjejiyjn1,

  input  gf33atgy,  
  input  ru_wi
  );

  localparam f16zrowg1s1f5 = (1+nm_fj+onr7l+(onr7l/8)+1+1+3+2+2+s3xvyho);

  wire [f16zrowg1s1f5-1:0] vwuqk746df8rzf = {
                                 ogvavqa7ta836s, 
                                 aw0a19a967dn7n0x25w, 
                                 sc169gxpr38lpe8, 
                                 hg1g2yh6yktfe_btdst7,
                                 h6hn_gz20krea1,
                                 l089k6vccrfphrtw,
                                 leieaos4fnc5s_81kr,
                                 j4d0rl87t28yrb94i,
                                 k994rox28a17feu,
                                 qku53_e41ce0r6rtb};

  wire [f16zrowg1s1f5-1:0] f1lo32g6mtt5xv;

  assign {
                                 xiyx61_yd314uojrls, 
                                 k68zoq6vpu0olvs99f, 
                                 m63rlc2ixlaphiq, 
                                 drdtbfa60cpn5ihc,
                                 da5mm7z1qer9hx385ck,
                                 tg7q7ezs0lgu3bv36l4,
                                 hycxa49k327vm1ncjh,
                                 rnrkzgtukyiil52jqbp7,
                                 wta_51f6oa6zy5t,
                                 vzw7nivk4j2idd} = f1lo32g6mtt5xv;

  wire g2tqgfxuk3a_ininxip0; 
  wire oesnimkjbwlow8m2tt7jix; 

  wire eawl4k3d3kw4r0ijlw8y9; 
  wire r_ka1cs6ztb7tu2j; 
  assign eawl4k3d3kw4r0ijlw8y9 = v9ov1b3vn5k4ctkb; 
  assign ub9pjiu4juf6nuqoq2w6  = r_ka1cs6ztb7tu2j; 

  wire ouxa7qfp_oicc4wo30tx3;

  vq28fpkbg0dxljs8bf0k # (
    .hejad2_b4dywimoxw5 (hejad2_b4dywimoxw5),
    .evi4vkasjp742kf4 (evi4vkasjp742kf4),
    .mhdlk  (xrvos0msri0),
    .onr7l  (f16zrowg1s1f5)
  ) apgmwplppfmc5zlbz8pb2 (
    .i0lklnhw28rc7dj(ouxa7qfp_oicc4wo30tx3),
    .geml8twgru(aqamddt_moiuy),
    .bw6ftrau0(eawl4k3d3kw4r0ijlw8y9),
    .eef2g8(r_ka1cs6ztb7tu2j),
    .qbjvs30wtb(vwuqk746df8rzf ),
    .td5hjljc_(rlwva_uzdseg),
    .wqljp(g2tqgfxuk3a_ininxip0),
    .h9378(oesnimkjbwlow8m2tt7jix),  
    .dqgck5s(f1lo32g6mtt5xv ),  

    .gf33atgy  (gf33atgy),
    .ru_wi(ru_wi)
  );

  wire xivnbyfcz0ixh;

  generate 
    if(w1ztl72rp0snpfsmgyhg == 1) begin: loll76014dqv_bk0654z9_jk
      assign me2s8h5yw65ail5     = xivnbyfcz0ixh & g2tqgfxuk3a_ininxip0; 
      assign oesnimkjbwlow8m2tt7jix = xivnbyfcz0ixh & dtyl4o87hqhm03wj57; 
    end
    else begin: llgd5y_nnmt70jc425enmt
      assign me2s8h5yw65ail5     = g2tqgfxuk3a_ininxip0; 
      assign oesnimkjbwlow8m2tt7jix = dtyl4o87hqhm03wj57; 
    end
  endgenerate



  localparam mp26klefy4v2f = (2+onr7l+s3xvyho);
  wire [mp26klefy4v2f-1:0] i2pk7kg6dmy2u8yk = {
                                 nkx3bwv604xt1,
                                 db9kwedxc8ekbwcenl8s9,
                                 lbvrc0jeu6t70bw, 
                                 wxjl9xtjejiyjn1};

  wire [mp26klefy4v2f-1:0] pq28r_0p1z8tuc;

  assign {
                                 uzwj715coelxmfqs,
                                 sihcnyg6z96riwnnw_np,
                                 dek0xt7q6guk2vf6, 
                                 efi4ga746crcrx} = pq28r_0p1z8tuc;



      vq28fpkbg0dxljs8bf0k # (
        .hejad2_b4dywimoxw5 (evi4vkasjp742kf4),
        .evi4vkasjp742kf4 (hejad2_b4dywimoxw5),
        .mhdlk  (b8vod12),
        .onr7l  (mp26klefy4v2f)
      ) csn98uaoatfnyzyk5x_ksl_ (
        .geml8twgru(rlwva_uzdseg),
        .bw6ftrau0(mg6xxata423v5aaikz4v),
        .eef2g8(yuew3x5jdkrr87g),
        .qbjvs30wtb(i2pk7kg6dmy2u8yk ),
        .td5hjljc_(aqamddt_moiuy),
        .wqljp(dy9ll1o6t6ytby71hf4),
        .h9378(ow4hbh48f0mt6le4o),  
        .dqgck5s(pq28r_0p1z8tuc ),  

        .i0lklnhw28rc7dj(),
        .gf33atgy  (gf33atgy),
        .ru_wi(ru_wi)
      );

































  wire kouhyfs99s2xt8qfr = v9ov1b3vn5k4ctkb & ub9pjiu4juf6nuqoq2w6 & aqamddt_moiuy;
  wire yk4t8yu2epj8 = dy9ll1o6t6ytby71hf4 & ow4hbh48f0mt6le4o & aqamddt_moiuy;

  wire r8axmur45uwwts_z = kouhyfs99s2xt8qfr ^ yk4t8yu2epj8;

  wire [ys68i6_dw7b2m2-1:0] ta6v7ss882s4;
  wire [ys68i6_dw7b2m2-1:0] w71i8osb89s79fy = kouhyfs99s2xt8qfr ? (ta6v7ss882s4 + 1'b1) : (ta6v7ss882s4 - 1'b1);
  ux607_gnrl_dfflr #(ys68i6_dw7b2m2) hh67nplqgwfr382l5y7 (r8axmur45uwwts_z, w71i8osb89s79fy, ta6v7ss882s4, gf33atgy, ru_wi);

  assign zmzpuim70lsljt2ccu2c1 = 

      v9ov1b3vn5k4ctkb | ouxa7qfp_oicc4wo30tx3 | (~(ta6v7ss882s4 == {ys68i6_dw7b2m2{1'b0}}));

  wire ac9xzowkbfofvivbgld = me2s8h5yw65ail5 & dtyl4o87hqhm03wj57 & rlwva_uzdseg;
  wire d52ga4eujifacqz3fm = dy9ll1o6t6ytby71hf4 & ow4hbh48f0mt6le4o & aqamddt_moiuy;

  wire gxnrnqvawiublwaex = ac9xzowkbfofvivbgld ^ d52ga4eujifacqz3fm;

  wire [ys68i6_dw7b2m2-1:0] xocrolyqnx55w9_l;
  wire [ys68i6_dw7b2m2-1:0] rap64cg93y4vrhfxj = ac9xzowkbfofvivbgld ? (xocrolyqnx55w9_l + 1'b1) : (xocrolyqnx55w9_l - 1'b1);
  ux607_gnrl_dfflr #(ys68i6_dw7b2m2) dzj2_y_jf3ro_xh1g489 (gxnrnqvawiublwaex, rap64cg93y4vrhfxj, xocrolyqnx55w9_l, gf33atgy, ru_wi);

  wire [ys68i6_dw7b2m2-1:0] wdg0cf05gpk_lf = gxnrnqvawiublwaex ? rap64cg93y4vrhfxj : xocrolyqnx55w9_l;

  wire g_t9p4x3pll74onz2sntrv = ~(xocrolyqnx55w9_l   == b8vod12[ys68i6_dw7b2m2-1:0]);
  wire ia6qzifxfp1274kvu3_ = ~(wdg0cf05gpk_lf == b8vod12[ys68i6_dw7b2m2-1:0]);


    wire l2kwhv43umaib = gxnrnqvawiublwaex; 
    wire kun4jk6p0x4b2bao34n;
    wire y9phf0tdehb0aev83ri = (l2kwhv43umaib && !rlwva_uzdseg);
    wire tr_pczcm87014ah6h9 = (kun4jk6p0x4b2bao34n && rlwva_uzdseg);
    wire w5tjv7yt39rnigu_u_l = y9phf0tdehb0aev83ri || tr_pczcm87014ah6h9;
    wire lmanup378q1qzwldb5 = y9phf0tdehb0aev83ri;
    ux607_gnrl_dfflr  #(1) bgspwk95kxsppsiarqazq7sm    (w5tjv7yt39rnigu_u_l, lmanup378q1qzwldb5, kun4jk6p0x4b2bao34n,     gf33atgy, ru_wi);

    wire k0wzgi364_3y212iy5;
    wire cp1fvdzzdqmx4y9v30_ = rlwva_uzdseg && (l2kwhv43umaib || kun4jk6p0x4b2bao34n);
    wire ssfq6skirzz69ut3wyr0 = (l2kwhv43umaib ? ia6qzifxfp1274kvu3_ : g_t9p4x3pll74onz2sntrv);
    ux607_gnrl_dfflrs  #(1) c6wpvkjomo5ivtwng5u2_g9ks    (cp1fvdzzdqmx4y9v30_, ssfq6skirzz69ut3wyr0, k0wzgi364_3y212iy5,     gf33atgy, ru_wi);

  assign xivnbyfcz0ixh = k0wzgi364_3y212iy5;

endmodule







module ux607_gnrl_icb_n2w # (
  parameter AW = 32,
  parameter USR_W = 1,
  parameter FIFO_OUTS_NUM = 8,
  parameter FIFO_CUT_READY = 0,
  parameter X_W = 32,
  parameter Y_W = 64
) (
  input              i_icb_cmd_valid, 
  output             i_icb_cmd_ready, 
  input              i_icb_cmd_read, 
  input  [AW-1:0]    i_icb_cmd_addr, 
  input  [X_W-1:0]   i_icb_cmd_wdata, 
  input  [(X_W/8-1):0] i_icb_cmd_wmask,
  input              i_icb_cmd_lock,
  input              i_icb_cmd_excl,
  input  [1:0]       i_icb_cmd_size,
  input  [2:0]       i_icb_cmd_burst,
  input  [1:0]       i_icb_cmd_beat,
  input  [USR_W-1:0] i_icb_cmd_usr,

  output             i_icb_rsp_valid, 
  input              i_icb_rsp_ready, 
  output             i_icb_rsp_err,
  output             i_icb_rsp_excl_ok,
  output [X_W-1:0]   i_icb_rsp_rdata, 
  output [USR_W-1:0] i_icb_rsp_usr,

  output             o_icb_cmd_valid, 
  input              o_icb_cmd_ready, 
  output             o_icb_cmd_read, 
  output [AW-1:0]    o_icb_cmd_addr, 
  output [Y_W-1:0]   o_icb_cmd_wdata, 
  output [(Y_W/8-1):0] o_icb_cmd_wmask,
  output             o_icb_cmd_lock,
  output             o_icb_cmd_excl,
  output [1:0]       o_icb_cmd_size,
  output [2:0]       o_icb_cmd_burst,
  output [1:0]       o_icb_cmd_beat,
  output [USR_W-1:0] o_icb_cmd_usr,

  input              o_icb_rsp_valid, 
  output             o_icb_rsp_ready, 
  input              o_icb_rsp_err,
  input              o_icb_rsp_excl_ok,
  input  [Y_W-1:0]   o_icb_rsp_rdata, 
  input  [USR_W-1:0] o_icb_rsp_usr,

  input  clk,  
  input  rst_n
  );


    wire de3xfv8sfos;
    wire t7xhkpciv6y402;

    wire hjqolsbb2pa6l = i_icb_cmd_valid & i_icb_cmd_ready;
    wire pt2bqzd5hnjcqv8m = i_icb_rsp_valid & i_icb_rsp_ready;

    wire ujjep82dtrl30kuula;
    wire bf85rp4zf2u_u3lz = hjqolsbb2pa6l;
    wire c6c2z53fscne3    = (~ujjep82dtrl30kuula);
    wire ecz8evddhu0z67ft0w7az ;
    wire fa1tx7irukwu_oa4j5nj = pt2bqzd5hnjcqv8m;
    wire q60zgikcwu82o2   = (~ecz8evddhu0z67ft0w7az);

  generate
    if(FIFO_OUTS_NUM == 1) begin:axug194an99bql_f8e
      ux607_gnrl_pipe_stage # (
        .CUT_READY (FIFO_CUT_READY),
        .DP  (1),
        .DW  (1)
      ) f6qervsn6byr85ihnxbr (
        .i_vld(bf85rp4zf2u_u3lz),
        .i_rdy(ujjep82dtrl30kuula),
        .i_dat(de3xfv8sfos ),
        .o_vld(ecz8evddhu0z67ft0w7az),
        .o_rdy(fa1tx7irukwu_oa4j5nj),  
        .o_dat(t7xhkpciv6y402 ),  

        .clk  (clk),
        .rst_n(rst_n)
      );

    end
    else begin: ayrjh6ok2h5s8a98q
      ux607_gnrl_fifo # (
        .CUT_READY (FIFO_CUT_READY),
        .MSKO      (0),
        .DP  (FIFO_OUTS_NUM),
        .DW  (1)
      ) f6qervsn6byr85ihnxbr (
        .i_vld(bf85rp4zf2u_u3lz),
        .i_rdy(ujjep82dtrl30kuula),
        .i_dat(de3xfv8sfos ),
        .o_vld(ecz8evddhu0z67ft0w7az),
        .o_rdy(fa1tx7irukwu_oa4j5nj),  
        .o_dat(t7xhkpciv6y402 ),  

        .clk  (clk),
        .rst_n(rst_n)
      );
    end
  endgenerate



  generate
    if(X_W == 32) begin: nj8x4m3p1g
      if(Y_W == 64) begin: fqo8yh5gosrncjf
        assign de3xfv8sfos = i_icb_cmd_addr[2]; 
      end
    end
  endgenerate

  assign o_icb_cmd_valid = (~c6c2z53fscne3) & i_icb_cmd_valid; 
  assign i_icb_cmd_ready = (~c6c2z53fscne3) & o_icb_cmd_ready; 
  assign o_icb_cmd_read  = i_icb_cmd_read ;
  assign o_icb_cmd_addr  = i_icb_cmd_addr ;
  assign o_icb_cmd_lock  = i_icb_cmd_lock ;
  assign o_icb_cmd_excl  = i_icb_cmd_excl ;
  assign o_icb_cmd_size  = i_icb_cmd_size ;
  assign o_icb_cmd_burst = i_icb_cmd_burst;
  assign o_icb_cmd_beat  = i_icb_cmd_beat ;
  assign o_icb_cmd_usr   = i_icb_cmd_usr  ;

  assign o_icb_cmd_wdata = {i_icb_cmd_wdata,i_icb_cmd_wdata};
  assign o_icb_cmd_wmask = de3xfv8sfos ?  {i_icb_cmd_wmask,  {X_W/8{1'b0}}} : {  {X_W/8{1'b0}},i_icb_cmd_wmask};

  assign i_icb_rsp_valid = o_icb_rsp_valid ;
  assign i_icb_rsp_err   = o_icb_rsp_err   ;
  assign i_icb_rsp_excl_ok   = o_icb_rsp_excl_ok   ;
  assign i_icb_rsp_rdata = t7xhkpciv6y402 ?  o_icb_rsp_rdata[Y_W-1:X_W] : o_icb_rsp_rdata[X_W-1:0] ;
  assign i_icb_rsp_usr   = o_icb_rsp_usr   ;
  assign o_icb_rsp_ready = i_icb_rsp_ready;  

endmodule







module ux607_gnrl_icb_w2n # (
  parameter LATE_READY = 0,
  parameter ZEROCYC_RSP = 0,
  parameter AW = 64,
  parameter USR_W = 1,
  parameter FIFO_OUTS_NUM = 8,
  parameter FIFO_CUT_READY = 0,
  parameter X_W = 64,
  parameter Y_W = 32 
) (
  input              i_icb_cmd_valid, 
  output             i_icb_cmd_ready, 
  input              i_icb_cmd_read, 
  input  [AW-1:0]    i_icb_cmd_addr, 
  input  [X_W-1:0]   i_icb_cmd_wdata, 
  input  [(X_W/8-1):0] i_icb_cmd_wmask,
  input              i_icb_cmd_lock,
  input              i_icb_cmd_excl,
  input  [1:0]       i_icb_cmd_size,
  input  [2:0]       i_icb_cmd_burst,
  input  [1:0]       i_icb_cmd_beat,
  input  [USR_W-1:0] i_icb_cmd_usr,

  output             i_icb_rsp_valid, 
  input              i_icb_rsp_ready, 
  output             i_icb_rsp_err,
  output             i_icb_rsp_excl_ok,
  output [X_W-1:0]   i_icb_rsp_rdata, 
  output [USR_W-1:0] i_icb_rsp_usr,

  output             o_icb_cmd_valid, 
  input              o_icb_cmd_ready, 
  output             o_icb_cmd_read, 
  output [AW-1:0]    o_icb_cmd_addr, 
  output [Y_W-1:0]   o_icb_cmd_wdata, 
  output [(Y_W/8-1):0] o_icb_cmd_wmask,
  output             o_icb_cmd_lock,
  output             o_icb_cmd_excl,
  output [1:0]       o_icb_cmd_size,
  output [2:0]       o_icb_cmd_burst,
  output [1:0]       o_icb_cmd_beat,
  output [USR_W-1:0] o_icb_cmd_usr,

  input              o_icb_rsp_valid, 
  output             o_icb_rsp_ready, 
  input              o_icb_rsp_err,
  input              o_icb_rsp_excl_ok,
  input  [Y_W-1:0]   o_icb_rsp_rdata, 
  input  [USR_W-1:0] o_icb_rsp_usr,

  input  clk,  
  input  rst_n
  );

  wire skq4j6qdkmbvs1k9lufa = (i_icb_cmd_size[1:0] == 2'b11);
  wire rg2wqryxlxihjmh4v  = i_icb_cmd_addr[2];

  wire j635vgr56_1t4_a8j = i_icb_cmd_valid & i_icb_cmd_ready;
  wire ci10vymorrqh8a = i_icb_rsp_valid & i_icb_rsp_ready;

  wire cyags_6gth1ma8wjx896 = j635vgr56_1t4_a8j;  
  wire y1l45u9lhj0l_z8ry7s_4;
  wire mw8igz4fx7cd12mg;
  wire x43j9vfjtxotxnel20jv = ci10vymorrqh8a;
  wire dutd07_i3co2w2978g = ~y1l45u9lhj0l_z8ry7s_4;   
  wire dyryg74kmrh9updbc = ~mw8igz4fx7cd12mg;
  wire m_ycdgre0ehecyndcdud;
  wire qaorcvxc0rrtus17;

generate
if (ZEROCYC_RSP == 1) begin:lt6a02wdfsh074vb99
  ux607_gnrl_bypbuf #(
          .DP  (FIFO_OUTS_NUM),
          .DW  (2)
  )  yfou_i2ygia41t_nhj75iftch(
      .i_vld(cyags_6gth1ma8wjx896),
      .i_rdy(y1l45u9lhj0l_z8ry7s_4),
      .i_dat({skq4j6qdkmbvs1k9lufa,rg2wqryxlxihjmh4v}),
      .o_vld(mw8igz4fx7cd12mg),
      .o_rdy(x43j9vfjtxotxnel20jv),
      .o_dat({m_ycdgre0ehecyndcdud,qaorcvxc0rrtus17}),

      .clk(clk),
      .rst_n(rst_n)
  );
end
else begin :gueeox0z90gbmx7
  if(FIFO_OUTS_NUM == 1) begin:axug194an99bql_f8e
      ux607_gnrl_pipe_stage #(
          .CUT_READY(FIFO_CUT_READY),
          .DP(1),
          .DW(2)
      ) x3q7avo94mkdoysyezegqn (
          .i_vld(cyags_6gth1ma8wjx896),
          .i_rdy(y1l45u9lhj0l_z8ry7s_4),
          .i_dat({skq4j6qdkmbvs1k9lufa,rg2wqryxlxihjmh4v}),
          .o_vld(mw8igz4fx7cd12mg),
          .o_rdy(x43j9vfjtxotxnel20jv),
          .o_dat({m_ycdgre0ehecyndcdud,qaorcvxc0rrtus17}),

          .clk(clk),
          .rst_n(rst_n)
      );
  end
  else begin:ayrjh6ok2h5s8a98q
      ux607_gnrl_fifo #(
          .CUT_READY (FIFO_CUT_READY),
          .MSKO      (0),
          .DP  (FIFO_OUTS_NUM),
          .DW  (2)
      )  x3q7avo94mkdoysyezegqn(
          .i_vld(cyags_6gth1ma8wjx896),
          .i_rdy(y1l45u9lhj0l_z8ry7s_4),
          .i_dat({skq4j6qdkmbvs1k9lufa,rg2wqryxlxihjmh4v}),
          .o_vld(mw8igz4fx7cd12mg),
          .o_rdy(x43j9vfjtxotxnel20jv),
          .o_dat({m_ycdgre0ehecyndcdud,qaorcvxc0rrtus17}),

          .clk(clk),
          .rst_n(rst_n)
      );
  end
end
endgenerate

  wire             n6uge82egdm_cw6aokw48;
  wire             ajfmeb_o6x5e11tp7ab4klcani;  
  wire             jpp4f0jj2yb2ud0b0stpyvy_zt;
  wire             rynrau0l_icpe8ztaqtcn;
  wire             vxv6yqxral28zu3xvv7oc;
  wire             kpz5lejuqu2xxcuj9opfwmau9nq;

  wire jm3dko31uqsmxc06awx4  = o_icb_cmd_valid & o_icb_cmd_ready;

  generate
  if (LATE_READY) begin :j8688n5of827
  assign rynrau0l_icpe8ztaqtcn = skq4j6qdkmbvs1k9lufa & jm3dko31uqsmxc06awx4 & (~n6uge82egdm_cw6aokw48);
  assign vxv6yqxral28zu3xvv7oc = skq4j6qdkmbvs1k9lufa & jm3dko31uqsmxc06awx4 & n6uge82egdm_cw6aokw48;
  assign kpz5lejuqu2xxcuj9opfwmau9nq = skq4j6qdkmbvs1k9lufa ? n6uge82egdm_cw6aokw48 : 1'b1;


  assign o_icb_cmd_valid = (~dutd07_i3co2w2978g) & i_icb_cmd_valid;
  assign o_icb_cmd_addr  = (skq4j6qdkmbvs1k9lufa & n6uge82egdm_cw6aokw48) ? {i_icb_cmd_addr[X_W-1:3],3'b100}
                                                                               : i_icb_cmd_addr;
  assign o_icb_cmd_read  = i_icb_cmd_read;                      
  assign o_icb_cmd_wdata = (skq4j6qdkmbvs1k9lufa & n6uge82egdm_cw6aokw48) ? i_icb_cmd_wdata[X_W-1:Y_W] : 
                           (rg2wqryxlxihjmh4v                       ) ? i_icb_cmd_wdata[X_W-1:Y_W] :
                                                                     i_icb_cmd_wdata[Y_W-1:0]
                                                                   ;
  assign o_icb_cmd_wmask = (skq4j6qdkmbvs1k9lufa & n6uge82egdm_cw6aokw48) ? i_icb_cmd_wmask[(X_W/8-1):(Y_W/8)] : 
                           (rg2wqryxlxihjmh4v                       ) ? i_icb_cmd_wmask[(X_W/8-1):(Y_W/8)] : 
                                                                     i_icb_cmd_wmask[(Y_W/8-1):0]
                                                                   ;
  assign o_icb_cmd_usr  = i_icb_cmd_usr;
  assign o_icb_cmd_beat = i_icb_cmd_beat[1:0];
  assign o_icb_cmd_size = skq4j6qdkmbvs1k9lufa ? 2'b10 : i_icb_cmd_size;
  end
  else begin :hmk5jwx4rw0ec10m
  assign rynrau0l_icpe8ztaqtcn     = skq4j6qdkmbvs1k9lufa      & jm3dko31uqsmxc06awx4;
  assign vxv6yqxral28zu3xvv7oc     = n6uge82egdm_cw6aokw48  & jm3dko31uqsmxc06awx4;
  assign kpz5lejuqu2xxcuj9opfwmau9nq = !n6uge82egdm_cw6aokw48; 

  wire             s8v498gn7d3w8gqr9q8;
  wire [AW-1:3]    tl3408q3kji1gyhpe9b12;
  wire [Y_W-1:0]   g306qzqxu0m2b5_se_w;
  wire [Y_W/8-1:0] ab9u834d1_y168o5ot4up;
  wire [USR_W-1:0] tv39u69w2zg7qly4kq_32r;
  wire [1:0]       g0mruv4nlr6uz8ghmp4n6lb;
  ux607_gnrl_dfflr #(1)     a7e04grbsp51zchg   (rynrau0l_icpe8ztaqtcn, i_icb_cmd_read, s8v498gn7d3w8gqr9q8, clk, rst_n);
  ux607_gnrl_dfflr #(AW-3)  i5g67bnjzxc1sgz3rnl   (rynrau0l_icpe8ztaqtcn, i_icb_cmd_addr[AW-1:3], tl3408q3kji1gyhpe9b12, clk, rst_n);
  ux607_gnrl_dfflr #(Y_W)   f3m0unt8ok7ruf2wt41x  (rynrau0l_icpe8ztaqtcn, i_icb_cmd_wdata[X_W-1:Y_W], g306qzqxu0m2b5_se_w, clk, rst_n);
  ux607_gnrl_dfflr #(Y_W/8) hrbnxkhon_lowwlfo5fi5s  (rynrau0l_icpe8ztaqtcn, i_icb_cmd_wmask[X_W/8-1:Y_W/8], ab9u834d1_y168o5ot4up, clk, rst_n);
  ux607_gnrl_dfflr #(USR_W) crqfamud9ajdv84    (rynrau0l_icpe8ztaqtcn, i_icb_cmd_usr, tv39u69w2zg7qly4kq_32r, clk, rst_n);
  ux607_gnrl_dfflr #(2)     qyaqvpwar993xu710o8   (rynrau0l_icpe8ztaqtcn, i_icb_cmd_beat[1:0], g0mruv4nlr6uz8ghmp4n6lb, clk, rst_n);


  assign o_icb_cmd_valid = (~dutd07_i3co2w2978g) & i_icb_cmd_valid || n6uge82egdm_cw6aokw48;

  assign o_icb_cmd_addr = n6uge82egdm_cw6aokw48 ? {tl3408q3kji1gyhpe9b12[AW-1:3],3'b100}
                                              :  i_icb_cmd_addr;
  assign o_icb_cmd_read = n6uge82egdm_cw6aokw48 ? s8v498gn7d3w8gqr9q8
                                              : i_icb_cmd_read;                      
  assign o_icb_cmd_wdata = n6uge82egdm_cw6aokw48 ? g306qzqxu0m2b5_se_w : 
                           rg2wqryxlxihjmh4v      ? i_icb_cmd_wdata[X_W-1:Y_W] :
                                                 i_icb_cmd_wdata[Y_W-1:0];

  assign o_icb_cmd_wmask = n6uge82egdm_cw6aokw48 ? ab9u834d1_y168o5ot4up : 
                           rg2wqryxlxihjmh4v      ? i_icb_cmd_wmask[(X_W/8-1):(Y_W/8)] : 
                                                 i_icb_cmd_wmask[(Y_W/8-1):0];

  assign o_icb_cmd_usr  = n6uge82egdm_cw6aokw48 ? tv39u69w2zg7qly4kq_32r
                                              : i_icb_cmd_usr;
  assign o_icb_cmd_beat = n6uge82egdm_cw6aokw48 ? g0mruv4nlr6uz8ghmp4n6lb
                                              : i_icb_cmd_beat[1:0];
  assign o_icb_cmd_size = (skq4j6qdkmbvs1k9lufa || n6uge82egdm_cw6aokw48)  ? 2'b10 : i_icb_cmd_size;
  end
  endgenerate

  assign ajfmeb_o6x5e11tp7ab4klcani = rynrau0l_icpe8ztaqtcn | vxv6yqxral28zu3xvv7oc;  
  assign jpp4f0jj2yb2ud0b0stpyvy_zt = rynrau0l_icpe8ztaqtcn & (~vxv6yqxral28zu3xvv7oc);
  ux607_gnrl_dfflr #(1)     y8t7_x8t91kcrz98gbbz  (ajfmeb_o6x5e11tp7ab4klcani, jpp4f0jj2yb2ud0b0stpyvy_zt, n6uge82egdm_cw6aokw48, clk, rst_n);

  wire n9lr4wk9te5d7rq1gklvi  = o_icb_rsp_valid & o_icb_rsp_ready;
  wire zpru6vd3zypnlwdarcg8  = i_icb_rsp_valid & i_icb_rsp_ready;

  wire maw39vt1c25mcyrh4wxm9g;
  wire q0kjpsn6gup6dnnoir08k = m_ycdgre0ehecyndcdud & n9lr4wk9te5d7rq1gklvi & (~maw39vt1c25mcyrh4wxm9g);
  wire f_9rnxzpm4fz5pptm3owiinepb = m_ycdgre0ehecyndcdud & n9lr4wk9te5d7rq1gklvi & maw39vt1c25mcyrh4wxm9g;
  wire miei12dtt5oc3lb1iduifvne = q0kjpsn6gup6dnnoir08k | f_9rnxzpm4fz5pptm3owiinepb;  
  wire kb380o8k74e8gwhc1ulhj = q0kjpsn6gup6dnnoir08k & (~f_9rnxzpm4fz5pptm3owiinepb);
  ux607_gnrl_dfflr #(1) egg_sec15307xgnxhp18gfeocj(miei12dtt5oc3lb1iduifvne, kb380o8k74e8gwhc1ulhj, maw39vt1c25mcyrh4wxm9g, clk, rst_n);



  wire c_iwfr81byy1o33srnue7 = m_ycdgre0ehecyndcdud &  n9lr4wk9te5d7rq1gklvi & (~maw39vt1c25mcyrh4wxm9g);
  wire [Y_W-1:0] mhjxzdjjzzimwz3fqigi7zujmdkki = o_icb_rsp_rdata[Y_W-1:0];
  wire [Y_W-1:0] s9qasvbuqbbeavzvhh2iuww3phepa; 
  ux607_gnrl_dfflr #(Y_W) m0rm43qj_27eg13nhc9l7rkuc298a4jc(c_iwfr81byy1o33srnue7, mhjxzdjjzzimwz3fqigi7zujmdkki, s9qasvbuqbbeavzvhh2iuww3phepa, clk, rst_n);

  wire l4cn27lciatju8nnkgrfavg0w = o_icb_rsp_err;
  wire sa9f3o18lj6m1utkqlfdo2w; 
  ux607_gnrl_dfflr #(1) icq8_w9fcb46g_fa3jrvlt0krh(c_iwfr81byy1o33srnue7, l4cn27lciatju8nnkgrfavg0w, sa9f3o18lj6m1utkqlfdo2w, clk, rst_n);


  wire uimr_wbkcfb6lws3k5a7 = maw39vt1c25mcyrh4wxm9g; 

  assign i_icb_cmd_ready = (~dutd07_i3co2w2978g) & kpz5lejuqu2xxcuj9opfwmau9nq & o_icb_cmd_ready;  
  assign o_icb_cmd_burst = 3'b0; 
  assign o_icb_cmd_lock = 1'b0;
  assign o_icb_cmd_excl = 1'b0;


  wire zvucw4f7m96zfihivkrut = m_ycdgre0ehecyndcdud ? maw39vt1c25mcyrh4wxm9g : 1'b1;


  assign i_icb_rsp_valid =  zvucw4f7m96zfihivkrut & o_icb_rsp_valid;
  assign i_icb_rsp_rdata = uimr_wbkcfb6lws3k5a7 ? {o_icb_rsp_rdata, s9qasvbuqbbeavzvhh2iuww3phepa} : 
                           qaorcvxc0rrtus17       ? {o_icb_rsp_rdata, {Y_W{1'b0}}}              :
                                                  {{Y_W{1'b0}}, o_icb_rsp_rdata}
                                                ;
  assign o_icb_rsp_ready = i_icb_rsp_ready; 
  assign i_icb_rsp_err   = uimr_wbkcfb6lws3k5a7 ? |{sa9f3o18lj6m1utkqlfdo2w, o_icb_rsp_err} : o_icb_rsp_err;
  assign i_icb_rsp_excl_ok = 1'b0;
  assign i_icb_rsp_usr   = o_icb_rsp_usr;


endmodule







module ux607_gnrl_icb_splt # (
  parameter AW = 32,
  parameter DW = 64,
  parameter USE_ALL_READY = 0,

  parameter FIFO_OUTS_NUM = 8,
  parameter FIFO_CUT_READY = 0,

  parameter SPLT_NUM = 4,
  parameter SPLT_PTR_1HOT = 1,

  parameter SPLT_PTR_W = 4,
  parameter ALLOW_DIFF = 1,
  parameter ALLOW_0CYCL_RSP = 1,
  parameter VLD_MSK_PAYLOAD = 0,
  parameter USR_W = 1 
) (
  input  [SPLT_NUM-1:0] i_icb_splt_indic,        

  output splt_active,

  input  i_icb_cmd_valid, 
  output i_icb_cmd_ready, 
  input             i_icb_cmd_read, 
  input  [AW-1:0]   i_icb_cmd_addr, 
  input  [DW-1:0]   i_icb_cmd_wdata, 
  input  [(DW/8-1):0] i_icb_cmd_wmask,
  input  [2:0]      i_icb_cmd_burst,
  input  [1:0]      i_icb_cmd_beat,
  input             i_icb_cmd_lock,
  input             i_icb_cmd_excl,
  input  [1:0]      i_icb_cmd_size,
  input  [USR_W-1:0]i_icb_cmd_usr,

  output i_icb_rsp_valid, 
  input  i_icb_rsp_ready, 
  output i_icb_rsp_err,
  output i_icb_rsp_excl_ok,
  output [DW-1:0] i_icb_rsp_rdata, 
  output [USR_W-1:0] i_icb_rsp_usr, 

  input  [SPLT_NUM*1-1:0]    o_bus_icb_cmd_ready, 
  output [SPLT_NUM*1-1:0]    o_bus_icb_cmd_valid, 
  output [SPLT_NUM*1-1:0]    o_bus_icb_cmd_read, 
  output [SPLT_NUM*AW-1:0]   o_bus_icb_cmd_addr, 
  output [SPLT_NUM*DW-1:0]   o_bus_icb_cmd_wdata, 
  output [(SPLT_NUM*DW/8-1):0] o_bus_icb_cmd_wmask,
  output [SPLT_NUM*3-1:0]    o_bus_icb_cmd_burst,
  output [SPLT_NUM*2-1:0]    o_bus_icb_cmd_beat,
  output [SPLT_NUM*1-1:0]    o_bus_icb_cmd_lock,
  output [SPLT_NUM*1-1:0]    o_bus_icb_cmd_excl,
  output [SPLT_NUM*2-1:0]    o_bus_icb_cmd_size,
  output [SPLT_NUM*USR_W-1:0]o_bus_icb_cmd_usr,

  input  [SPLT_NUM*1-1:0]  o_bus_icb_rsp_valid, 
  output [SPLT_NUM*1-1:0]  o_bus_icb_rsp_ready, 
  input  [SPLT_NUM*1-1:0]  o_bus_icb_rsp_err,
  input  [SPLT_NUM*1-1:0]  o_bus_icb_rsp_excl_ok,
  input  [SPLT_NUM*DW-1:0] o_bus_icb_rsp_rdata, 
  input  [SPLT_NUM*USR_W-1:0] o_bus_icb_rsp_usr, 

  input  clk,  
  input  rst_n
  );


    wire pjisa4vlo9u0rtnt1whf8;       

generate 
  if(SPLT_NUM == 1) begin:zyyh4gsu1mivdipl43
    assign i_icb_cmd_ready     = o_bus_icb_cmd_ready; 
    assign o_bus_icb_cmd_valid = i_icb_cmd_valid; 
    assign o_bus_icb_cmd_read  = i_icb_cmd_read ; 
    assign o_bus_icb_cmd_addr  = i_icb_cmd_addr ; 
    assign o_bus_icb_cmd_wdata = i_icb_cmd_wdata; 
    assign o_bus_icb_cmd_wmask = i_icb_cmd_wmask;
    assign o_bus_icb_cmd_burst = i_icb_cmd_burst;
    assign o_bus_icb_cmd_beat  = i_icb_cmd_beat ;
    assign o_bus_icb_cmd_lock  = i_icb_cmd_lock ;
    assign o_bus_icb_cmd_excl  = i_icb_cmd_excl ;
    assign o_bus_icb_cmd_size  = i_icb_cmd_size ;
    assign o_bus_icb_cmd_usr   = i_icb_cmd_usr  ;

    assign o_bus_icb_rsp_ready = i_icb_rsp_ready; 
    assign i_icb_rsp_valid     = o_bus_icb_rsp_valid; 
    assign i_icb_rsp_err       = o_bus_icb_rsp_err  ;
    assign i_icb_rsp_excl_ok   = o_bus_icb_rsp_excl_ok  ;
    assign i_icb_rsp_rdata     = o_bus_icb_rsp_rdata;
    assign i_icb_rsp_usr       = o_bus_icb_rsp_usr;

    assign pjisa4vlo9u0rtnt1whf8    = 1'b1;       
  end
  else begin:x_be1k_xipx5pgftxq1

    genvar i;
    genvar nzd5e;
    integer j;

    wire [SPLT_NUM-1:0] me2s8h5yw65ail5; 
    wire [SPLT_NUM-1:0] dtyl4o87hqhm03wj57; 

    wire            xiyx61_yd314uojrls [SPLT_NUM-1:0]; 
    wire [AW-1:0]   k68zoq6vpu0olvs99f [SPLT_NUM-1:0]; 
    wire [DW-1:0]   m63rlc2ixlaphiq[SPLT_NUM-1:0]; 
    wire [(DW/8-1):0] drdtbfa60cpn5ihc[SPLT_NUM-1:0];
    wire [2:0]      rnrkzgtukyiil52jqbp7[SPLT_NUM-1:0];
    wire [1:0]      wta_51f6oa6zy5t [SPLT_NUM-1:0];
    wire            da5mm7z1qer9hx385ck [SPLT_NUM-1:0];
    wire            tg7q7ezs0lgu3bv36l4 [SPLT_NUM-1:0];
    wire [1:0]      hycxa49k327vm1ncjh [SPLT_NUM-1:0];
    wire [USR_W-1:0]vzw7nivk4j2idd  [SPLT_NUM-1:0];

    wire [SPLT_NUM-1:0] mg6xxata423v5aaikz4v; 
    wire [SPLT_NUM-1:0] yuew3x5jdkrr87g; 
    wire [SPLT_NUM-1:0] nkx3bwv604xt1  ;
    wire [SPLT_NUM-1:0] db9kwedxc8ekbwcenl8s9  ;
    wire [DW-1:0] lbvrc0jeu6t70bw  [SPLT_NUM-1:0];
    wire [USR_W-1:0] wxjl9xtjejiyjn1 [SPLT_NUM-1:0];

    wire [SPLT_NUM-1:0] t20655hp_wcz_dzflgifw9xah_2g1 [SPLT_NUM-1:0];

    wire yuy8ms35qeu8m4f4rwz9wpc;

    wire djmbzt1843lpcet2xr1d1b;
    wire gp0lafw7tngumfeqku5;
    wire m3ho2mulswsyi6r_r;

    wire [SPLT_PTR_W-1:0] gelhdm56emraair2nv;

    wire jxqrb_9po4b1mxj0al90g;
    wire kbtixer0amhrz2dzvhe;
    wire wr80zcrpu3t413geuk;
    wire nhqlx69jse016ld9w87kjm7;
    wire [SPLT_PTR_W-1:0] ibsurazp9nyl3c3a;
    wire [SPLT_PTR_W-1:0] uogk6x1xf6j9v5w;

    wire ns807okp2nn628yu3u;       
    reg [SPLT_PTR_W-1:0] syio1sc28rnpat8cala;

    wire xp2vrz0kfqlv21fb4ce;
    wire l60xdkct0g8mjsykqp71f9ti;

    wire gyig5xdgz_v1h18gkcrz_j1; 
    wire jcxgswikiw_3vq65p8jdb;


    for(i = 0; i < SPLT_NUM; i = i+1)
    begin:s9dy2pie07n9wcw_a
      assign dtyl4o87hqhm03wj57[i]                             = o_bus_icb_cmd_ready[(i+1)*1     -1 : (i)*1     ]; 
      assign o_bus_icb_cmd_valid[(i+1)*1     -1 : i*1     ] = me2s8h5yw65ail5[i];
      assign o_bus_icb_cmd_read [(i+1)*1     -1 : i*1     ] = xiyx61_yd314uojrls [i];
      assign o_bus_icb_cmd_addr [(i+1)*AW    -1 : i*AW    ] = k68zoq6vpu0olvs99f [i];
      assign o_bus_icb_cmd_wdata[(i+1)*DW    -1 : i*DW    ] = m63rlc2ixlaphiq[i];
      assign o_bus_icb_cmd_wmask[(i+1)*(DW/8)-1 : i*(DW/8)] = drdtbfa60cpn5ihc[i];
      assign o_bus_icb_cmd_burst[(i+1)*3     -1 : i*3     ] = rnrkzgtukyiil52jqbp7[i];
      assign o_bus_icb_cmd_beat [(i+1)*2     -1 : i*2     ] = wta_51f6oa6zy5t [i];
      assign o_bus_icb_cmd_lock [(i+1)*1     -1 : i*1     ] = da5mm7z1qer9hx385ck [i];
      assign o_bus_icb_cmd_excl [(i+1)*1     -1 : i*1     ] = tg7q7ezs0lgu3bv36l4 [i];
      assign o_bus_icb_cmd_size [(i+1)*2     -1 : i*2     ] = hycxa49k327vm1ncjh [i];
      assign o_bus_icb_cmd_usr  [(i+1)*USR_W -1 : i*USR_W ] = vzw7nivk4j2idd  [i];

      assign o_bus_icb_rsp_ready[(i+1)*1-1 :i*1 ] = yuew3x5jdkrr87g[i]; 
      assign mg6xxata423v5aaikz4v[i]                   = o_bus_icb_rsp_valid[(i+1)*1-1 :i*1 ]; 
      assign nkx3bwv604xt1  [i]                   = o_bus_icb_rsp_err  [(i+1)*1-1 :i*1 ];
      assign db9kwedxc8ekbwcenl8s9  [i]               = o_bus_icb_rsp_excl_ok  [(i+1)*1-1 :i*1 ];
      assign lbvrc0jeu6t70bw[i]                   = o_bus_icb_rsp_rdata[(i+1)*DW-1:i*DW];
      assign wxjl9xtjejiyjn1  [i]                   = o_bus_icb_rsp_usr  [(i+1)*USR_W-1:i*USR_W];
    end





    if(USE_ALL_READY == 1) begin:u393d5_r1r_efen5ak
      assign yuy8ms35qeu8m4f4rwz9wpc = (&dtyl4o87hqhm03wj57);
    end
    else begin:wpjtermhv2o0ch3tw83sqm
      reg  kozxvnx2573ftzsqsd8mov36c;
      always @ (*) begin : lh82_td_rnhybm4y5zqrzzru2jbcd
        kozxvnx2573ftzsqsd8mov36c = 1'b0;
          for(j = 0; j < SPLT_NUM; j = j+1) begin
            kozxvnx2573ftzsqsd8mov36c = kozxvnx2573ftzsqsd8mov36c | (i_icb_splt_indic[j] & dtyl4o87hqhm03wj57[j]);
          end
      end
      assign yuy8ms35qeu8m4f4rwz9wpc = kozxvnx2573ftzsqsd8mov36c;
    end

    assign xp2vrz0kfqlv21fb4ce = yuy8ms35qeu8m4f4rwz9wpc;

    if(ALLOW_DIFF == 1) begin:ec1olcpuy6vur03
       assign l60xdkct0g8mjsykqp71f9ti = i_icb_cmd_valid     & (~ns807okp2nn628yu3u);
       assign i_icb_cmd_ready     = xp2vrz0kfqlv21fb4ce & (~ns807okp2nn628yu3u);
    end
    else begin:djynwdimydwsxgit7_bqy7


       wire csr6ull36_jpsgz3o2al = (~pjisa4vlo9u0rtnt1whf8) & (~(uogk6x1xf6j9v5w == ibsurazp9nyl3c3a));
       assign l60xdkct0g8mjsykqp71f9ti = i_icb_cmd_valid     & (~csr6ull36_jpsgz3o2al) & (~ns807okp2nn628yu3u);
       assign i_icb_cmd_ready     = xp2vrz0kfqlv21fb4ce & (~csr6ull36_jpsgz3o2al) & (~ns807okp2nn628yu3u);
    end


    if(SPLT_PTR_1HOT == 1) begin:g8c3ly7vmyb0r
       always @ (*) begin : yzw7sa9icrhk0xwc1mp1rw7v
         syio1sc28rnpat8cala = i_icb_splt_indic;
       end
    end
    else begin:hsawddfz6jvn5kzgl
       always @ (*) begin : yzw7sa9icrhk0xwc1mp1rw7v
         syio1sc28rnpat8cala = {SPLT_PTR_W{1'b0}};
         for(j = 0; j < SPLT_NUM; j = j+1) begin
           syio1sc28rnpat8cala = syio1sc28rnpat8cala | ({SPLT_PTR_W{i_icb_splt_indic[j]}} & $unsigned(j[SPLT_PTR_W-1:0]));
         end
       end
    end

    assign gp0lafw7tngumfeqku5 = i_icb_cmd_valid & i_icb_cmd_ready;
    assign m3ho2mulswsyi6r_r = i_icb_rsp_valid & i_icb_rsp_ready;

    if(ALLOW_0CYCL_RSP == 1) begin: ywf24098_gi8bfyn2w
        assign djmbzt1843lpcet2xr1d1b = pjisa4vlo9u0rtnt1whf8 & gp0lafw7tngumfeqku5 & m3ho2mulswsyi6r_r;
        assign gelhdm56emraair2nv = pjisa4vlo9u0rtnt1whf8 ? uogk6x1xf6j9v5w : ibsurazp9nyl3c3a;

        assign i_icb_rsp_valid     = jcxgswikiw_3vq65p8jdb;
        assign gyig5xdgz_v1h18gkcrz_j1 = i_icb_rsp_ready;
    end
    else begin: ss_g5sktytsbln200rqk
        assign djmbzt1843lpcet2xr1d1b = 1'b0;
        assign gelhdm56emraair2nv = ibsurazp9nyl3c3a;
        assign i_icb_rsp_valid     = (~pjisa4vlo9u0rtnt1whf8) & jcxgswikiw_3vq65p8jdb;
        assign gyig5xdgz_v1h18gkcrz_j1 = (~pjisa4vlo9u0rtnt1whf8) & i_icb_rsp_ready;
    end

    assign jxqrb_9po4b1mxj0al90g = gp0lafw7tngumfeqku5 & (~djmbzt1843lpcet2xr1d1b);
    assign ns807okp2nn628yu3u    = (~wr80zcrpu3t413geuk);
    assign nhqlx69jse016ld9w87kjm7 = m3ho2mulswsyi6r_r & (~djmbzt1843lpcet2xr1d1b);
    assign pjisa4vlo9u0rtnt1whf8   = (~kbtixer0amhrz2dzvhe);

    assign uogk6x1xf6j9v5w   = syio1sc28rnpat8cala;

    if(FIFO_OUTS_NUM == 1) begin:axug194an99bql_f8e
      ux607_gnrl_pipe_stage # (
        .CUT_READY (FIFO_CUT_READY),
        .DP  (1),
        .DW  (SPLT_PTR_W)
      ) ahkryar1lc8lsjv5v1c_6ce6 (
        .i_vld(jxqrb_9po4b1mxj0al90g),
        .i_rdy(wr80zcrpu3t413geuk),
        .i_dat(uogk6x1xf6j9v5w ),
        .o_vld(kbtixer0amhrz2dzvhe),
        .o_rdy(nhqlx69jse016ld9w87kjm7),  
        .o_dat(ibsurazp9nyl3c3a ),  

        .clk  (clk),
        .rst_n(rst_n)
      );

    end
    else begin: ayrjh6ok2h5s8a98q
      ux607_gnrl_fifo # (
        .CUT_READY (FIFO_CUT_READY),
        .MSKO      (0),
        .DP  (FIFO_OUTS_NUM),
        .DW  (SPLT_PTR_W)
      ) ahkryar1lc8lsjv5v1c_6ce6 (
        .i_vld(jxqrb_9po4b1mxj0al90g),
        .i_rdy(wr80zcrpu3t413geuk),
        .i_dat(uogk6x1xf6j9v5w ),
        .o_vld(kbtixer0amhrz2dzvhe),
        .o_rdy(nhqlx69jse016ld9w87kjm7),  
        .o_dat(ibsurazp9nyl3c3a ),  

        .clk  (clk),
        .rst_n(rst_n)
      );
    end



    for(i = 0; i < SPLT_NUM; i = i+1)
    begin:dud1pqnswdrsex1ymzb4xux

      for(nzd5e = 0; nzd5e < SPLT_NUM; nzd5e = nzd5e+1)
      begin:ldo1tu4qfgp98k1pwxo5_a4dbwpb
         if(i == nzd5e) begin: c_qzobhog39
           assign t20655hp_wcz_dzflgifw9xah_2g1[i][nzd5e] = 1'b1;
         end
         else begin: t2dfftioa6dhr9y
           assign t20655hp_wcz_dzflgifw9xah_2g1[i][nzd5e] = dtyl4o87hqhm03wj57[nzd5e];
         end
      end

      if(USE_ALL_READY == 1) begin:u393d5_r1r_efen5ak
         assign me2s8h5yw65ail5[i] = i_icb_splt_indic[i] & l60xdkct0g8mjsykqp71f9ti & (&t20655hp_wcz_dzflgifw9xah_2g1[i]);         
      end
      else begin:wpjtermhv2o0ch3tw83sqm
         assign me2s8h5yw65ail5[i] = i_icb_splt_indic[i] & l60xdkct0g8mjsykqp71f9ti;         
      end
      if(VLD_MSK_PAYLOAD == 0) begin: uxdupicf1j93739ktjcbjka_3fd
          assign xiyx61_yd314uojrls [i] = i_icb_cmd_read ;
          assign k68zoq6vpu0olvs99f [i] = i_icb_cmd_addr ;
          assign m63rlc2ixlaphiq[i] = i_icb_cmd_wdata;
          assign drdtbfa60cpn5ihc[i] = i_icb_cmd_wmask;
          assign rnrkzgtukyiil52jqbp7[i] = i_icb_cmd_burst;
          assign wta_51f6oa6zy5t [i] = i_icb_cmd_beat ;
          assign da5mm7z1qer9hx385ck [i] = i_icb_cmd_lock ;
          assign tg7q7ezs0lgu3bv36l4 [i] = i_icb_cmd_excl ;
          assign hycxa49k327vm1ncjh [i] = i_icb_cmd_size ;
          assign vzw7nivk4j2idd  [i] = i_icb_cmd_usr  ;
      end
      else begin: j5_ymxr1x20ah4dcw0ypt3
          assign xiyx61_yd314uojrls [i] = {1    {me2s8h5yw65ail5[i]}} & i_icb_cmd_read ;
          assign k68zoq6vpu0olvs99f [i] = {AW   {me2s8h5yw65ail5[i]}} & i_icb_cmd_addr ;
          assign m63rlc2ixlaphiq[i] = {DW   {me2s8h5yw65ail5[i]}} & i_icb_cmd_wdata;
          assign drdtbfa60cpn5ihc[i] = {DW/8 {me2s8h5yw65ail5[i]}} & i_icb_cmd_wmask;
          assign rnrkzgtukyiil52jqbp7[i] = {3    {me2s8h5yw65ail5[i]}} & i_icb_cmd_burst;
          assign wta_51f6oa6zy5t [i] = {2    {me2s8h5yw65ail5[i]}} & i_icb_cmd_beat ;
          assign da5mm7z1qer9hx385ck [i] = {1    {me2s8h5yw65ail5[i]}} & i_icb_cmd_lock ;
          assign tg7q7ezs0lgu3bv36l4 [i] = {1    {me2s8h5yw65ail5[i]}} & i_icb_cmd_excl ;
          assign hycxa49k327vm1ncjh [i] = {2    {me2s8h5yw65ail5[i]}} & i_icb_cmd_size ;
          assign vzw7nivk4j2idd  [i] = {USR_W{me2s8h5yw65ail5[i]}} & i_icb_cmd_usr  ;
      end
    end





    if(SPLT_PTR_1HOT == 1) begin:saq1sh16t3q3w7y7_hl5_

        for(i = 0; i < SPLT_NUM; i = i+1)
        begin:y5k3_r0ccgeuxsjc688hv5o
          assign yuew3x5jdkrr87g[i] = (gelhdm56emraair2nv[i] & gyig5xdgz_v1h18gkcrz_j1);
        end

        assign jcxgswikiw_3vq65p8jdb = |({SPLT_PTR_W{mg6xxata423v5aaikz4v}} & gelhdm56emraair2nv);


        reg p7ejtrejd40jkasujx;
        reg s8izkgasvh31dc67zdh_1dz2;
        reg [DW-1:0] ddeyuzlw7mltu69morzvy7; 
        reg [USR_W-1:0] iiafqgjhrh58_l69wwni; 

        always @ (*) begin : oe9tqryz7wdpms9syhz
          p7ejtrejd40jkasujx   = 1'b0;
          s8izkgasvh31dc67zdh_1dz2   = 1'b0;
          ddeyuzlw7mltu69morzvy7 = {DW   {1'b0}};
          iiafqgjhrh58_l69wwni   = {USR_W{1'b0}};
          for(j = 0; j < SPLT_NUM; j = j+1) begin
            p7ejtrejd40jkasujx     = p7ejtrejd40jkasujx     | (       gelhdm56emraair2nv[j]   & nkx3bwv604xt1[j]);
            s8izkgasvh31dc67zdh_1dz2 = s8izkgasvh31dc67zdh_1dz2 | (       gelhdm56emraair2nv[j]   & db9kwedxc8ekbwcenl8s9[j]);
            ddeyuzlw7mltu69morzvy7   = ddeyuzlw7mltu69morzvy7   | ({DW   {gelhdm56emraair2nv[j]}} & lbvrc0jeu6t70bw[j]);
            iiafqgjhrh58_l69wwni     = iiafqgjhrh58_l69wwni     | ({USR_W{gelhdm56emraair2nv[j]}} & wxjl9xtjejiyjn1[j]);
          end
        end

        assign i_icb_rsp_err   = p7ejtrejd40jkasujx  ;
        assign i_icb_rsp_excl_ok   = s8izkgasvh31dc67zdh_1dz2  ;
        assign i_icb_rsp_rdata = ddeyuzlw7mltu69morzvy7;
        assign i_icb_rsp_usr   = iiafqgjhrh58_l69wwni  ;

    end
    else begin:n9cey7fhfge6_6xc7jpn

        for(i = 0; i < SPLT_NUM; i = i+1)
        begin:y5k3_r0ccgeuxsjc688hv5o
          assign yuew3x5jdkrr87g[i] = (gelhdm56emraair2nv == i[SPLT_PTR_W-1:0]) & gyig5xdgz_v1h18gkcrz_j1;
        end

        assign jcxgswikiw_3vq65p8jdb = mg6xxata423v5aaikz4v[gelhdm56emraair2nv]; 


        assign i_icb_rsp_err     = nkx3bwv604xt1    [gelhdm56emraair2nv]; 
        assign i_icb_rsp_excl_ok = db9kwedxc8ekbwcenl8s9[gelhdm56emraair2nv]; 
        assign i_icb_rsp_rdata   = lbvrc0jeu6t70bw  [gelhdm56emraair2nv]; 
        assign i_icb_rsp_usr     = wxjl9xtjejiyjn1    [gelhdm56emraair2nv]; 
    end

  end
  endgenerate 

  assign splt_active = (i_icb_cmd_valid) | (~pjisa4vlo9u0rtnt1whf8);

endmodule














































































































































































































































































































module ux607_gnrl_icb2ahbl
  #(
    parameter SUPPORT_LOCK = 0,


    parameter MON_DATA_WIDTH = 2,
    parameter AW = 32,
    parameter DW = 32 
    )
  (

  input              icb_cmd_valid, 
  output             icb_cmd_ready, 
  input              icb_cmd_read, 
  input  [AW-1:0]    icb_cmd_addr, 
  input  [DW-1:0]    icb_cmd_wdata, 
  input  [(DW/8-1):0]  icb_cmd_wmask,
  input  [1:0]       icb_cmd_size,
  input              icb_cmd_lock,
  input              icb_cmd_excl,
  input  [3-1:0]     icb_cmd_burst, 
  input  [3:0]       icb_cmd_hprot, 
  input  [1:0]       icb_cmd_attri, 
  input              icb_cmd_dmode, 
  input              icb_cmd_hseq,

  output             icb_rsp_valid, 

  output             icb_rsp_err,
  output             icb_rsp_excl_ok,
  output [DW-1:0]    icb_rsp_rdata, 

  output [1:0]       ahbl_htrans,   
  output             ahbl_hwrite,   
  output [AW    -1:0]ahbl_haddr,    
  output [2:0]       ahbl_hsize,    
  output             ahbl_hlock,   
  output             ahbl_hexcl,   
  output [2:0]       ahbl_hburst,   
  output [DW    -1:0]ahbl_hwdata,   
  output [3:0]       ahbl_hprot, 
  output [1:0]       ahbl_hattri,
  output [1:0]       ahbl_master,
  input  [DW    -1:0]ahbl_hrdata,   
  input  [1:0]       ahbl_hresp,    
  input              ahbl_hresp_exok,    
  input              ahbl_hready,   

  input              bus_clk_en,

  output             icb2ahbl_pend_active,

  input              clk,          
  input              rst_n         
  );

  wire wy36iirxspfw56864 = 1'b1;



  wire tx75ny_me9b15mo9 = ahbl_hready & bus_clk_en;


  wire xpoxafcifn9bt7d4;

  wire o0mpts6_n;
  wire bzrj54k7l7llo;
  wire y29zeznmb9;
  wire rcp39kxzwzrujoq;
  wire v77j9kx662fjy8;

  wire a1n_156c8l6j3t;
  wire lujkjdlze9ir0fkzi5j;
  wire w_cvn_004iq_92cu;
  wire rjb0ake6bkvi_uexrp;
  wire s5toprsofbaca65lg78g1;

  wire arl3n7ckluqs5vkij;































      assign xpoxafcifn9bt7d4  = 1'b0;
      assign o0mpts6_n   = 1'b0;
      assign bzrj54k7l7llo = 1'b0;
      assign y29zeznmb9 = 1'b0;
      assign rcp39kxzwzrujoq = 1'b0;
      assign v77j9kx662fjy8 = 1'b0;

      assign arl3n7ckluqs5vkij = 1'b0;

      assign a1n_156c8l6j3t   = 1'b0;
      assign lujkjdlze9ir0fkzi5j = 1'b0;
      assign w_cvn_004iq_92cu = 1'b0;
      assign rjb0ake6bkvi_uexrp = 1'b0;
      assign s5toprsofbaca65lg78g1 = 1'b0;










  wire v706iusq08t42dr9;
  wire r6sgqz3qozop_78f;


  wire bap6f5epfkrw1qc = tx75ny_me9b15mo9 & ahbl_htrans[1];

 wire bov6iggub5nn246qx = bap6f5epfkrw1qc;  
 wire rln9rwa2epujlx = bus_clk_en & (ahbl_htrans == 2'b0);
 wire ftuhlxrh0247tw = bov6iggub5nn246qx | rln9rwa2epujlx;
 wire ud5em0ounnh90859 = rln9rwa2epujlx ? 1'b0 : (~(ahbl_hburst == 3'b0));
 wire s1vlx4vpc6x9a7z;

 ux607_gnrl_dfflr #(1) nx2pkh44k874l468 (ftuhlxrh0247tw, ud5em0ounnh90859, s1vlx4vpc6x9a7z, clk, rst_n);






















  assign icb_cmd_ready  = tx75ny_me9b15mo9   & (~v706iusq08t42dr9);
  assign ahbl_htrans[1] = icb_cmd_valid & (~v706iusq08t42dr9);


  assign ahbl_htrans[0] = s1vlx4vpc6x9a7z ? icb_cmd_hseq : 1'b0;




  localparam qet2jodq6p  = 2;
  localparam vvgygupma0 = 2'b00; 
  localparam ay22jhu = 2'b01;
  localparam me7m0orwjhi = 2'b10;

  wire[qet2jodq6p-1:0] avzmm87w3kglnb5;
  wire[qet2jodq6p-1:0] it5ozza4tacg;

  wire z0rei8ewbehy = bap6f5epfkrw1qc & ahbl_hwrite;
  wire y8jt5vaziqir7j = bap6f5epfkrw1qc & (~ahbl_hwrite);
  wire i_sml2_3euhg2h = tx75ny_me9b15mo9 & (~ahbl_htrans[1]);

  wire  u49jscbid_zl7e = (avzmm87w3kglnb5 == vvgygupma0);


  assign it5ozza4tacg = tx75ny_me9b15mo9 ?  (
                               {qet2jodq6p{i_sml2_3euhg2h}} & (vvgygupma0) 
                             | {qet2jodq6p{z0rei8ewbehy}} & (ay22jhu)
                             | {qet2jodq6p{y8jt5vaziqir7j}} & (me7m0orwjhi)
                         ) : avzmm87w3kglnb5;


  ux607_gnrl_dffr #(qet2jodq6p) maqgcj2hln_86h (it5ozza4tacg, avzmm87w3kglnb5, clk, rst_n);

  wire [DW-1:0]fns8_auk6bx1mp;
  wire nazlbbvkmagsapws043 = z0rei8ewbehy;
  ux607_gnrl_dfflr #(DW) oewvhqfu6k29ioq2ji (nazlbbvkmagsapws043, icb_cmd_wdata, fns8_auk6bx1mp, clk, rst_n);




  assign ahbl_hwrite = ~icb_cmd_read;    
  assign ahbl_haddr  = icb_cmd_addr;    
  assign ahbl_hsize  = {1'b0,icb_cmd_size};    
  assign ahbl_hexcl  = icb_cmd_excl;    
  assign ahbl_hburst = icb_cmd_burst;
  assign ahbl_hwdata = fns8_auk6bx1mp;

  assign ahbl_hprot  = icb_cmd_hprot ;
  assign ahbl_hattri = icb_cmd_attri;


  wire qzk27vwr9nlli9n  = (~icb_cmd_dmode) & (~icb_cmd_hprot[0]);
  wire vffty9dks1z4369 = (~icb_cmd_dmode) & icb_cmd_hprot[0];
  wire hx1s4cyg43_yuo  = icb_cmd_dmode;

  wire [1:0] g9nt_7hlbzbpwfh6 = 
                        vffty9dks1z4369 ? 2'b00 :
                        hx1s4cyg43_yuo ? 2'b01 :
                        qzk27vwr9nlli9n ? 2'b10 :
                                      2'b11;
  assign ahbl_master = g9nt_7hlbzbpwfh6;

  assign icb_rsp_valid = ahbl_hready & (~u49jscbid_zl7e);  
  assign icb_rsp_rdata = ahbl_hrdata;   
  assign icb_rsp_err   = ahbl_hresp[0];
  assign icb_rsp_excl_ok   = ahbl_hresp_exok;


  wire uwy7_yj98jvt2txl8;
  wire jv36i_7i91oi6z0_1;
  wire j4m355hz01jwcc4z;
  wire m_mn82s6u2u75_yuh2;

  wire kj8wwsv34og24o;
  wire cjkp0r7a6b75zxi;
  wire fkwb0t7wf_xcl;
  wire btn06r3ay0ydt76s;






  generate

    if(SUPPORT_LOCK == 1) begin:dwylazwt1o
      assign ahbl_hlock    = ((icb_cmd_lock & icb_cmd_valid) | r6sgqz3qozop_78f) 
                           & (~v706iusq08t42dr9)  
                           & (~(
                                  ((~icb_cmd_lock) & icb_cmd_valid)
                               )
                             );



      assign uwy7_yj98jvt2txl8 = cjkp0r7a6b75zxi;

      assign jv36i_7i91oi6z0_1 = v706iusq08t42dr9 & i_sml2_3euhg2h;
      assign j4m355hz01jwcc4z = uwy7_yj98jvt2txl8 | jv36i_7i91oi6z0_1;
      assign m_mn82s6u2u75_yuh2 = uwy7_yj98jvt2txl8 & (~jv36i_7i91oi6z0_1);
      ux607_gnrl_dfflr #(1) kn2qnj_4g3axckorsu (j4m355hz01jwcc4z, m_mn82s6u2u75_yuh2, v706iusq08t42dr9, clk, rst_n);











      assign kj8wwsv34og24o = (bap6f5epfkrw1qc & icb_cmd_lock);




      assign cjkp0r7a6b75zxi = r6sgqz3qozop_78f & (
                             (bap6f5epfkrw1qc & (~icb_cmd_lock))

                           )
                           ;
      assign fkwb0t7wf_xcl = kj8wwsv34og24o | cjkp0r7a6b75zxi;
      assign btn06r3ay0ydt76s = kj8wwsv34og24o & (~cjkp0r7a6b75zxi);
      ux607_gnrl_dfflr #(1) arrc4fx9g7ji4ds (fkwb0t7wf_xcl, btn06r3ay0ydt76s, r6sgqz3qozop_78f, clk, rst_n);
    end

    else begin: ovaieqiabzlow61
      assign uwy7_yj98jvt2txl8 = 1'b0;
      assign jv36i_7i91oi6z0_1 = 1'b0;
      assign j4m355hz01jwcc4z = 1'b0;
      assign m_mn82s6u2u75_yuh2 = 1'b0;

      assign kj8wwsv34og24o = 1'b0;
      assign cjkp0r7a6b75zxi = 1'b0;
      assign fkwb0t7wf_xcl = 1'b0;
      assign btn06r3ay0ydt76s = 1'b0;


      assign ahbl_hlock    = 1'b0;
      assign v706iusq08t42dr9   = 1'b0;
      assign r6sgqz3qozop_78f   = 1'b0;
    end

  endgenerate




  assign icb2ahbl_pend_active = v706iusq08t42dr9 | s1vlx4vpc6x9a7z;

endmodule 










module ux607_gnrl_ahbl2icb
  #(
    parameter AW = 32,
    parameter DW = 32 
    )
  (

  output             ahbl2icb_active,



  input              ahbl_hsel,   
  input              ahbl_hexcl,   
  input  [1:0]       ahbl_htrans,   
  input              ahbl_hwrite,   
  input  [AW    -1:0]ahbl_haddr,    
  input  [2:0]       ahbl_hsize,    
  input  [DW    -1:0]ahbl_hwdata,
  input              ahbl_huser,



  output  [DW   -1:0]ahbl_hrdata,   
  output  [1:0]      ahbl_hresp,    
  output             ahbl_hresp_exok,    
  input              ahbl_hready_in,   
  output             ahbl_hready_out,   

  output             icb_cmd_sel, 

  output             icb_cmd_valid, 
  input              icb_cmd_ready, 
  output             icb_cmd_read, 
  output  [AW-1:0]   icb_cmd_addr,
  output             icb_cmd_user,
  output  [DW-1:0]   icb_cmd_wdata, 
  output  [(DW/8-1):0] icb_cmd_wmask,
  output  [1:0]      icb_cmd_size,
  output             icb_cmd_excl,   



  input              icb_rsp_valid, 
  output             icb_rsp_ready, 
  input              icb_rsp_err,
  input              icb_rsp_excl_ok,
  input  [DW-1:0]    icb_rsp_rdata, 

  input              clk,          
  input              rst_n         
  );



  wire  v9ov1b3vn5k4ctkb;
  wire  ub9pjiu4juf6nuqoq2w6;
  wire  ogvavqa7ta836s;
  wire  l089k6vccrfphrtw;
  wire  [AW-1:0] aw0a19a967dn7n0x25w; 
  wire  qc9p77b285nqot; 
  wire  [DW-1:0] sc169gxpr38lpe8; 
  wire  [(DW/8-1):0] hg1g2yh6yktfe_btdst7; 
  wire  [2-1:0] leieaos4fnc5s_81kr; 

  localparam hv5mlbfaebnkypctu = (AW+DW+(DW/8)+4+1);
  wire [hv5mlbfaebnkypctu-1:0] ez0jkdg20o7_ib;
  wire [hv5mlbfaebnkypctu-1:0] djfdd4cy1d_i5vg =  {
                      ogvavqa7ta836s, 
                      l089k6vccrfphrtw, 
                      aw0a19a967dn7n0x25w,
                      qc9p77b285nqot,
                      sc169gxpr38lpe8, 
                      hg1g2yh6yktfe_btdst7, 
                      leieaos4fnc5s_81kr  
                    };
  assign {
                      icb_cmd_read, 
                      icb_cmd_excl, 
                      icb_cmd_addr,
					  icb_cmd_user,
                      icb_cmd_wdata, 
                      icb_cmd_wmask, 
                      icb_cmd_size  
                    } = ez0jkdg20o7_ib;


  ux607_gnrl_bypbuf # (
   .DP(1),
   .DW(hv5mlbfaebnkypctu)
  ) lquetohr9xd39fj_d(
    .i_vld(v9ov1b3vn5k4ctkb), 
    .i_rdy(ub9pjiu4juf6nuqoq2w6), 
    .i_dat(djfdd4cy1d_i5vg),
    .o_vld(icb_cmd_valid), 
    .o_rdy(icb_cmd_ready), 
    .o_dat(ez0jkdg20o7_ib),

    .clk  (clk  ),
    .rst_n(rst_n)  
   );




  wire dy9ll1o6t6ytby71hf4;
  wire ow4hbh48f0mt6le4o;
  wire uzwj715coelxmfqs;
  wire sihcnyg6z96riwnnw_np;
  wire [DW-1:0] dek0xt7q6guk2vf6; 

  wire [DW+2-1:0]ziubvvomv2nddezv;
  wire [DW+2-1:0]kgh1znd6ahvjhj;

  assign kgh1znd6ahvjhj = {
                          icb_rsp_excl_ok,
                          icb_rsp_err,
                          icb_rsp_rdata
                          };

  assign {
                          sihcnyg6z96riwnnw_np,
                          uzwj715coelxmfqs,
                          dek0xt7q6guk2vf6
                          } = ziubvvomv2nddezv;

  ux607_gnrl_bypbuf # (
    .DP(1),
    .DW(DW+2) 
  ) oakf7pdt8qf2ffmokrq8s0a(
      .i_vld   (icb_rsp_valid),
      .i_rdy   (icb_rsp_ready),

      .o_vld   (dy9ll1o6t6ytby71hf4),
      .o_rdy   (ow4hbh48f0mt6le4o),

      .i_dat   (kgh1znd6ahvjhj),
      .o_dat   (ziubvvomv2nddezv),

      .clk     (clk  ),
      .rst_n   (rst_n)
  );


  wire k22p5hfn4flvvrsx = ahbl_hready_out & ahbl_hready_in;

  wire vho3hf4e5c_jie2e5num  =

        ahbl_hsel

      & ahbl_htrans[1] 
      ;

  wire tk6k_fy7j7yzlulnx  = vho3hf4e5c_jie2e5num

      & k22p5hfn4flvvrsx;

  wire [1:0] ysp4qylgpi14tq5ei;

  wire gskbfu9e5zjcbwxum  = 

        ysp4qylgpi14tq5ei[1] 

      & k22p5hfn4flvvrsx;

  wire a2cfz2uuae81g;
  wire wfldzwh25ntc3ageaue = k22p5hfn4flvvrsx;
  wire f9pxtpa_6gspdp8xz0q8 = tk6k_fy7j7yzlulnx;
  ux607_gnrl_dfflr #(1) n1psx12qleb9ys88b_as (wfldzwh25ntc3ageaue, f9pxtpa_6gspdp8xz0q8, a2cfz2uuae81g, clk, rst_n);






  wire jx0jqq_arfubsf7 = k22p5hfn4flvvrsx;
  wire [1:0] j30cmax5pajkly7 = ahbl_htrans;
  ux607_gnrl_dfflr #(2) ocm6bg3vsj4il4wlfs (jx0jqq_arfubsf7, j30cmax5pajkly7, ysp4qylgpi14tq5ei, clk, rst_n);

  wire fl2hafaygmmow65h;
  wire i60nitrgupy7qze = k22p5hfn4flvvrsx;
  wire owu8qejj04lh6evkn5a = ahbl_hexcl;
  ux607_gnrl_dfflr #(1) sw3ya5n7uxb5xtgcqi60g (i60nitrgupy7qze, owu8qejj04lh6evkn5a, fl2hafaygmmow65h, clk, rst_n);

  wire [1:0] r2po5xb39zit;
  wire xcwx9l0wizjfmim = k22p5hfn4flvvrsx;
  wire [1:0] gj5bkqu_442yx1n40yu = ahbl_hsize[1:0];
  ux607_gnrl_dfflr #(2) uojogcss2zfo5lx2g (xcwx9l0wizjfmim, gj5bkqu_442yx1n40yu, r2po5xb39zit, clk, rst_n);

  wire xtqy0z3x6f47a5xlk2 = k22p5hfn4flvvrsx;
  wire [AW-1:0] w490nquvx0gj_;
  wire [AW-1:0] fbtq6gbc7jmb29i9ul = ahbl_haddr;
  ux607_gnrl_dfflr #(AW) spc3le_lqt1vat6f48c15 (xtqy0z3x6f47a5xlk2, fbtq6gbc7jmb29i9ul, w490nquvx0gj_, clk, rst_n);

  wire z8pbhqxqlco954rhg = k22p5hfn4flvvrsx;
  wire wm4ctwhlq7abl9vb;
  wire wrxky4n1bsmcm1p = ahbl_huser;
  ux607_gnrl_dfflr #(1) pyrp6o9g1d8x3_5vw (z8pbhqxqlco954rhg, wrxky4n1bsmcm1p, wm4ctwhlq7abl9vb, clk, rst_n);


  wire sbfb89ar9g4e;

  assign ogvavqa7ta836s = sbfb89ar9g4e ? 1'b0 : 1'b1;  
  assign aw0a19a967dn7n0x25w = sbfb89ar9g4e ? w490nquvx0gj_ : ahbl_haddr;
  assign qc9p77b285nqot = sbfb89ar9g4e ? wm4ctwhlq7abl9vb : ahbl_huser;
  assign leieaos4fnc5s_81kr = sbfb89ar9g4e ? r2po5xb39zit[1:0] : ahbl_hsize[1:0];
  assign l089k6vccrfphrtw = sbfb89ar9g4e ? fl2hafaygmmow65h : ahbl_hexcl;
  assign sc169gxpr38lpe8 = ahbl_hwdata; 


  wire [(DW/8-1):0] xh1ov17gxap8xp967;
  wire [(DW/8-1):0] gykofhynkgdwyada3h5;

  wire ovbw2ge12bcjlsrib3t1 = k22p5hfn4flvvrsx;
  wire [(DW/8-1):0] ww1q8kqrai87lkg9mq = xh1ov17gxap8xp967;
  ux607_gnrl_dfflr #(DW/8) wlj5hmz9l32pn_j7gxm6gw (ovbw2ge12bcjlsrib3t1, ww1q8kqrai87lkg9mq, gykofhynkgdwyada3h5, clk, rst_n);

  assign hg1g2yh6yktfe_btdst7 = gykofhynkgdwyada3h5; 

  generate 

  if(DW == 64) begin:bh9h6t0g5q_n
     assign xh1ov17gxap8xp967 = 
         (ahbl_hsize == 3'b000) ? (4'b1 << ahbl_haddr[2:0])
       : (ahbl_hsize == 3'b001) ? (4'b11 << {ahbl_haddr[2:1],1'b0})
       : (ahbl_hsize == 3'b010) ? (4'b1111 << {ahbl_haddr[2],2'b0})

       : (8'b1111_1111)
       ;
  end

  if(DW == 32) begin:r_5ssyvcqw9
     assign xh1ov17gxap8xp967 = 
         (ahbl_hsize == 3'b000) ? (4'b1 << ahbl_haddr[1:0])
       : (ahbl_hsize == 3'b001) ? (4'b11 << {ahbl_haddr[1:1],1'b0})

       : (ahbl_hsize == 3'b010) ? (4'b1111)

       : (4'b1111)
       ;
  end

  endgenerate

  wire m38dev21ov3pe8jjqun4;
  wire yzg5met0xqgc6lduitq3n;
  wire d0qh365dtr6viqwzpncyg0ct = dy9ll1o6t6ytby71hf4 & yzg5met0xqgc6lduitq3n;
  wire ry__6funfjr6nf6w5dun = m38dev21ov3pe8jjqun4 & k22p5hfn4flvvrsx;
  wire wolj0jptzljq4g03n1l9q = d0qh365dtr6viqwzpncyg0ct | ry__6funfjr6nf6w5dun; 
  wire rhrkou30g8ou2w3ylm3_x42q4 = d0qh365dtr6viqwzpncyg0ct | (~ry__6funfjr6nf6w5dun); 
  ux607_gnrl_dfflr #(1) nntmqm7mh256au_noe9iq27qp (wolj0jptzljq4g03n1l9q, rhrkou30g8ou2w3ylm3_x42q4, m38dev21ov3pe8jjqun4, clk, rst_n);

  wire l5_854x2xqxvorikov = (vho3hf4e5c_jie2e5num & ahbl_hwrite);

  wire smgh49vlhb87z6ewet = wfldzwh25ntc3ageaue & l5_854x2xqxvorikov;
  wire z6on__qyneteip28 = v9ov1b3vn5k4ctkb & ub9pjiu4juf6nuqoq2w6 & (~ogvavqa7ta836s);
  wire zkhfflrkgf_rlcopt5o = smgh49vlhb87z6ewet | z6on__qyneteip28; 
  wire es0s1yfvc84zifhrs_ = smgh49vlhb87z6ewet | (~z6on__qyneteip28); 
  ux607_gnrl_dfflr #(1) qzegzxdk67g30hxu0g (zkhfflrkgf_rlcopt5o, es0s1yfvc84zifhrs_, sbfb89ar9g4e, clk, rst_n);

  wire cjaplq_da70txumt;
  wire h2rmo3o27yvs5bcfsu = v9ov1b3vn5k4ctkb & ub9pjiu4juf6nuqoq2w6 & ogvavqa7ta836s;
  wire iujuu3i8nradk6qrv0s = dy9ll1o6t6ytby71hf4 & ow4hbh48f0mt6le4o & cjaplq_da70txumt;
  wire z87owt3w5r7vjueu = h2rmo3o27yvs5bcfsu | iujuu3i8nradk6qrv0s; 
  wire askhpywchgt7f5mca = h2rmo3o27yvs5bcfsu | (~iujuu3i8nradk6qrv0s); 
  ux607_gnrl_dfflr #(1) vbgb0hmg7xqagzgu7d0y1 (z87owt3w5r7vjueu, askhpywchgt7f5mca, cjaplq_da70txumt, clk, rst_n);

  wire a1n_156c8l6j3t;
  wire kouhyfs99s2xt8qfr = v9ov1b3vn5k4ctkb & ub9pjiu4juf6nuqoq2w6;
  wire yk4t8yu2epj8 = dy9ll1o6t6ytby71hf4 & ow4hbh48f0mt6le4o;
  wire r8axmur45uwwts_z = kouhyfs99s2xt8qfr ^ yk4t8yu2epj8;
  wire [2-1:0] ta6v7ss882s4;
  wire [2-1:0] w71i8osb89s79fy = kouhyfs99s2xt8qfr ? (ta6v7ss882s4 + 1'b1) : (ta6v7ss882s4 - 1'b1);
  ux607_gnrl_dfflr #(2) hh67nplqgwfr382l5y7 (r8axmur45uwwts_z, w71i8osb89s79fy, ta6v7ss882s4, clk, rst_n);

  assign a1n_156c8l6j3t = (~(ta6v7ss882s4 == {2{1'b0}}));


  wire gbjm5za8l9etp;
  wire u7d126psw95_0fj = kouhyfs99s2xt8qfr;
  wire c1pxt2sk9rzorz63_6 = ogvavqa7ta836s;
  ux607_gnrl_dfflr #(1) fsdkrikspmvveulc06ooi (u7d126psw95_0fj, c1pxt2sk9rzorz63_6, gbjm5za8l9etp, clk, rst_n);

  wire t20grifz_pud7_1cmugvs = (vho3hf4e5c_jie2e5num & (~ahbl_hwrite));
  wire btw1d72vb49b1v4wv;
  assign v9ov1b3vn5k4ctkb = (
                 (t20grifz_pud7_1cmugvs & btw1d72vb49b1v4wv)
               | sbfb89ar9g4e) 
               ;

  assign icb_cmd_sel = vho3hf4e5c_jie2e5num | sbfb89ar9g4e | a1n_156c8l6j3t; 

  assign yzg5met0xqgc6lduitq3n = (uzwj715coelxmfqs & gbjm5za8l9etp) ? (~m38dev21ov3pe8jjqun4) : 1'b0;

  wire   gcngsz_zjod7bh = (a1n_156c8l6j3t & (~gbjm5za8l9etp)); 

  assign btw1d72vb49b1v4wv = 
                (a1n_156c8l6j3t ? ((ta6v7ss882s4 == 2'b1) & dy9ll1o6t6ytby71hf4) : 1'b1) & 
                ((gcngsz_zjod7bh & (~ahbl_hwrite)) ? dy9ll1o6t6ytby71hf4 : 1'b1) & 
                ((gcngsz_zjod7bh & ahbl_hwrite & ahbl_hexcl) ? dy9ll1o6t6ytby71hf4 : 1'b1) & 
                (

                  (~a2cfz2uuae81g) ? 1'b1 : 

                  cjaplq_da70txumt ? (~yzg5met0xqgc6lduitq3n) : 


                  sbfb89ar9g4e ? (ahbl_hwrite & (~ahbl_hexcl)) : 
                  1'b1);
  assign ahbl_hready_out = ub9pjiu4juf6nuqoq2w6 & btw1d72vb49b1v4wv; 

  assign ow4hbh48f0mt6le4o = (ahbl_hready_in & (~yzg5met0xqgc6lduitq3n)) 

                         | gcngsz_zjod7bh;

  assign ahbl_hrdata = dek0xt7q6guk2vf6;


  assign ahbl_hresp[0]  = 1'b0;
  assign ahbl_hresp[1]  = 1'b0;
  assign ahbl_hresp_exok  = sihcnyg6z96riwnnw_np;

  assign ahbl2icb_active = v9ov1b3vn5k4ctkb | icb_cmd_valid | a1n_156c8l6j3t | ahbl_htrans[1];

endmodule 











module ux607_gnrl_icb_active # (

  parameter OUTS_CNT_W = 1
) (

  output             icb_active,

  input              icb_cmd_valid, 
  input              icb_cmd_ready, 

  input              icb_rsp_valid, 
  input              icb_rsp_ready, 

  input              clk,          
  input              rst_n         
  );


  wire kouhyfs99s2xt8qfr = icb_cmd_valid & icb_cmd_ready;
  wire yk4t8yu2epj8 = icb_rsp_valid & icb_rsp_ready;

  wire r8axmur45uwwts_z = kouhyfs99s2xt8qfr ^ yk4t8yu2epj8;

  wire [OUTS_CNT_W-1:0] ta6v7ss882s4;
  wire [OUTS_CNT_W-1:0] w71i8osb89s79fy = kouhyfs99s2xt8qfr ? (ta6v7ss882s4 + 1'b1) : (ta6v7ss882s4 - 1'b1);
  ux607_gnrl_dfflr #(OUTS_CNT_W) hh67nplqgwfr382l5y7 (r8axmur45uwwts_z, w71i8osb89s79fy, ta6v7ss882s4, clk, rst_n);

  assign icb_active = icb_cmd_valid | (~(ta6v7ss882s4 == {OUTS_CNT_W{1'b0}}));


endmodule 












module ux607_gnrl_icb2apb # (
  parameter CUT_READY = 1,
  parameter AW = 32,
  parameter DW = 32 
) (
  input              icb_cmd_valid, 
  output             icb_cmd_ready, 
  input              icb_cmd_read, 
  input  [AW-1:0]    icb_cmd_addr, 
  input  [DW-1:0]    icb_cmd_wdata, 
  input  [(DW/8-1):0]  icb_cmd_wmask,
  input  [1:0]       icb_cmd_size,
  input              icb_cmd_dmode,
  input              icb_cmd_mmode,
  input              icb_cmd_smode,

  output             icb_rsp_valid, 
  input              icb_rsp_ready, 
  output             icb_rsp_err,
  output [DW-1:0]    icb_rsp_rdata, 
  
  output [AW-1:0] apb_paddr,
  output          apb_pwrite,
  output          apb_psel,
  output          apb_dmode,
  output [2:0]    apb_pprot,
  output [3:0]    apb_pstrobe,
  output          apb_penable,
  output [DW-1:0] apb_pwdata,
  input  [DW-1:0] apb_prdata,
  input           apb_pready,
  input           apb_pslverr,

  input  clk,  
  input  rst_n
  );


  
  
  
  
  
  
  wire e3k3c6jyr1wjx;

  wire v9ov1b3vn5k4ctkb;
  wire ub9pjiu4juf6nuqoq2w6;
  wire dy9ll1o6t6ytby71hf4;
  wire ow4hbh48f0mt6le4o;
  wire uzwj715coelxmfqs;
  wire sihcnyg6z96riwnnw_np;
  wire [DW-1:0] dek0xt7q6guk2vf6; 
  wire [DW+1-1:0]ziubvvomv2nddezv;


  wire bx5dmny2mt_9zz3an8f;
  wire p203154jjq0bymz90k3t;
  
  wire [DW+1-1:0] xw4ju3m2k6rsjtoipo;

  wire [DW+1-1:0] kgh1znd6ahvjhj;

  wire a1n_156c8l6j3t;
  wire lujkjdlze9ir0fkzi5j = icb_cmd_valid & icb_cmd_ready;
  wire w_cvn_004iq_92cu = bx5dmny2mt_9zz3an8f & p203154jjq0bymz90k3t;
  wire rjb0ake6bkvi_uexrp = lujkjdlze9ir0fkzi5j | w_cvn_004iq_92cu; 
  wire s5toprsofbaca65lg78g1 = lujkjdlze9ir0fkzi5j | (~w_cvn_004iq_92cu); 
  ux607_gnrl_dfflr #(1) j9j9tnqhq8oep38tws6n(rjb0ake6bkvi_uexrp, s5toprsofbaca65lg78g1, a1n_156c8l6j3t, clk, rst_n);

  
  wire kbje5ox2409b4x4 =  (~a1n_156c8l6j3t) | w_cvn_004iq_92cu;

  assign v9ov1b3vn5k4ctkb = kbje5ox2409b4x4 & icb_cmd_valid;
  assign icb_cmd_ready   = kbje5ox2409b4x4 & ub9pjiu4juf6nuqoq2w6;


  assign ziubvvomv2nddezv = {
                          uzwj715coelxmfqs,
                          dek0xt7q6guk2vf6
                          };

  assign {
                          icb_rsp_err,
                          icb_rsp_rdata
                          } = kgh1znd6ahvjhj;


  ux607_gnrl_bypbuf # (
    .DP(1),
    .DW(DW+1) 
  ) o16j4hr_n43azd_dlwb6y71(
      .i_vld   (dy9ll1o6t6ytby71hf4),
      .i_rdy   (ow4hbh48f0mt6le4o),

      .o_vld   (bx5dmny2mt_9zz3an8f),
      .o_rdy   (p203154jjq0bymz90k3t),

      .i_dat   (ziubvvomv2nddezv),
      .o_dat   (xw4ju3m2k6rsjtoipo),
  
      .clk     (clk  ),
      .rst_n   (rst_n)
  );

  generate

  if(CUT_READY==1) begin:sktrpd6lnp4mrgz

  ux607_gnrl_bypbuf # (
    .DP(1),
    .DW(DW+1) 
  ) ydvjiz1qsgdhh8lnj6sdc6me(
      .i_vld   (bx5dmny2mt_9zz3an8f),
      .i_rdy   (p203154jjq0bymz90k3t),

      .o_vld   (icb_rsp_valid),
      .o_rdy   (icb_rsp_ready),

      .i_dat   (xw4ju3m2k6rsjtoipo),
      .o_dat   (kgh1znd6ahvjhj),
  
      .clk     (clk  ),
      .rst_n   (rst_n)
  );
  end
  else begin:euls1i3brh416bq
    assign kgh1znd6ahvjhj = xw4ju3m2k6rsjtoipo;
    assign icb_rsp_valid = bx5dmny2mt_9zz3an8f;
    assign p203154jjq0bymz90k3t = icb_rsp_ready;
  end

  endgenerate
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  assign dy9ll1o6t6ytby71hf4 = ub9pjiu4juf6nuqoq2w6;
  assign dek0xt7q6guk2vf6 = apb_prdata;

  assign uzwj715coelxmfqs = apb_pslverr;

    
         
         
  
  
  wire vkfariivah1kji = (~e3k3c6jyr1wjx) & icb_cmd_valid;
  assign ub9pjiu4juf6nuqoq2w6 = (e3k3c6jyr1wjx & apb_pready);
    
  wire xwrv9k91pl5yps3l = ub9pjiu4juf6nuqoq2w6;
  wire tx7u7gk_9k8c886r1 = vkfariivah1kji | xwrv9k91pl5yps3l;
  wire xk84via5umyd392 = vkfariivah1kji & (~xwrv9k91pl5yps3l);
  ux607_gnrl_dfflr #(1) t6y3u6tg2i4dd51kga8 (tx7u7gk_9k8c886r1, xk84via5umyd392, e3k3c6jyr1wjx, clk, rst_n);


  assign apb_paddr  = icb_cmd_addr;
  assign apb_pwrite = (~icb_cmd_read);
  assign apb_dmode  = icb_cmd_dmode;

  assign apb_pprot[0] = icb_cmd_mmode | icb_cmd_smode;
  assign apb_pprot[1] = 1'b1         ;
  assign apb_pprot[2] = 1'b0         ;

  assign apb_psel    = icb_cmd_valid;
  assign apb_penable = e3k3c6jyr1wjx;
  assign apb_pwdata  = icb_cmd_wdata;
  assign apb_pstrobe = icb_cmd_read ? {DW/8{1'b0}} : icb_cmd_wmask;

endmodule










module ux607_gnrl_apb2icb # (
  parameter AW = 32,
  parameter DW = 64 
) (
  output              icb_cmd_valid, 
  input               icb_cmd_ready, 
  output              icb_cmd_read, 
  output  [AW-1:0]    icb_cmd_addr, 
  output  [DW-1:0]    icb_cmd_wdata, 
  output  [(DW/8-1):0]  icb_cmd_wmask,
  output  [1:0]       icb_cmd_size,

  input               icb_rsp_valid, 
  
  input               icb_rsp_err,
  input   [DW-1:0]    icb_rsp_rdata, 
  
  input   [AW-1:0] apb_paddr,
  input            apb_pwrite,
  input            apb_psel ,
  input            apb_penable,
  input   [DW-1:0] apb_pwdata,
  output  [DW-1:0] apb_prdata,
  output           apb_pready,
  output           apb_pslverr,

  input  clk,  
  input  rst_n
  );

  assign apb_prdata  = icb_rsp_rdata;
  assign apb_pslverr = icb_rsp_err;

  assign apb_pready    = icb_cmd_ready;
  assign icb_cmd_valid = apb_psel & apb_penable;

  assign icb_cmd_read  = ~apb_pwrite;
  assign icb_cmd_addr  = apb_paddr;
  assign icb_cmd_wdata = apb_pwdata;
  assign icb_cmd_wmask = {DW/8{1'b1}};

  generate 
    if(DW == 8) begin:mapaysj
      assign icb_cmd_size = 2'b00;
    end
    if(DW == 16) begin:ryf5iemp_la8
      assign icb_cmd_size = 2'b01;
    end
    if(DW == 32) begin:kmwu2hcx3znc
      assign icb_cmd_size = 2'b10;
    end
    if(DW == 64) begin:qa954o41la5
      assign icb_cmd_size = 2'b11;
    end
  endgenerate

endmodule



















































































































































































































































































module ux607_gnrl_rbin4 # (
    parameter ARBT_NUM = 4
)(
  output[ARBT_NUM-1:0] grt_vec,  
  input [ARBT_NUM-1:0] req_vec,  
  input arbt_ena,   
  input clk,        
  input rst_n
);

  wire [ARBT_NUM-1:0] an03ge2t2lnqokt;
  wire [ARBT_NUM-1:0] c0_fjr1ekbr;

  genvar i;

  generate
      for(i = 0; i < ARBT_NUM; i = i+1)
      begin:shr0zu2xtqr9_iq9psn

        if(i==0) begin: xvpcp9wjmb99kn

          assign grt_vec[i] =  ~an03ge2t2lnqokt[0];
        end
        else if(i==(ARBT_NUM-1)) begin: w57_9w73hrvp6nndf

          assign grt_vec[i] =  (~(|req_vec[i-1:0])) | an03ge2t2lnqokt[0];
        end
        else begin:ccs98kfg22q4r73kas1les21q6a
          assign grt_vec[i] =  (~(|req_vec[i-1:0])) & (~an03ge2t2lnqokt[i]);
        end

      end
  endgenerate

  localparam a65wkc = 2;
  localparam p5qxocb = 3;
  wire [a65wkc-1:0] pb_3hk9ea0;

  wire ajgbfq66r4 = req_vec[ARBT_NUM-1] & (~grt_vec[ARBT_NUM-1]) & arbt_ena;

  wire yh750xgqgxwx =  req_vec[ARBT_NUM-1] & grt_vec[ARBT_NUM-1] & arbt_ena; 
  wire kv09wlfd =  yh750xgqgxwx & (|pb_3hk9ea0);
  wire v3vd66_q9 = ajgbfq66r4 | kv09wlfd;
  wire [a65wkc-1:0] ov6927s7pq8 = ajgbfq66r4 ? (pb_3hk9ea0 + 1'b1) : {a65wkc{1'b0}};
  ux607_gnrl_dfflr #(a65wkc) bwli31sfcrd (v3vd66_q9, ov6927s7pq8, pb_3hk9ea0, clk, rst_n);

  wire qvgk14nlz = (pb_3hk9ea0 == p5qxocb[a65wkc-1:0]);


  wire d8_oitpk = qvgk14nlz & ajgbfq66r4;

  wire iq56_qt5shnc4 = (|c0_fjr1ekbr) & yh750xgqgxwx;
  wire pjd96vtarupx = d8_oitpk | iq56_qt5shnc4;

  wire [ARBT_NUM-1:0] fyawtijy0_mr = d8_oitpk ? {1'b0,{ARBT_NUM-1{1'b1}}} : {ARBT_NUM{1'b0}};
  ux607_gnrl_dfflr #(ARBT_NUM) vazepyge_wr (pjd96vtarupx, fyawtijy0_mr, c0_fjr1ekbr, clk, rst_n);

  assign an03ge2t2lnqokt = c0_fjr1ekbr;

endmodule







































module as9e9kibsg2lccbbj9 #(
    parameter onr7l = 32
)(
    input [onr7l-1:0] ta7wib,
    input [onr7l-1:0] g35wi_,
    input [onr7l-1:0] h_kg5l,
    output ig1wj,

    input gf33atgy,
    input ru_wi
);

wire [onr7l:0] frgfco = {ta7wib[onr7l-1], ta7wib};
wire [onr7l:0] ii = {g35wi_[onr7l-1], g35wi_};
wire [onr7l:0] fij51v = ~{h_kg5l[onr7l-1],h_kg5l};

wire [onr7l:0] s = (frgfco ^ ii) ^ fij51v;

wire [onr7l:0] oz7_y5 = (frgfco & ii) | (frgfco & fij51v) | (ii & fij51v);

wire [onr7l:0] c = {oz7_y5[onr7l-1:0], 1'b0};

assign ig1wj = ((c ^ s) == {(onr7l+1){1'b1}});

endmodule




















module gdyqy_u6w0mpgo (
  input  pp7hxkc1fr9z2qqw,
  input  i_x3a8jgmo8qd81tcr,

  input  nvyp85muxi8p9u1y8brs,

  input  f48_2zc1qro_3dodmk8,
  input  vaiscz5bqo4k6ql0519,
  input  w93is2iaq5aikcpaqxg3,
  input  uuuoq6te8sq6lj_e02iqoc,
  output azqy5qfm4kwm7vkwu6e,
  output ig7796duzb8wqodp,

  input  qmd94avv02av64cbwaj42,
  output hv9e7_hu5oyc6e87832pmb,
  input  m4ndmqnlr5eisc8m2k6fd,
  input  [27-1:0] jcczlhzxqzl5dx51l,
  input  nkdn__tk5pvp4nczp7xysy5,
  input  [16-1:0] fhzpp1p52pmfd3syoo,
 
  output j8cjhcuf0m6xjvemdaz,
  output umc_2tn6um_9xaiy7_ksg0w,
  output uiyh4da4134sjv7gnmc,
  output q7ru87fmzxczveihcxcwh,
  input  s_eowfyzlvx7gjv542upo,
 
  output d40pep591l63yhmefp7i,

  output t57d026x085pay,
  input  k5th293qdrtsytaehbsk,
  output g6gwjq519o1w1m3csgrrf3,
  output [27-1:0] lo_2ny7_v71by78q3,
  output hbdj3fcr8qkfkgzq58o1o2ozh,
  output [16-1:0] m_k_n75bb0f_im9fu_,

  
  
  
  input                                    jgm2b78on4di5vswgsdt,           
  input  [74-1:0]       tuui0ewt7j2chov1tdfd,          
  output                                   u_g5yts7tlcxo7ykedbqiv4ji0,         
  output                                   qdiqiuzopx36bi3s6fbh7mc16h2cj0,     
  output [5:0]                             urdbh4qug0s4u_dxqek3ejkxxgejj,      

  
  
  
  input  dep51yq,
  
  output                                   wk9s3wmc2q0yaa13,                
  output  [27-1:0]     s7re1eyp36bjvie,                 
  output  [1:0]                            a1pnq3ko2aaldi7h3xwme,          
  
  input                                    oq4nxgat71_rnebbasjmv9,          
  input                                    rj1ewmv16hujp9xlnpm6a3hhu9y8ml,     
  input                                    ryfblq1f8us1a8u3gy2gijl12x085ja,   
  input  [51-1:0]       j6q7tn13h_mjup45od1mu,           
  input                                    x81uu_gb6esoi095hudjgylqn,         
  input                                    ql2if76ihe_ppb4rp3buw7,         



  input  th06du2c8e2_b7k, 
  output irjoi8wvo25u209f_5,
  input  [64-1:0] zvk11dhgg2s67mkq, 
  input  r8nzx6_1no31zeloft,
  input  fbzs0o4ysyuzeg_qdj,
  input  me1n4pvwxa7n3u8l05,
  input  qaidts35dk5jcji0n, 

  output phzkntckzzbndu4wevf1o6, 
  output bpyef3a0dnkkyqdpymy, 
  output wv442dsr_nxty0qoldk7qmqg, 
  output b2loifdzo9b2smec06r0t, 
  output tx07brh7_ullbwlubonaqwg2,   
  output [64-1:0] ba1ucnyekcm68i9wuqwmn, 


  output                           ldqpjrsj9dp8yg3uc,  
  output                           s70e4xdis3p67ndpn6fbx,  
  output [7-1:0] h9zlka3j3ih8ihpvwvky1, 
  
  output [54-1:0] tf_tmpul8i8qbm_djvtl5f,          
  input  [54-1:0] qtsqtuxyont41a7h7i6,

  output                           w0ve66vjdz8lzwws3ic,  
  output                           df775k2ts6dn4528iq_ce5,  
  output [9-1:0] k3dychuj1pv4vw7cfj01ft8v, 
  
  output [64-1:0] jh4zf96qrsb31j072n,          
  input  [64-1:0] vfvtxk4jkkc3ql7_rqd,

  output                           hv6xxz3oswj4wy4j46,  
  output                           q6p7kcdd9o7j3e2c886,  
  output [7-1:0] ee_yaeclihal4dht69liwy6z, 
  
  output [54-1:0] thl4cxcuzntax8hnsn9bl4,          
  input  [54-1:0] mysqpp41yovfcis6f2dza47,

  
  output                           vp3x08mx4e27x4k26n,  
  output                           a7b829uahvy2i28yzgg,  
  output [9-1:0] kzxrmeg90fb06oya08h1, 
  
  output [64-1:0] kl5wycr14v5ukl7oqfhwe6,          
  input  [64-1:0] wt6c82_zmqgmt7if41t698,



  output  rinamilgle00i5xmx_vt, 
  input   j8wlfupbw25hdmohz5q0,
  output  [64-1:0] z64bwdr23steb7s9y9j, 
  output  bg1spy6_v2kbo75pz1d6,
  output  [2:0] b7aet1zp_fcfxn8h7rw0u1,
  output  [1:0] t3szwnvfo2nj3wk6r5kvt,
  output  cneu8a119tg3vmie6zr2h_,
  output  jw2dzv9gi7gygudyqql6fz,
  output  ybcilssdlw64sqj1jf2uuk,
  output  o_7kpry6inkqpqi1bf1nd,
  output  znotwr53pu47f5m1agm   ,
  output [1:0] bngbyv57e7juc0vkk2y8i   ,

  input   ze2bfnigu62i9937pcxnjc, 
  input   dm5b92mx0redfbuhs1u3d, 
  input   [64-1:0] c3vtv1izxu7rm5646jsmmke,

  input [8*32-1:0] pcr4upio7_tx37, 
  input [8*1-1:0] uzklqlncpqqm1rav,
  input [8*1-1:0] ortueunvnkx_l5m_j,
  input [8*1-1:0] hwuhtb7ucto_utk56,
  input [8*2-1:0] i1env2kmns7qvvuuc,
  input [8*1-1:0] g3s3vpafvy3i,


  input  c4ughu0qm5sfai,
  input  gc4b3kdcan6do88ta_,

  output wz_if_2q_23jhl2,
  input  gf33atgy,
  input  ru_wi
  );

  localparam wq7_4t7xmr99 = 2;


  wire tlmb65lrny6own    = jgm2b78on4di5vswgsdt;
  wire qqz76r4390y_pzoug  = tuui0ewt7j2chov1tdfd[5];
  wire r96xqbs4rp4ud91vy  = tuui0ewt7j2chov1tdfd[6];
  wire ha3mzwrvohf1v4m9  = tuui0ewt7j2chov1tdfd[7];
  wire c4197epxq1j27j_    = tuui0ewt7j2chov1tdfd[1] & ~tuui0ewt7j2chov1tdfd[0];
  wire vkt5l8auhc9hkqf   = tuui0ewt7j2chov1tdfd[2];
  wire h8yhw0bhacd77xw = tuui0ewt7j2chov1tdfd[3];
  wire wzrv89a8lbkafx2qdx = tuui0ewt7j2chov1tdfd[0];
  wire [64-1:0] nkj14m5ilghbj = tuui0ewt7j2chov1tdfd[74-1:10];  

  wire zla7uqbb3yfvop1ja9 = c4ughu0qm5sfai;
  wire fnjtncb80f_1t9v1mn5;
  wire gf3aiywpsjayl9nw6y_rl_r;
  wire hsv3kgrb3c_k_9x6hb;
  wire syeryna6edz5he27_zgkify;
  
  ux607_gnrl_dffr #(1) k1twmto5d66302213o849gk (zla7uqbb3yfvop1ja9    , fnjtncb80f_1t9v1mn5, gf33atgy, ru_wi);
  ux607_gnrl_dffr #(1) kex7m81u0yuh1l9_kxujrpg3oh (fnjtncb80f_1t9v1mn5, gf3aiywpsjayl9nw6y_rl_r, gf33atgy, ru_wi);
  ux607_gnrl_dffr #(1) sy5z2392vbppdpknt27b1m6oph (gf3aiywpsjayl9nw6y_rl_r, hsv3kgrb3c_k_9x6hb, gf33atgy, ru_wi);
  ux607_gnrl_dffr #(1) uqzb7645ng6kxy8kb_a0knchg (hsv3kgrb3c_k_9x6hb, syeryna6edz5he27_zgkify, gf33atgy, ru_wi);
 
  wire raha4wzwsh_g_zg = (~nvyp85muxi8p9u1y8brs) & syeryna6edz5he27_zgkify;
  
  wire nywm0kv90g64r5310wz = 
                 fnjtncb80f_1t9v1mn5 
               | gf3aiywpsjayl9nw6y_rl_r 
               | hsv3kgrb3c_k_9x6hb 
               | syeryna6edz5he27_zgkify ;

  wire jlihkmvsqt_p1_x;
  wire e4exh90ggokeh;
  wire uz8uoctou96a_0m95zx = 
                 zla7uqbb3yfvop1ja9 
               | nywm0kv90g64r5310wz
               | e4exh90ggokeh;
  
  wire vyneby1uawco;
  wire lh8ggdb3m21qvo0q;
  wire lm7s5990gmfb;
  
  
  wire n8hk7_wggv11dp5_wcn7kn;
  wire fb2yieg4ys3p19gmk96ooyq66 =   n8hk7_wggv11dp5_wcn7kn
                               | (lh8ggdb3m21qvo0q)
                               ;

  
  
  
  
  
  
  
  
  
  wire gysg24e47c3aqwd9wkc7m;
  wire ce4pb74pw07ylxuf649mb4j = f48_2zc1qro_3dodmk8 & ~gysg24e47c3aqwd9wkc7m;
  ux607_gnrl_dffr #(1) e1qlnzm32b2h97m_4y2xywur (f48_2zc1qro_3dodmk8, gysg24e47c3aqwd9wkc7m, gf33atgy, ru_wi);

  
  wire jtl_350sxkk00uc2pqvyi24m = (ce4pb74pw07ylxuf649mb4j & ~pp7hxkc1fr9z2qqw) ? 1'b1 : lm7s5990gmfb; 
  wire bpzgy4h2_6osq44grnr60fj_kng = ce4pb74pw07ylxuf649mb4j & pp7hxkc1fr9z2qqw;                       
  wire roq7q8s1jcx19fzuzj42rq6 = n8hk7_wggv11dp5_wcn7kn & jtl_350sxkk00uc2pqvyi24m;
  wire tzwjirxlpok2de1pf4b0dv_sm = bpzgy4h2_6osq44grnr60fj_kng |  roq7q8s1jcx19fzuzj42rq6;
  wire p64hlk6qolmw7ptxce4ugpk = bpzgy4h2_6osq44grnr60fj_kng & ~roq7q8s1jcx19fzuzj42rq6;

  ux607_gnrl_dfflr #(1) nxgldtq251ikmlber37oxh8b_ (tzwjirxlpok2de1pf4b0dv_sm, p64hlk6qolmw7ptxce4ugpk, n8hk7_wggv11dp5_wcn7kn, gf33atgy, ru_wi);

  
  wire x2kr_spj9bwej2jxuua6zok2f5qsb6;
  wire y05m1a51kn2mjz3v1oglw;
  wire ztn79u83h27c1ybfi1uepsxdd = jtl_350sxkk00uc2pqvyi24m;
  wire wxwqnheoa144a8sw669v7yqvf9sl = x2kr_spj9bwej2jxuua6zok2f5qsb6;
  wire mtkvvaodp2cx34eyqxb6dhfr9s3e3i = ztn79u83h27c1ybfi1uepsxdd |  wxwqnheoa144a8sw669v7yqvf9sl;
  wire pvb8v8oubjqouvl48q19jqdzrqa3l = ztn79u83h27c1ybfi1uepsxdd & ~wxwqnheoa144a8sw669v7yqvf9sl;

  ux607_gnrl_dfflr #(1) dzhq525ffai0j0ooq6kzhnfgq50np_l (mtkvvaodp2cx34eyqxb6dhfr9s3e3i, pvb8v8oubjqouvl48q19jqdzrqa3l, y05m1a51kn2mjz3v1oglw, gf33atgy, ru_wi);

  
  wire qkwe_e7cchwb2sjj71c9;
  
  
  wire esgt1gkpa42bbzbwk1u = s_eowfyzlvx7gjv542upo;                                                     
  wire qpmgoal00ptp1ossymtbzuwb = ce4pb74pw07ylxuf649mb4j;                                                
  wire y3v8ih3fb0uruvpaks8f2yyjo = qkwe_e7cchwb2sjj71c9 & esgt1gkpa42bbzbwk1u;
  wire mqb46555ry_d67lk0zwhczfz8 = qpmgoal00ptp1ossymtbzuwb |  y3v8ih3fb0uruvpaks8f2yyjo;
  wire tdmarmur2ohf42egko550xgk = qpmgoal00ptp1ossymtbzuwb & ~y3v8ih3fb0uruvpaks8f2yyjo;

  ux607_gnrl_dfflr #(1) v2k_gixm14cspb7etoo33_6r1_ (mqb46555ry_d67lk0zwhczfz8, tdmarmur2ohf42egko550xgk, qkwe_e7cchwb2sjj71c9, gf33atgy, ru_wi);

  assign j8cjhcuf0m6xjvemdaz = qkwe_e7cchwb2sjj71c9;

  
  wire tvs6nbhqtgdbo_xpu1idjg7;
  wire jyjwqrh40xmfk23zxmtctz0ba4dvn4 = esgt1gkpa42bbzbwk1u;
  wire qxa6k5fdycf_ibc01y494sz03h22 = x2kr_spj9bwej2jxuua6zok2f5qsb6;
  wire hgblpuifivioqo4zbadjuo_jsv = jyjwqrh40xmfk23zxmtctz0ba4dvn4 |  qxa6k5fdycf_ibc01y494sz03h22;
  wire lnqtwnxj6osgnyrbzbu953tzlpt_ = jyjwqrh40xmfk23zxmtctz0ba4dvn4 & ~qxa6k5fdycf_ibc01y494sz03h22;

  ux607_gnrl_dfflr #(1) i2prukk8rt9n9vmjs1odbuxj3ikp24wu (hgblpuifivioqo4zbadjuo_jsv, lnqtwnxj6osgnyrbzbu953tzlpt_, tvs6nbhqtgdbo_xpu1idjg7, gf33atgy, ru_wi);

  assign umc_2tn6um_9xaiy7_ksg0w = vaiscz5bqo4k6ql0519;
  assign q7ru87fmzxczveihcxcwh = uuuoq6te8sq6lj_e02iqoc;
  assign uiyh4da4134sjv7gnmc = w93is2iaq5aikcpaqxg3;

  
  assign x2kr_spj9bwej2jxuua6zok2f5qsb6 =   y05m1a51kn2mjz3v1oglw
                                        & tvs6nbhqtgdbo_xpu1idjg7
                                         ;

  assign azqy5qfm4kwm7vkwu6e =   x2kr_spj9bwej2jxuua6zok2f5qsb6;


  
  
  
  
  
  
  
  
  
  
  wire jzqhfc_ru__vhwkz46_3 = qmd94avv02av64cbwaj42 & ~t57d026x085pay & ~vyneby1uawco; 

  
  wire y75xeozj0wna88fi2;
  wire nstpz1tj94vlp30tb2ue = jzqhfc_ru__vhwkz46_3;
  wire iqr6gddiie5aaaztsgvdsbxs = y75xeozj0wna88fi2;
  wire bpyvvs5gutks6ssip3qajy6 = nstpz1tj94vlp30tb2ue | iqr6gddiie5aaaztsgvdsbxs;
  wire jrqc49ty9zwxqm2biw0g2q8 = nstpz1tj94vlp30tb2ue & ~iqr6gddiie5aaaztsgvdsbxs;

  ux607_gnrl_dfflr #(1) j4o8xuw6t3hkf_x5k8_tk17gim (bpyvvs5gutks6ssip3qajy6, jrqc49ty9zwxqm2biw0g2q8, y75xeozj0wna88fi2, gf33atgy, ru_wi);

  
  assign d40pep591l63yhmefp7i = y75xeozj0wna88fi2;

  
  wire nyft8x6dvpm34sgx0ay0 = jzqhfc_ru__vhwkz46_3;
  wire ez6a1xb6d192zis12z5ra = k5th293qdrtsytaehbsk;
  wire f78v5l7opria5y3pjhti = nyft8x6dvpm34sgx0ay0 |  ez6a1xb6d192zis12z5ra;
  wire y68n1g03hkb7ehwwagr1 = nyft8x6dvpm34sgx0ay0 & ~ez6a1xb6d192zis12z5ra;

  ux607_gnrl_dfflr #(1) jui86zege1565jl_8e6gcm8gt (f78v5l7opria5y3pjhti, y68n1g03hkb7ehwwagr1, t57d026x085pay, gf33atgy, ru_wi);

  
  assign g6gwjq519o1w1m3csgrrf3   = t57d026x085pay & m4ndmqnlr5eisc8m2k6fd;
  assign lo_2ny7_v71by78q3         = jcczlhzxqzl5dx51l;
  assign hbdj3fcr8qkfkgzq58o1o2ozh = t57d026x085pay & nkdn__tk5pvp4nczp7xysy5;
  assign m_k_n75bb0f_im9fu_       = fhzpp1p52pmfd3syoo;

  assign hv9e7_hu5oyc6e87832pmb    = k5th293qdrtsytaehbsk;


  wire kva0dtfrzw769eb = (fb2yieg4ys3p19gmk96ooyq66 & (~lm7s5990gmfb) & (~vyneby1uawco)); 

  wire [7-1:0] e1a8llu4i0eq;
  wire rofqn5vmqgj3 = (~jlihkmvsqt_p1_x) & ( 
      
         raha4wzwsh_g_zg
      
         | kva0dtfrzw769eb
         );
  wire wb2d7lcanso_if = jlihkmvsqt_p1_x;
  wire e76n14px0ratq4_ = rofqn5vmqgj3 | wb2d7lcanso_if;
  wire [7-1:0] wg62qey3bgbqfj3d5 = 
                                   rofqn5vmqgj3 ? {7{1'b0}}
                                 : wb2d7lcanso_if ? (e1a8llu4i0eq + {{7-1{1'b0}},1'b1})
                                 : e1a8llu4i0eq;
  
  ux607_gnrl_dfflr #(7) qboluq6i0kgda042d0s (e76n14px0ratq4_, wg62qey3bgbqfj3d5, e1a8llu4i0eq, gf33atgy, ru_wi);
  
  localparam x_g7_amp9xm4fxdr52ks60ap = (128 -1);
  wire tgvigiz1id3yq74ap7a = rofqn5vmqgj3;
  wire wx1aad1kfoyvalpt74 = (e1a8llu4i0eq == x_g7_amp9xm4fxdr52ks60ap[7-1:0]);
  wire r79h9xnmvtiwcs5 = tgvigiz1id3yq74ap7a |   wx1aad1kfoyvalpt74;
  wire dda72ysm66bqae = tgvigiz1id3yq74ap7a | (~wx1aad1kfoyvalpt74);
  ux607_gnrl_dfflr #(1) g1f9nu4pykh3rvv70 (r79h9xnmvtiwcs5, dda72ysm66bqae, jlihkmvsqt_p1_x, gf33atgy, ru_wi);
  
  wire su138bbockj4qe1u = fb2yieg4ys3p19gmk96ooyq66 & wx1aad1kfoyvalpt74;
  wire fbm89oqzpf485u = lm7s5990gmfb;
  wire crmc1rsdybc9ge4qsr5 = su138bbockj4qe1u |   fbm89oqzpf485u;
  wire lfpcr5qjru5aaf8y3 = su138bbockj4qe1u | (~fbm89oqzpf485u);
  ux607_gnrl_dfflr #(1) vp5qn6e7y0_so4m9yo (crmc1rsdybc9ge4qsr5, lfpcr5qjru5aaf8y3, lm7s5990gmfb, gf33atgy, ru_wi);
  
  assign e4exh90ggokeh = tgvigiz1id3yq74ap7a | jlihkmvsqt_p1_x;
  
  wire xqihtrwb2rux = wb2d7lcanso_if;
  wire zm10o_ok84f1a2a = 1'b1;
  wire [7-1:0] hkzt7_zvbwxs8pg = e1a8llu4i0eq;
  wire [54-1:0] twcou1u_kor0c6xc  = {54{1'b0}};
  

  wire klkflmsyyf5w7ar; 
  wire wy36iirxspfw56864;
  wire lkjqs6kiuyj; 
  wire sxxoah7zbvh8noti; 
  wire wgls7kw8r0vwnfoaa5; 
  wire rxb8t16amctwwc; 
  wire [64-1:0] h7f6k_ims_9p3; 

  wire  c86b14qr2qo45_qw2ns;

  wire h5maomnmovgqtb7 = th06du2c8e2_b7k & irjoi8wvo25u209f_5;

  wire [64-1:0]           r74gcroj00so8fhld15kw;
  wire                                 m79e4y4bxjv8wjf92v;
  wire                                 sdiutxggk1c2ak7ktdrdb;
  wire                                 cc6qwrad4apslaurcpws7k;
  wire                                 yvi4x0op9l363_sn0wyyawr;
  assign r74gcroj00so8fhld15kw  = tlmb65lrny6own ? nkj14m5ilghbj  : zvk11dhgg2s67mkq;
  assign sdiutxggk1c2ak7ktdrdb = tlmb65lrny6own ? qqz76r4390y_pzoug : qaidts35dk5jcji0n;
  assign cc6qwrad4apslaurcpws7k = tlmb65lrny6own ? r96xqbs4rp4ud91vy : fbzs0o4ysyuzeg_qdj;
  assign yvi4x0op9l363_sn0wyyawr = tlmb65lrny6own ? ha3mzwrvohf1v4m9 : me1n4pvwxa7n3u8l05;
  assign m79e4y4bxjv8wjf92v = tlmb65lrny6own ? 1'b0           : r8nzx6_1no31zeloft;

  wire [5-1:0]      o44qsljzqi70j2c9ld    = r74gcroj00so8fhld15kw[4:0];
  wire [59-1:0]   gep338whtkvmcn2qzgt_7rp = r74gcroj00so8fhld15kw[(64-1):5];

  wire [7-1:0]      nrpgu15ovg_qfow2s14 = gep338whtkvmcn2qzgt_7rp[7-1:0];
  wire [52-1:0]        c2whp6v0rnjcid3g9gf = gep338whtkvmcn2qzgt_7rp[59-1:7];

  wire aoteh1s7gdbchnl8m;

  wire dcj485cah5;
  wire peo2y31x_joi;

  wire e0ccmihftf2h7qp1bb4m;
  wire pexht3mjwe9iclbm;
  
  wire xd1hp6jei8rpmhpkg_sl =  1'b0 
                             
                             ;
  wire zudemjr0ci807luhc;
  wire vz5nhqfrpq1hoj;
  wire [7-1:0] kqqo4t7wgbicepuzlzgoe8;
  wire [54-1:0] bg33yeiaa_koh0mtr7f2;

  wire z983juq6oh_0wb;
  wire fi44ix6nhyef6;
  
  
  
  
  
  
  assign e0ccmihftf2h7qp1bb4m = z983juq6oh_0wb;
  assign pexht3mjwe9iclbm = fi44ix6nhyef6;
  



  wire [7-1:0] jm9hjt3oqbob590sdfe;
  wire [54-1:0] wb4vwdrejqmlx7swh7a_0b;

  wire rjy1mb7tnflt7ea;  
  wire hxztlrjkqickn6urw;

  wire eckc0ni49znxd84c2epuu3v = (~aoteh1s7gdbchnl8m) &  
                            (~dcj485cah5) &         
                            h5maomnmovgqtb7;          
  wire ex9kj5aqz1c8t_s5qt32 =   h5maomnmovgqtb7 
                             & (~dcj485cah5) 
                             ;
  wire [9-1:0] twci9ec7780eeo = {nrpgu15ovg_qfow2s14,o44qsljzqi70j2c9ld[5-1:3]};
  
  wire [59-1:0]   yalj29s91xhsqm2mjvz9dtnq39t = zvk11dhgg2s67mkq[(64-1):5];
  wire [7-1:0]      vbbu0tudbtb03g7jz78r4gu = yalj29s91xhsqm2mjvz9dtnq39t[7-1:0];
  wire [7-1:0]   bnxmgh9k7tgknk6p1yl8g = vbbu0tudbtb03g7jz78r4gu;

  
  wire [59-1:0]   cchx3mkgg7dd8kkwcg3f7enkvsy = nkj14m5ilghbj[(64-1):5];
  wire [7-1:0]      vmrcuch33vluqwki8tsnvmbli8 = cchx3mkgg7dd8kkwcg3f7enkvsy[7-1:0];
  wire [7-1:0]   bqoquiu_sr0myw0y4tow = vmrcuch33vluqwki8tsnvmbli8;

  wire l7sauvhwo7orvwq0tz6tql;
  wire gsf_5l61c1nvvp_;
  wire [7-1:0] akg6apmoz04bjkagrh;
  wire [54-1:0] fxu0h92n3g4evsus;
  
  
  wire b88tuttz2asy0vv3oo4x0k =  ~(e4exh90ggokeh | l7sauvhwo7orvwq0tz6tql | e0ccmihftf2h7qp1bb4m | pexht3mjwe9iclbm | peo2y31x_joi);
  assign ldqpjrsj9dp8yg3uc   = e4exh90ggokeh ? xqihtrwb2rux   : (l7sauvhwo7orvwq0tz6tql | eckc0ni49znxd84c2epuu3v | e0ccmihftf2h7qp1bb4m | pexht3mjwe9iclbm | peo2y31x_joi);
  assign s70e4xdis3p67ndpn6fbx   = b88tuttz2asy0vv3oo4x0k ? 1'b0                            : e4exh90ggokeh ? zm10o_ok84f1a2a   :  l7sauvhwo7orvwq0tz6tql ? gsf_5l61c1nvvp_   : e0ccmihftf2h7qp1bb4m ? 1'b0          : peo2y31x_joi ? rjy1mb7tnflt7ea       : zudemjr0ci807luhc;
  assign h9zlka3j3ih8ihpvwvky1 = b88tuttz2asy0vv3oo4x0k ? bnxmgh9k7tgknk6p1yl8g              : e4exh90ggokeh ? hkzt7_zvbwxs8pg :  l7sauvhwo7orvwq0tz6tql ? akg6apmoz04bjkagrh : e0ccmihftf2h7qp1bb4m ? bqoquiu_sr0myw0y4tow : peo2y31x_joi ? jm9hjt3oqbob590sdfe : kqqo4t7wgbicepuzlzgoe8;
  assign tf_tmpul8i8qbm_djvtl5f  = b88tuttz2asy0vv3oo4x0k ? {54{1'b0}} : e4exh90ggokeh ? twcou1u_kor0c6xc  :  l7sauvhwo7orvwq0tz6tql ? fxu0h92n3g4evsus  : e0ccmihftf2h7qp1bb4m ? {54{1'b0}} : peo2y31x_joi ? wb4vwdrejqmlx7swh7a_0b : bg33yeiaa_koh0mtr7f2;
  
  
  wire rj69sa3044rb1cz6lvd6;
  wire atpyq4kwa38ur5a1v4jxl;

  wire r5947sq0alkh4q;
  wire [9-1:0] g7c1415q8kv_x6ed0;
  wire [64-1:0] dkn8bvcvpdmu34 ;
  

  
  assign w0ve66vjdz8lzwws3ic   = (rj69sa3044rb1cz6lvd6 | ex9kj5aqz1c8t_s5qt32);
  assign df775k2ts6dn4528iq_ce5   = rj69sa3044rb1cz6lvd6 ? r5947sq0alkh4q   : 1'b0;
  assign k3dychuj1pv4vw7cfj01ft8v = rj69sa3044rb1cz6lvd6 ? g7c1415q8kv_x6ed0 : twci9ec7780eeo;
  assign jh4zf96qrsb31j072n  = rj69sa3044rb1cz6lvd6 ? dkn8bvcvpdmu34  : {64{1'b0}};
  
  
  
  wire d3j_g8wp81xd22uqe66u;  
  
  wire gnvikxdm0vcpzqnzpygul5o45 =  ~(e4exh90ggokeh | d3j_g8wp81xd22uqe66u | e0ccmihftf2h7qp1bb4m | pexht3mjwe9iclbm | peo2y31x_joi);
  assign hv6xxz3oswj4wy4j46   = e4exh90ggokeh ? xqihtrwb2rux   : (d3j_g8wp81xd22uqe66u | eckc0ni49znxd84c2epuu3v | e0ccmihftf2h7qp1bb4m | pexht3mjwe9iclbm);
  assign q6p7kcdd9o7j3e2c886   = gnvikxdm0vcpzqnzpygul5o45 ? 1'b0                            : e4exh90ggokeh ? zm10o_ok84f1a2a   :  d3j_g8wp81xd22uqe66u ? gsf_5l61c1nvvp_   : e0ccmihftf2h7qp1bb4m ? 1'b0          : peo2y31x_joi ? hxztlrjkqickn6urw       : vz5nhqfrpq1hoj;
  assign ee_yaeclihal4dht69liwy6z = gnvikxdm0vcpzqnzpygul5o45 ? bnxmgh9k7tgknk6p1yl8g              : e4exh90ggokeh ? hkzt7_zvbwxs8pg :  d3j_g8wp81xd22uqe66u ? akg6apmoz04bjkagrh : e0ccmihftf2h7qp1bb4m ? bqoquiu_sr0myw0y4tow : peo2y31x_joi ? jm9hjt3oqbob590sdfe : kqqo4t7wgbicepuzlzgoe8;
  assign thl4cxcuzntax8hnsn9bl4  = gnvikxdm0vcpzqnzpygul5o45 ? {54{1'b0}} : e4exh90ggokeh ? twcou1u_kor0c6xc  :  d3j_g8wp81xd22uqe66u ? fxu0h92n3g4evsus  : e0ccmihftf2h7qp1bb4m ? {54{1'b0}} : peo2y31x_joi ? wb4vwdrejqmlx7swh7a_0b : bg33yeiaa_koh0mtr7f2;
  
  
  assign vp3x08mx4e27x4k26n   = (atpyq4kwa38ur5a1v4jxl | ex9kj5aqz1c8t_s5qt32);
  assign a7b829uahvy2i28yzgg   = atpyq4kwa38ur5a1v4jxl ? r5947sq0alkh4q   : 1'b0;
  assign kzxrmeg90fb06oya08h1 = atpyq4kwa38ur5a1v4jxl ? g7c1415q8kv_x6ed0 : twci9ec7780eeo;
  assign kl5wycr14v5ukl7oqfhwe6  = atpyq4kwa38ur5a1v4jxl ? dkn8bvcvpdmu34  : {64{1'b0}};
  
  


 wire x00j30a6s29yi = 
               | nywm0kv90g64r5310wz
               | e4exh90ggokeh        
               | f48_2zc1qro_3dodmk8  
               | qmd94avv02av64cbwaj42 
               ;
     
     



 wire zs89k7qgupd1xlvx63l2r;
 wire v43e726lsk4q8y4jnic;
 wire mz_exhb6gtbcmmad884;
 assign wz_if_2q_23jhl2 = uz8uoctou96a_0m95zx | vyneby1uawco | th06du2c8e2_b7k  
                      | f48_2zc1qro_3dodmk8  
                      | gysg24e47c3aqwd9wkc7m  
                      | zs89k7qgupd1xlvx63l2r  
                      | (~mz_exhb6gtbcmmad884)  
                      | (~v43e726lsk4q8y4jnic)  
                      | qmd94avv02av64cbwaj42  
                      | tlmb65lrny6own  
                      ;

 wire k1by1np3;
 wire ax1mncgjkrzn;
 wire cu3vv6uz5iff;

 wire jy8uskaamz5hsuj8mmvvc; 
 wire k6crim9kra7e8x1l; 
 wire ub__mzukp2wlfwg; 
 wire lh5iofwlh72_4 = ~jy8uskaamz5hsuj8mmvvc;
 wire kdkn39pg0ldyc23un = tlmb65lrny6own & k6crim9kra7e8x1l;  
 assign k1by1np3      = (~x00j30a6s29yi) & ((th06du2c8e2_b7k & (~tlmb65lrny6own)) | kdkn39pg0ldyc23un) & (~peo2y31x_joi);
 assign irjoi8wvo25u209f_5 = (~x00j30a6s29yi) & ax1mncgjkrzn & (~peo2y31x_joi)
                      & (~tlmb65lrny6own)                     
                        ;

 wire s9hgy6syn2arl9fxs8kb0 = rinamilgle00i5xmx_vt & j8wlfupbw25hdmohz5q0;
 wire jetszpnn_3n3x0k4d = klkflmsyyf5w7ar & wy36iirxspfw56864;
 wire v_x8q3x575_d2wk1peosi7 = ze2bfnigu62i9937pcxnjc & c86b14qr2qo45_qw2ns;

 
 wire tadam78rmm5zsv = cc6qwrad4apslaurcpws7k | sdiutxggk1c2ak7ktdrdb | dep51yq;





 assign dcj485cah5 = lh5iofwlh72_4 ? 1'b0 : (~pp7hxkc1fr9z2qqw) ? 1'b1 : sdiutxggk1c2ak7ktdrdb ? 1'b1 : 1'b0;
 localparam bu7gxwekpym = 64+5+1
                         + 1
                         + 1
                       ;

 wire [bu7gxwekpym-1:0] hgv6e1dphu;
 wire [bu7gxwekpym-1:0] xbookicei5na;
 wire t3tudcq0j;
 wire vcalsdo6q;
 wire gj5_lf5d5ejxyzhli9;
 wire v3aoq66fpdwia80or5l;
 wire v5wwz2lnt_lzr76xz2;
 wire ucjjrmorqafl;
 wire z5oodn6lsltcchb6;
 wire w_45r8lsw7umpt;
 wire dd8s8azwnmm78;
 wire mu_grj5_po0a4ek;
 wire ik4xc_1hh4vb;
 wire p8jjix1l0zn0yr760;
 wire [64-1:0] dm_t8xh6s80cssm; 
 wire [7-1:0] pkmbkt_zq0yhlemrgi;
 wire [52-1:0]   jcbv86t6ccbny9um2sm;
 assign hgv6e1dphu = {
                    lh5iofwlh72_4,
                    tadam78rmm5zsv,
                    dcj485cah5,
                    m79e4y4bxjv8wjf92v,
                    cc6qwrad4apslaurcpws7k,
                    sdiutxggk1c2ak7ktdrdb,
                    yvi4x0op9l363_sn0wyyawr,
                    aoteh1s7gdbchnl8m,
                    r74gcroj00so8fhld15kw};
 assign {
     ub__mzukp2wlfwg,
     t3tudcq0j,
     gj5_lf5d5ejxyzhli9,
     mu_grj5_po0a4ek,
     z5oodn6lsltcchb6,
     ik4xc_1hh4vb,
     w_45r8lsw7umpt,
     p8jjix1l0zn0yr760,
     dm_t8xh6s80cssm} = xbookicei5na;
  wire o1w7damum_chn0d2y;

  wire [64-1:0] axng6pw6x_ngow1o7_7e;

wc2lipjaiimwuy7fx9zp32mr  lbpbwc1x5lhcs71rg3inpdi1d2xu(
     .e98zc_xde8d   (axng6pw6x_ngow1o7_7e[32-1:0]),
     .lms849k     (v3aoq66fpdwia80or5l),
     .dhzk00cwbk (v5wwz2lnt_lzr76xz2)
  );

  assign ucjjrmorqafl = v5wwz2lnt_lzr76xz2 & (~ik4xc_1hh4vb);


  wire aknbc4862andzqg1530a;
  assign vcalsdo6q =   gj5_lf5d5ejxyzhli9 
                    | (v3aoq66fpdwia80or5l & (t3tudcq0j ? 1'b1 : aknbc4862andzqg1530a))
                    ;

  
  
    localparam xio4kx7ep1ojwa_r = 51;
    localparam cmnocc9r2aiw8za  = 8;
    localparam xholqktr732apzsv8d0 = 3;

    wire                           hq6v70g7_oxcoxo;
    wire                           tshed5u3v36qsn;
    wire [27-1:0] scyket9x073uq5f;
    
    
    wire [20-1:0] wp81q9t8ggv2_3x2;
    
    
    wire                           kobvr2up44i45y3z;
    wire                           mi1x48jare2xkb4w8p550kcadl6;
    wire                           oqf10y60u0sj6773kobz81we1znk;
    wire                           ylm6yo9kkk2s745bw1ay;
    wire                           x_lssc66vaunqx1;
    wire                           wal48n0a3elwnwyud8i3jmv;
    wire                           x3vfczxmitp90acekkojua;
    wire                           dnlcindr8ja4jikk;
    wire [26-1:0]  k7nob8irhm5ucjhtgm230et; 
    wire                           ebjxpmm7zy2qjn994pkq3d;
    wire [1:0]                     n0c39kkvp4h6ula91p; 

    assign hq6v70g7_oxcoxo = k1by1np3 & ax1mncgjkrzn;
    assign tshed5u3v36qsn = hq6v70g7_oxcoxo & (~tadam78rmm5zsv);
    assign scyket9x073uq5f = r74gcroj00so8fhld15kw[64-26 : 64-26-27+1]; 

    assign k7nob8irhm5ucjhtgm230et = dm_t8xh6s80cssm[64-1: 64-26];
    assign ebjxpmm7zy2qjn994pkq3d =   (k7nob8irhm5ucjhtgm230et != {26{1'b1}}) 
                                    & (k7nob8irhm5ucjhtgm230et != {26{1'b0}})
                                    ;

    
    
    
    
    
    
    assign wal48n0a3elwnwyud8i3jmv =   mi1x48jare2xkb4w8p550kcadl6 
                                | (~z5oodn6lsltcchb6 & ~w_45r8lsw7umpt & ~ik4xc_1hh4vb & ~kobvr2up44i45y3z & ~oqf10y60u0sj6773kobz81we1znk) 
                                | (~z5oodn6lsltcchb6 &  w_45r8lsw7umpt & ~ik4xc_1hh4vb &  kobvr2up44i45y3z & ~oqf10y60u0sj6773kobz81we1znk) 
                                | (ebjxpmm7zy2qjn994pkq3d)
                                ;
    
    
    
    assign x3vfczxmitp90acekkojua = oqf10y60u0sj6773kobz81we1znk;
    
    
    
    
    
    assign dnlcindr8ja4jikk = vcalsdo6q;
    
    
    
    
    assign n0c39kkvp4h6ula91p = {1'b0,yvi4x0op9l363_sn0wyyawr}; 

  hpwm3nya3 #(
   .xio4kx7ep1ojwa_r     (xio4kx7ep1ojwa_r),
   .cmnocc9r2aiw8za      (cmnocc9r2aiw8za),
   .xholqktr732apzsv8d0 (xholqktr732apzsv8d0)
  )  tf8tyherihphzj2 (
    .mv5to8v6                            (y75xeozj0wna88fi2                    ),
    .k3n1uuckanw669a                    (tshed5u3v36qsn                         ),
    .qfy7pr76nvqld1f                    (scyket9x073uq5f                         ),
    .nowfs1y75z9hmhv6r0ppp6vjly             (n0c39kkvp4h6ula91p                  ),
    .f_8ecse5wf0jrndlozy2070bja             (aknbc4862andzqg1530a                  ),
    
    .c_lxwlogrc590ejlmhjdrmfmj               (wp81q9t8ggv2_3x2                    ),
    
    
    .ugixcggahb26m1glzpuqvpq              (kobvr2up44i45y3z                   ),
    .vbpz6tidsg3o93kih6nmamlyg9wmr1zz        (mi1x48jare2xkb4w8p550kcadl6             ),
    .j2dtuvq0m4iir947lery9tpxqwhjj2g3      (oqf10y60u0sj6773kobz81we1znk           ),
    .wo834bx1b9sidvkaqiq_b7jk             (ylm6yo9kkk2s745bw1ay                  ),
    .faamp7iz46_jj1ci8a                  (x_lssc66vaunqx1                       ),
    .v66ux9ovjkzt3jn                     (wk9s3wmc2q0yaa13                    ),
    .cd3lo77nievm4v3                      (s7re1eyp36bjvie                     ),
    .rgnht1zljy67subvhyua_               (a1pnq3ko2aaldi7h3xwme              ),
    .nmlix317bu48vgct7x02m7vgn               (oq4nxgat71_rnebbasjmv9              ),
    .s6zb15tq6xjiqgce5nwjcg7be4          (rj1ewmv16hujp9xlnpm6a3hhu9y8ml         ),
    .ry0rypry86op3l_hqbwk8pe32ena3e        (ryfblq1f8us1a8u3gy2gijl12x085ja       ), 
    .h4zmq2srkdf5iaeagd8d7i87                (j6q7tn13h_mjup45od1mu               ),
    .dzo70vq3_1_kyxyiurxy1d20ed              (x81uu_gb6esoi095hudjgylqn             ), 
    .b0c0o6unssb9h3tgqck870              (ql2if76ihe_ppb4rp3buw7             ), 
    .c2_546oy8pb0vifo                    (v43e726lsk4q8y4jnic                   ), 
    .gf33atgy                                (gf33atgy                                ),
    .ru_wi                              (ru_wi                              ),
    .gc4b3kdcan6do88ta_                     (gc4b3kdcan6do88ta_                     ) 
  );


  wire [64-1:0] xb37vggkwqec73o   = {{(64-20-12){1'b0}},wp81q9t8ggv2_3x2,dm_t8xh6s80cssm[11:0]};
  assign axng6pw6x_ngow1o7_7e = t3tudcq0j ? dm_t8xh6s80cssm : xb37vggkwqec73o;

  wire gdc31z_ah0g;
  wire vldo6rbn;
  wire vh2j7b0kt7n2s59;
  wire b24yx4ictsbkcpj;
  wire xvnxfgnlx05;
  wire b293miy3ig80jz;
  wire h6yap55ubdbc2;
  wire yz14ncxfv0;
  wire iaaolhc_afh_9est07sqv;

  
  
  

  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  

  localparam v8lpuviyaayisob6gd6b  = 4;
  
  localparam afsd_3qtyoxr7r3 = 4'd0;
  
  localparam rnvbydgv9rjrawrwvg   = 4'd1;
  
  localparam vlpwcdyr8gjljrzocaj  = 4'd2;
  
  localparam np8lmm9f0lgm38   = 4'd3;
  
  localparam mlfpumkewbr06h9 = 4'd4;
  
  localparam daw0j4ce5dqq6tac_3x = 4'd5;
  
  localparam zj5oy4mazgo9wh9x = 4'd6;
  
  localparam as0gdykns7qp74p1v5 = 4'd7;
  
  localparam a84dgj1l2pfccyw_ = 4'd8;

  
  
  wire [v8lpuviyaayisob6gd6b-1:0] bgzt_rw45yxhq99rb36;
  wire [v8lpuviyaayisob6gd6b-1:0] o7fmwngroif0;
  wire ud7a052bl2cgx_;

  wire [v8lpuviyaayisob6gd6b-1:0] u1kckrxxhwuxkfspvd59yq;
  wire [v8lpuviyaayisob6gd6b-1:0] rl1wtat2cxs2ev3eb55;
  wire [v8lpuviyaayisob6gd6b-1:0] da3_gntbvgqv_zwnh76a1;
  wire [v8lpuviyaayisob6gd6b-1:0] afbx7t4n5uyitw02ia5;
  wire [v8lpuviyaayisob6gd6b-1:0] wbboo1t2jqvlu7hvq2shmztb;
  wire [v8lpuviyaayisob6gd6b-1:0] ttdas42zc03dc75jdvgc;
  wire [v8lpuviyaayisob6gd6b-1:0] d7aeg8a362uouq00q0nf7;
  wire [v8lpuviyaayisob6gd6b-1:0] k_vqilrpwrrf3i35kqqor6l;
  wire [v8lpuviyaayisob6gd6b-1:0] pnina70evcktcnps9z4w2k;
  wire b9hc1gjej65emhg1dwdfsbnc;
  wire n0_f6p9ntm2jqlpigf_32wptq3;
  wire sgx0qmcequsitomfo73r_yn;
  wire llpn9i5u8xn1zuk7riwmx3_cgog_;
  wire oyjswan269wye8llb20w4ffe;
  wire v6pcpcfd3o48r9ohc4q6fylq;
  wire dxf8_iddqbp7dzewb_gryj65;
  wire t66ja3ehz1sj30q598igq2x5t;
  wire kf0t5xhv8cyrwr47q76ax5mfyq;
  
  assign jy8uskaamz5hsuj8mmvvc = (o7fmwngroif0 == afsd_3qtyoxr7r3);
  assign k6crim9kra7e8x1l   = (o7fmwngroif0 == rnvbydgv9rjrawrwvg);
  wire cyjoizk175tz59s73g1    = (o7fmwngroif0 == vlpwcdyr8gjljrzocaj);
  wire jl11end_ebzc87k5v    = (o7fmwngroif0 == as0gdykns7qp74p1v5);
  wire s9tpwhywo_9533a_ux   = (o7fmwngroif0 == a84dgj1l2pfccyw_);
  wire cskxranfmzb5vjara58   = (o7fmwngroif0 == mlfpumkewbr06h9);
  wire vpb0cabpdsgj5tv_     = (o7fmwngroif0 == np8lmm9f0lgm38);
  wire h7psrqammllwnecuonz  = (o7fmwngroif0 == daw0j4ce5dqq6tac_3x);
  wire c6gjb7_uolsl4agll02   = (o7fmwngroif0 == zj5oy4mazgo9wh9x);
   
  assign b9hc1gjej65emhg1dwdfsbnc = jy8uskaamz5hsuj8mmvvc & tlmb65lrny6own & ~vyneby1uawco & ~x00j30a6s29yi;
  assign u1kckrxxhwuxkfspvd59yq = wzrv89a8lbkafx2qdx ? daw0j4ce5dqq6tac_3x : rnvbydgv9rjrawrwvg;
  
  assign n0_f6p9ntm2jqlpigf_32wptq3 = k6crim9kra7e8x1l;
  assign rl1wtat2cxs2ev3eb55 = vlpwcdyr8gjljrzocaj;
  
  wire smqoz2oj8ww5don;
  wire l_razgaao587019p;
  wire u7ja7msr33bxl;
  wire dh_clbn0o20fgf4;
  wire iq0t6kp6qfri0qe61w;

 wire [7-1:0] v94hbvyskjuea4n7wsw4d;
 wire [52-1:0]   wfvfwnnky0p7at5zp07vtk;
  wire egsj_v4pl_4;    
  wire wo2xz_n9y7nkzka;    
  wire vkhotkpp9yeqfbubp;    
  wire mhd_d53mz4u2o78ojq;    
  wire tqd1xxmvx9svwxcdh32;    
  wire fdjtu3kedjy4crxuyi;
  wire nd_hcfia24v6mp0zx;   
  wire z1gnqpih0tzo73j7opinl;
  wire va1c1blelsdo93uz;
  wire cwxkjxgleg8vuggc_nh2xt8c;
  
 wire [7-1:0] zug6nwomkc29qfxbzdpocn;
 wire [52-1:0]   d9hprjtpa534yd5p17wt33b9h;
  wire rng0m4_qo_00;    
  wire zbshs61j683bajzde;    
  wire zej0zy3isij_80da;    
  wire tr3x6j926x74p00e;    
  wire luex4fm_4zh4bo58e1b4l;    
  wire wtbx6tgxz2r4ze7xt;
  wire c3pqxq1ukkc352nk;   
  wire kw97mqedpw8dwl56q6_zx5;
  wire hkvmg02232a2c9zb;
  wire duy9wppkj4is5xqmehcjyu6;
  

  assign l_razgaao587019p = (smqoz2oj8ww5don & b293miy3ig80jz);
  assign iq0t6kp6qfri0qe61w = (dh_clbn0o20fgf4 & yz14ncxfv0);



















  assign u7ja7msr33bxl =   l_razgaao587019p
                       | iq0t6kp6qfri0qe61w
                       ;
  wire b0nb3z34fjl;
  wire h3gomfxna_id829ebe52k5a09 = cyjoizk175tz59s73g1 & (t3tudcq0j ? 1'b1 : aknbc4862andzqg1530a);

  
  assign sgx0qmcequsitomfo73r_yn = h3gomfxna_id829ebe52k5a09; 
  assign da3_gntbvgqv_zwnh76a1 = as0gdykns7qp74p1v5;

  
  assign llpn9i5u8xn1zuk7riwmx3_cgog_ = jl11end_ebzc87k5v;
  assign afbx7t4n5uyitw02ia5 = a84dgj1l2pfccyw_;

  
  assign oyjswan269wye8llb20w4ffe = s9tpwhywo_9533a_ux &
                                   (
                                     peo2y31x_joi | 
                                     rng0m4_qo_00 | 
                                     zej0zy3isij_80da | 
                                    (zbshs61j683bajzde & c4197epxq1j27j_)    |
                                    (zbshs61j683bajzde & vkt5l8auhc9hkqf)   |
                                    (zbshs61j683bajzde & h8yhw0bhacd77xw) 
                                   );
  assign wbboo1t2jqvlu7hvq2shmztb =
                              (rng0m4_qo_00  &  tr3x6j926x74p00e)                                                             ? zj5oy4mazgo9wh9x :
                              (zej0zy3isij_80da )                                                                             ? zj5oy4mazgo9wh9x :
                              (peo2y31x_joi )                                                                                  ? zj5oy4mazgo9wh9x : 
                              (rng0m4_qo_00  & ~tr3x6j926x74p00e & vkt5l8auhc9hkqf   & ~luex4fm_4zh4bo58e1b4l & ~wtbx6tgxz2r4ze7xt)   ? np8lmm9f0lgm38   :
                              (rng0m4_qo_00  & ~tr3x6j926x74p00e & vkt5l8auhc9hkqf   & ~luex4fm_4zh4bo58e1b4l &  wtbx6tgxz2r4ze7xt)   ? zj5oy4mazgo9wh9x :
                              (rng0m4_qo_00  & ~tr3x6j926x74p00e & vkt5l8auhc9hkqf   &  luex4fm_4zh4bo58e1b4l & ~wtbx6tgxz2r4ze7xt)   ? zj5oy4mazgo9wh9x :
                              (rng0m4_qo_00  & ~tr3x6j926x74p00e & vkt5l8auhc9hkqf   &  luex4fm_4zh4bo58e1b4l &  wtbx6tgxz2r4ze7xt)   ? zj5oy4mazgo9wh9x :
                              (zbshs61j683bajzde                    & vkt5l8auhc9hkqf   & ~luex4fm_4zh4bo58e1b4l)                       ? mlfpumkewbr06h9 :
                              (zbshs61j683bajzde                    & vkt5l8auhc9hkqf   &  luex4fm_4zh4bo58e1b4l)                       ? zj5oy4mazgo9wh9x :
                              (rng0m4_qo_00  & ~tr3x6j926x74p00e & c4197epxq1j27j_)                                              ? np8lmm9f0lgm38   :
                              (zbshs61j683bajzde                    & c4197epxq1j27j_)                                              ? zj5oy4mazgo9wh9x :
                              (rng0m4_qo_00  & ~tr3x6j926x74p00e & h8yhw0bhacd77xw &  wtbx6tgxz2r4ze7xt)                       ? np8lmm9f0lgm38   : 
                              (rng0m4_qo_00  & ~tr3x6j926x74p00e & h8yhw0bhacd77xw & ~wtbx6tgxz2r4ze7xt)                       ? zj5oy4mazgo9wh9x : 
                              (zbshs61j683bajzde                    & h8yhw0bhacd77xw)                                           ? zj5oy4mazgo9wh9x :
                              zj5oy4mazgo9wh9x;

  assign v6pcpcfd3o48r9ohc4q6fylq = cskxranfmzb5vjara58 & zs89k7qgupd1xlvx63l2r & iaaolhc_afh_9est07sqv;
  assign ttdas42zc03dc75jdvgc = zj5oy4mazgo9wh9x;
  
  assign dxf8_iddqbp7dzewb_gryj65 = vpb0cabpdsgj5tv_;
  assign d7aeg8a362uouq00q0nf7 = zj5oy4mazgo9wh9x;
  
  assign t66ja3ehz1sj30q598igq2x5t = h7psrqammllwnecuonz & lm7s5990gmfb;
  assign k_vqilrpwrrf3i35kqqor6l = zj5oy4mazgo9wh9x;
  assign lh8ggdb3m21qvo0q = h7psrqammllwnecuonz;
  
  assign kf0t5xhv8cyrwr47q76ax5mfyq = c6gjb7_uolsl4agll02;
  assign pnina70evcktcnps9z4w2k = afsd_3qtyoxr7r3;
  
  assign ud7a052bl2cgx_ =   b9hc1gjej65emhg1dwdfsbnc
                          | n0_f6p9ntm2jqlpigf_32wptq3
                          | sgx0qmcequsitomfo73r_yn
                          | llpn9i5u8xn1zuk7riwmx3_cgog_
                          | oyjswan269wye8llb20w4ffe
                          | v6pcpcfd3o48r9ohc4q6fylq
                          | dxf8_iddqbp7dzewb_gryj65
                          | t66ja3ehz1sj30q598igq2x5t
                          | kf0t5xhv8cyrwr47q76ax5mfyq
                          ;
  
  assign bgzt_rw45yxhq99rb36 =   ({v8lpuviyaayisob6gd6b{b9hc1gjej65emhg1dwdfsbnc  }} & u1kckrxxhwuxkfspvd59yq)
                          | ({v8lpuviyaayisob6gd6b{n0_f6p9ntm2jqlpigf_32wptq3    }} & rl1wtat2cxs2ev3eb55)               
                          | ({v8lpuviyaayisob6gd6b{sgx0qmcequsitomfo73r_yn   }} & da3_gntbvgqv_zwnh76a1)               
                          | ({v8lpuviyaayisob6gd6b{llpn9i5u8xn1zuk7riwmx3_cgog_   }} & afbx7t4n5uyitw02ia5)               
                          | ({v8lpuviyaayisob6gd6b{oyjswan269wye8llb20w4ffe  }} & wbboo1t2jqvlu7hvq2shmztb)               
                          | ({v8lpuviyaayisob6gd6b{v6pcpcfd3o48r9ohc4q6fylq  }} & ttdas42zc03dc75jdvgc)               
                          | ({v8lpuviyaayisob6gd6b{dxf8_iddqbp7dzewb_gryj65    }} & d7aeg8a362uouq00q0nf7)               
                          | ({v8lpuviyaayisob6gd6b{t66ja3ehz1sj30q598igq2x5t }} & k_vqilrpwrrf3i35kqqor6l)               
                          | ({v8lpuviyaayisob6gd6b{kf0t5xhv8cyrwr47q76ax5mfyq  }} & pnina70evcktcnps9z4w2k)               
                          ;
  
  ux607_gnrl_dfflr #(v8lpuviyaayisob6gd6b) dv22mdwcbadidwcw1cnoz (ud7a052bl2cgx_, bgzt_rw45yxhq99rb36, o7fmwngroif0, gf33atgy, ru_wi);
  
  
  
  
  
  assign u_g5yts7tlcxo7ykedbqiv4ji0 = c6gjb7_uolsl4agll02;
  
  
  
  
  
  
  wire z0me2kv52n1b2rtx3gulrbp3w = (s9tpwhywo_9533a_ux  & rng0m4_qo_00  & vkt5l8auhc9hkqf &  luex4fm_4zh4bo58e1b4l & ~wtbx6tgxz2r4ze7xt & ~tr3x6j926x74p00e);
  wire mtah0hwbkrxixd8lp7tdo021g6ge = (s9tpwhywo_9533a_ux  & zbshs61j683bajzde & vkt5l8auhc9hkqf &  luex4fm_4zh4bo58e1b4l & ~tr3x6j926x74p00e);
  
  wire fcum8eje8_3cdlx773gn9a =  z0me2kv52n1b2rtx3gulrbp3w
                               | mtah0hwbkrxixd8lp7tdo021g6ge
                               
                               ;
  wire g0i48rjigmu5_sioztkt8o80 = c6gjb7_uolsl4agll02;  
  wire laf_onfam7bjqrk6xs5sxis = fcum8eje8_3cdlx773gn9a | g0i48rjigmu5_sioztkt8o80;
  wire rmhn596kc4q_c_h1ooz76im = fcum8eje8_3cdlx773gn9a | (~g0i48rjigmu5_sioztkt8o80);
  wire r8zovw2or06kczmgdxhwpm03;
  
  ux607_gnrl_dfflr #(1) hmuonof1oan_22dfykkmahy8oj2 (laf_onfam7bjqrk6xs5sxis, rmhn596kc4q_c_h1ooz76im, r8zovw2or06kczmgdxhwpm03, gf33atgy, ru_wi);
  
  assign qdiqiuzopx36bi3s6fbh7mc16h2cj0 = r8zovw2or06kczmgdxhwpm03 | (|urdbh4qug0s4u_dxqek3ejkxxgejj);

  
  wire lgg2u7pece1k446wk = h3gomfxna_id829ebe52k5a09;
  
  wire bbty43k640bvzf8gmxzo6gtr = lgg2u7pece1k446wk;
  wire b0445ky_wlb2ppb03r4fyd6hnb = c6gjb7_uolsl4agll02;
  wire w943ko5nlylz_ptgccfgcp5a47 = bbty43k640bvzf8gmxzo6gtr | b0445ky_wlb2ppb03r4fyd6hnb;
  wire nz82079sh4nv2v_13hk6hk89_92v = bbty43k640bvzf8gmxzo6gtr ? sxxoah7zbvh8noti : 1'b0;
  wire g3cs02xc407ynr7417_2so6;
  
  ux607_gnrl_dfflr #(1) br3h351_on6_j1j90t99jdrlsc (w943ko5nlylz_ptgccfgcp5a47, nz82079sh4nv2v_13hk6hk89_92v, g3cs02xc407ynr7417_2so6, gf33atgy, ru_wi);
  
  wire a9_padjil63rulm7wwm4ph7wlur2d = g3cs02xc407ynr7417_2so6;


  
  wire ltpp_o9uj91l7ty9f_s0d9g5pm7 = lgg2u7pece1k446wk;
  wire kpfchgtnamutfgb8fpr3_0bo0 = c6gjb7_uolsl4agll02; 
  wire ldlbpkuggu593dncwrhv3n5txj = ltpp_o9uj91l7ty9f_s0d9g5pm7 | kpfchgtnamutfgb8fpr3_0bo0;
  wire nnf0zywkgcjvku61i6tp83msu = ltpp_o9uj91l7ty9f_s0d9g5pm7 ? rxb8t16amctwwc : 1'b0;
  wire gixbcam1z7t3vvzi1wur4yaxw79;
  
  ux607_gnrl_dfflr #(1) t0xz_8bnse22_8b6k_wxrc2ep03vyy (ldlbpkuggu593dncwrhv3n5txj, nnf0zywkgcjvku61i6tp83msu, gixbcam1z7t3vvzi1wur4yaxw79, gf33atgy, ru_wi);
  
  wire ts0keas6eynpk3l9byaw4fy0gkgy20vm = gixbcam1z7t3vvzi1wur4yaxw79;

  
  wire arl2u6_jf5shis627bfda = lgg2u7pece1k446wk;
  wire vbyj81wtowofn93e4a5u = c6gjb7_uolsl4agll02;
  wire ldxgv0ti0l19jdguro3dowfso = arl2u6_jf5shis627bfda | vbyj81wtowofn93e4a5u;
  wire t2lcm197g_w0z76vr6zjnqu = arl2u6_jf5shis627bfda ? vcalsdo6q : 1'b0;  
  wire n2ohn8ezswl65dhw_q6o6z;
  
  ux607_gnrl_dfflr #(1) vslchmehu5leet3e5m1ydydl (ldxgv0ti0l19jdguro3dowfso, t2lcm197g_w0z76vr6zjnqu, n2ohn8ezswl65dhw_q6o6z, gf33atgy, ru_wi);
  
  wire f3993odohbfdgg39mrvyhtz8 = n2ohn8ezswl65dhw_q6o6z;


  
  wire ioc0wmaekzh8ax6wb7o18n8i0h0 = lgg2u7pece1k446wk;
  wire bfeapps_jw_jdcv4eald34t7 = c6gjb7_uolsl4agll02; 
  wire loebzm7mohsm804in7c5ovvuj = ioc0wmaekzh8ax6wb7o18n8i0h0 | bfeapps_jw_jdcv4eald34t7;
  wire csgi8kqysmga0nuwgov9jd5ewkx = ioc0wmaekzh8ax6wb7o18n8i0h0 ? wgls7kw8r0vwnfoaa5 : 1'b0;
  wire xxg_m8not7n4l7wzpmimwu4p;
  
  ux607_gnrl_dfflr #(1) oqjr1cskoyol__v8mbezuagk6mx69 (loebzm7mohsm804in7c5ovvuj, csgi8kqysmga0nuwgov9jd5ewkx, xxg_m8not7n4l7wzpmimwu4p, gf33atgy, ru_wi);
  
  wire lnn96u93upk2ndw5t1ugdpkxr3ngc = xxg_m8not7n4l7wzpmimwu4p;

  
  wire pt7htj1sg7wvma4fcz3m6h45i1 = (cskxranfmzb5vjara58 & zbshs61j683bajzde & vkt5l8auhc9hkqf & ~luex4fm_4zh4bo58e1b4l  & jetszpnn_3n3x0k4d & (vh2j7b0kt7n2s59 & b24yx4ictsbkcpj));
  wire a8t24f6wi1hc8e44p2cwqog0vq = c6gjb7_uolsl4agll02;
  wire s2pau5_2qyovglq356jssxnd0qzb = pt7htj1sg7wvma4fcz3m6h45i1 | a8t24f6wi1hc8e44p2cwqog0vq;
  wire r1ypk8geeq3hvf94npy5w9q7cxs = pt7htj1sg7wvma4fcz3m6h45i1 ? vh2j7b0kt7n2s59 : 1'b0;
  wire seu840wl15adcq49hceoy7z;
  
  ux607_gnrl_dfflr #(1) j6_o_tdpunmonlv2hk5zs2idxm (s2pau5_2qyovglq356jssxnd0qzb, r1ypk8geeq3hvf94npy5w9q7cxs, seu840wl15adcq49hceoy7z, gf33atgy, ru_wi);
  
  wire ntcgludzi7yvanea2lpmzeab9a97 = seu840wl15adcq49hceoy7z;
  
  wire cxnxw5hdq3hknewrmd_3j8y6 = jl11end_ebzc87k5v;
  wire vf_7z446fg5wchupx3n9s75vfb4e = c6gjb7_uolsl4agll02;
  wire nio_p6ibwm0c7wsav14qfwl56y = cxnxw5hdq3hknewrmd_3j8y6 | vf_7z446fg5wchupx3n9s75vfb4e;
  wire o6j1ir4rxpqiv4vc01me6bp4 = cxnxw5hdq3hknewrmd_3j8y6 ? peo2y31x_joi : 1'b0;
  wire my9v93rnvz8cvl5idgdxmtold;
  
  ux607_gnrl_dfflr #(1) t3cj8h5pui0dl_59ez_u_d7y6qp (nio_p6ibwm0c7wsav14qfwl56y, o6j1ir4rxpqiv4vc01me6bp4, my9v93rnvz8cvl5idgdxmtold, gf33atgy, ru_wi);
  
  wire xsphv6i9o4qr9fr90ixku4ugnln7 = my9v93rnvz8cvl5idgdxmtold;


  assign urdbh4qug0s4u_dxqek3ejkxxgejj[0] = r8zovw2or06kczmgdxhwpm03;
  assign urdbh4qug0s4u_dxqek3ejkxxgejj[1] =   a9_padjil63rulm7wwm4ph7wlur2d
                                       | lnn96u93upk2ndw5t1ugdpkxr3ngc
                                       | ts0keas6eynpk3l9byaw4fy0gkgy20vm
                                       | f3993odohbfdgg39mrvyhtz8
                                       ;

  assign urdbh4qug0s4u_dxqek3ejkxxgejj[2] = ntcgludzi7yvanea2lpmzeab9a97;
  assign urdbh4qug0s4u_dxqek3ejkxxgejj[3] = 1'b0;
  assign urdbh4qug0s4u_dxqek3ejkxxgejj[4] = 1'b0;
  assign urdbh4qug0s4u_dxqek3ejkxxgejj[5] = 1'b0;

  
  
  
  
  
  
  
  
  
  
  
  
  
  assign z983juq6oh_0wb = k6crim9kra7e8x1l & ax1mncgjkrzn;
  assign fi44ix6nhyef6 = vpb0cabpdsgj5tv_; 
  
  
  wire j13hzcuptjizy7xbui0u = (cyjoizk175tz59s73g1 & gdc31z_ah0g & vkt5l8auhc9hkqf);
  wire g0dh581gl7ahy_ee9ux1k = (cyjoizk175tz59s73g1 & gdc31z_ah0g & h8yhw0bhacd77xw);
  wire g24q3a57abe1vjbd = (cyjoizk175tz59s73g1 & gdc31z_ah0g & c4197epxq1j27j_);
  wire t36loy84rtvhep1 = j13hzcuptjizy7xbui0u | g0dh581gl7ahy_ee9ux1k | g24q3a57abe1vjbd;
  wire o_zjuagysj4ekq4ov5 = t36loy84rtvhep1;
  wire y8ujfff8f61jrud07 =   (j13hzcuptjizy7xbui0u   & ~b0nb3z34fjl & ~l_razgaao587019p  & b293miy3ig80jz)
                        | (g0dh581gl7ahy_ee9ux1k                &  l_razgaao587019p  & b293miy3ig80jz)  
                        | (g24q3a57abe1vjbd                                      & b293miy3ig80jz)
                        ; 
  wire nzk6svvthgmp0;

  ux607_gnrl_dfflr #(1) u0r96zm6ow7vm_7x_ (o_zjuagysj4ekq4ov5, y8ujfff8f61jrud07, nzk6svvthgmp0, gf33atgy, ru_wi);

  assign zudemjr0ci807luhc = nzk6svvthgmp0;

 
  wire cncemk9avkao4_i28p = t36loy84rtvhep1;
  wire vpxhpom64ykpotd =   (j13hzcuptjizy7xbui0u   & ~b0nb3z34fjl & ~iq0t6kp6qfri0qe61w  & yz14ncxfv0)
                        | (g0dh581gl7ahy_ee9ux1k                &  iq0t6kp6qfri0qe61w  & yz14ncxfv0)  
                        | (g24q3a57abe1vjbd                                      & yz14ncxfv0)
                        ; 
  wire jhha03sfd60mcdpv;

  ux607_gnrl_dfflr #(1) e_j5me3wv61ggou1o (cncemk9avkao4_i28p, vpxhpom64ykpotd, jhha03sfd60mcdpv, gf33atgy, ru_wi);

  assign vz5nhqfrpq1hoj = jhha03sfd60mcdpv;



  
  assign kqqo4t7wgbicepuzlzgoe8 = zug6nwomkc29qfxbzdpocn;

  
  assign bg33yeiaa_koh0mtr7f2 = vkt5l8auhc9hkqf   ? {1'b1, 1'b1, d9hprjtpa534yd5p17wt33b9h} :  
                            h8yhw0bhacd77xw ? {1'b0, 1'b1, d9hprjtpa534yd5p17wt33b9h} :  
                            {1'b0, 1'b0, d9hprjtpa534yd5p17wt33b9h};                     
                            
  

 wire t64aa_wox4xm44t_p; 

  d7stl61zflp21cls1tg e64ki97s_fn9b3w4qea7si2uasbp6kvu (
      .pcr4upio7_tx37     (pcr4upio7_tx37   ), 
      .uzklqlncpqqm1rav  (uzklqlncpqqm1rav),
      .ortueunvnkx_l5m_j  (ortueunvnkx_l5m_j),
      .hwuhtb7ucto_utk56  (hwuhtb7ucto_utk56),
      .i1env2kmns7qvvuuc  (i1env2kmns7qvvuuc),
      .g3s3vpafvy3i  (g3s3vpafvy3i),

      .sxvvsxtbhyvt    (1'b0),
      .rm1dxjejhq7dh3q5m  (1'b0 ),
      .xatytj_r0fv14q  (1'b0 ),

      .oily7    (mu_grj5_po0a4ek),
      .ly3dor8    (1'b0),
      .p1m    (~mu_grj5_po0a4ek),

      .u2k4dyp52s_m(z5oodn6lsltcchb6),
      .bktu0z1mk56(ik4xc_1hh4vb),
      .e98zc_xde8d (axng6pw6x_ngow1o7_7e[32-1:0]),
      .foj6m18  (t64aa_wox4xm44t_p) 
  );

 assign o1w7damum_chn0d2y =   t64aa_wox4xm44t_p
                        & (ub__mzukp2wlfwg ? vkt5l8auhc9hkqf : 1'b1)  
                        ;





  assign dd8s8azwnmm78 = (t3tudcq0j ? o1w7damum_chn0d2y : (o1w7damum_chn0d2y | wal48n0a3elwnwyud8i3jmv | x3vfczxmitp90acekkojua))
                    | ucjjrmorqafl
                    | (t3tudcq0j ? 1'b0 : ylm6yo9kkk2s745bw1ay) 
                    ;

 ux607_gnrl_pipe_stage # (
  .CUT_READY(0),
  .DP(1),
  .DW(bu7gxwekpym)
 ) og14lb1p7094058rm4aft (
   .i_vld(k1by1np3),
   .i_rdy(ax1mncgjkrzn), 
   .i_dat(hgv6e1dphu),
   .o_vld(vyneby1uawco), 
   .o_rdy(cu3vv6uz5iff), 
   .o_dat(xbookicei5na),

   .clk  (gf33atgy  ),
   .rst_n(ru_wi)  
  );

  wire [5-1:0]    m603xpg5m7bwf6h1d    = axng6pw6x_ngow1o7_7e[4:0];
  wire [59-1:0] nf7a14kdh46q_gb4d27t5o = axng6pw6x_ngow1o7_7e[(64-1):5];

    
  wire afyql3m7n_e_;
  assign aoteh1s7gdbchnl8m = afyql3m7n_e_ &    
           (tadam78rmm5zsv == t3tudcq0j) &     
           (~y75xeozj0wna88fi2) &               
           (~dcj485cah5) & (~vcalsdo6q) &  
           (~lh5iofwlh72_4) & (~ub__mzukp2wlfwg) &  
           (~peo2y31x_joi) &                   
           (r74gcroj00so8fhld15kw[(64-1):5] == dm_t8xh6s80cssm[(64-1):5]);  
  
  assign pkmbkt_zq0yhlemrgi = nf7a14kdh46q_gb4d27t5o[7-1:0];
  assign jcbv86t6ccbny9um2sm = nf7a14kdh46q_gb4d27t5o[59-1:7];
  
  wire apmzaxtau_e4j8y = xvnxfgnlx05 & (jcbv86t6ccbny9um2sm == qtsqtuxyont41a7h7i6[52-1:0]);
  assign b293miy3ig80jz = vyneby1uawco & apmzaxtau_e4j8y;

  
  wire mrwckdg2xmt_g4e = h6yap55ubdbc2 & (jcbv86t6ccbny9um2sm == mysqpp41yovfcis6f2dza47[52-1:0]);
  assign yz14ncxfv0 = vyneby1uawco & mrwckdg2xmt_g4e;
  
  

  wire hfltsl05h0c161m131 = (
                                    apmzaxtau_e4j8y 
                                  | mrwckdg2xmt_g4e 
                                  | p8jjix1l0zn0yr760
                                  
                                  
                                  | dd8s8azwnmm78
                                  | (ub__mzukp2wlfwg & (c4197epxq1j27j_ | h8yhw0bhacd77xw | vcalsdo6q)) 
                       );

  assign vldo6rbn =   vyneby1uawco & (~hfltsl05h0c161m131) & mz_exhb6gtbcmmad884
                
                
                
                
                
                
                 & (t3tudcq0j ? (vcalsdo6q ? 1'b0 : 1'b1) : aknbc4862andzqg1530a & (dnlcindr8ja4jikk ? 1'b0 : 1'b1))
                 ; 

  assign gdc31z_ah0g  =   vyneby1uawco &   hfltsl05h0c161m131  & mz_exhb6gtbcmmad884
                
                
                
                
                
                
                 & (t3tudcq0j ? (vcalsdo6q ? dd8s8azwnmm78 | ub__mzukp2wlfwg : 1'b1) : aknbc4862andzqg1530a & (dnlcindr8ja4jikk ? dd8s8azwnmm78 | ub__mzukp2wlfwg : 1'b1))
                 ; 

  wire s2cclwenb  =   vyneby1uawco & mz_exhb6gtbcmmad884
                
                
                
                
                
                
                 & (t3tudcq0j ? (vcalsdo6q ? ~dd8s8azwnmm78 & ~ub__mzukp2wlfwg : 1'b0) : aknbc4862andzqg1530a & (dnlcindr8ja4jikk ? ~dd8s8azwnmm78 & ~ub__mzukp2wlfwg : 1'b0))
                 ; 

  wire rs9cr43eb36gq815zlxyw;
  wire gjkof2a42or0w  =  ze2bfnigu62i9937pcxnjc & rs9cr43eb36gq815zlxyw;

  wire bvs0w3jafe5oum96j06;
  wire swrbe70hp3wsvkt04;

  wire [wq7_4t7xmr99-1:0] y7_io5z_hoy7o_sd1g7q;

  wire ffd_fx0uggmz_c = 
      
          (gdc31z_ah0g & p8jjix1l0zn0yr760) ? bvs0w3jafe5oum96j06 :
      
               gdc31z_ah0g ? b293miy3ig80jz : 
      
               b24yx4ictsbkcpj ? (y7_io5z_hoy7o_sd1g7q[0] == 1'b1) :
                   1'b0;
  wire r2zjd7aqmv0bk_c4 = 
      
          (gdc31z_ah0g & p8jjix1l0zn0yr760) ? swrbe70hp3wsvkt04 :
      
               gdc31z_ah0g ? yz14ncxfv0 : 
      
               b24yx4ictsbkcpj ? (y7_io5z_hoy7o_sd1g7q[1] == 1'b1) :
                   1'b0;

  wire f79jnk8qx3ksw3fem4bpzvg = s9tpwhywo_9533a_ux & zbshs61j683bajzde & vkt5l8auhc9hkqf & ~peo2y31x_joi & ~tr3x6j926x74p00e & luex4fm_4zh4bo58e1b4l;

  assign klkflmsyyf5w7ar = 

                     gdc31z_ah0g
                     
                   | f79jnk8qx3ksw3fem4bpzvg

                   | gjkof2a42or0w

                   | b24yx4ictsbkcpj;

  assign lkjqs6kiuyj = (vh2j7b0kt7n2s59 & b24yx4ictsbkcpj) | (gdc31z_ah0g & dd8s8azwnmm78) | (s2cclwenb & dd8s8azwnmm78) | (gjkof2a42or0w & dm5b92mx0redfbuhs1u3d);

  assign sxxoah7zbvh8noti = t3tudcq0j ? o1w7damum_chn0d2y : 
                                   (
                                      o1w7damum_chn0d2y 
                                    | x3vfczxmitp90acekkojua
                                   ) & ~wal48n0a3elwnwyud8i3jmv; 

  assign rxb8t16amctwwc = (
                             t3tudcq0j ? ucjjrmorqafl & ~o1w7damum_chn0d2y : 
                           ( 
                             ucjjrmorqafl & ~o1w7damum_chn0d2y & ~x3vfczxmitp90acekkojua & ~wal48n0a3elwnwyud8i3jmv
                           ) 
                          ); 

  assign wgls7kw8r0vwnfoaa5 = (t3tudcq0j ? 1'b0 : wal48n0a3elwnwyud8i3jmv);

  assign cu3vv6uz5iff = jetszpnn_3n3x0k4d;

  
  wire [64-1:0] o_p_mo6kcgr0k = ffd_fx0uggmz_c ? vfvtxk4jkkc3ql7_rqd : wt6c82_zmqgmt7if41t698;
  
  wire [64-1:0] ikf61_i17b0iv = o_p_mo6kcgr0k[64-1:0]; 

  assign xvnxfgnlx05 = qtsqtuxyont41a7h7i6[52];
  assign h6yap55ubdbc2 = mysqpp41yovfcis6f2dza47[52];

  assign smqoz2oj8ww5don= xvnxfgnlx05 & qtsqtuxyont41a7h7i6[52+1];
  assign dh_clbn0o20fgf4= h6yap55ubdbc2 & mysqpp41yovfcis6f2dza47[52+1];
  assign b0nb3z34fjl = smqoz2oj8ww5don | dh_clbn0o20fgf4;







  localparam psxtg_0xr2lkj4049fu  = 3;

  localparam uk1oi33ntqrycsuxu = 3'd0;

  localparam dcmmvnhb4tmumn60lcp4  = 3'd1;

  localparam dsix6p9ipz7r85mja3fr  = 3'd2;

  localparam ulyzdpaocwknytnebndi  = 3'd3;

  localparam ojf5u64xjqjjuk3p  = 3'd4;

  localparam f6n2huuf8s7hdk3vb33gy  = 3'd5;

  wire [psxtg_0xr2lkj4049fu-1:0] bv6l6emrtk2jtqlt;
  wire [psxtg_0xr2lkj4049fu-1:0] kjlcok4umxxx55_7a;
  wire z34lqkyodsolv0ogf;

  wire [psxtg_0xr2lkj4049fu-1:0] u99tnldu986760c5;
  wire [psxtg_0xr2lkj4049fu-1:0] nb3914w6z5nmnlsmou;
  wire [psxtg_0xr2lkj4049fu-1:0] y5ramxcxkrqsz12gk;
  wire [psxtg_0xr2lkj4049fu-1:0] ry8d7x33kgj4n14g;
  wire [psxtg_0xr2lkj4049fu-1:0] bmoq17r3wc66qf26;
  wire [psxtg_0xr2lkj4049fu-1:0] xhsqvfdidt5pi73vflj;
  wire wfoen161d4r42bkqp34lj;
  wire ar7ss7g0h7o9d58_adekeyg;
  wire hln5byq3t_zxwy8c51dq;
  wire kw11y7fxacdlitoe4r8m;
  wire jen_u9yotkl41mh0z6i_;
  wire bx88i6bwlcax77b86ju78j9;

  wire bh0_09jdv_nabkpizd8n = ze2bfnigu62i9937pcxnjc & c86b14qr2qo45_qw2ns;


  assign mz_exhb6gtbcmmad884 = (kjlcok4umxxx55_7a == uk1oi33ntqrycsuxu);
  wire bmvfssucdy0r3n27ax8n0lk   = (kjlcok4umxxx55_7a == dcmmvnhb4tmumn60lcp4);
  wire vcmhu_hc1hyry96oi3iy   = (kjlcok4umxxx55_7a == dsix6p9ipz7r85mja3fr);
  wire pg1c74tginny3v957a   = (kjlcok4umxxx55_7a == ulyzdpaocwknytnebndi);
  wire soksz54m8dbj9im9wsptt   = (kjlcok4umxxx55_7a == ojf5u64xjqjjuk3p);
  assign rs9cr43eb36gq815zlxyw = (kjlcok4umxxx55_7a == f6n2huuf8s7hdk3vb33gy);



  assign wfoen161d4r42bkqp34lj = mz_exhb6gtbcmmad884 & s9hgy6syn2arl9fxs8kb0;
  assign u99tnldu986760c5      = vldo6rbn ? dcmmvnhb4tmumn60lcp4 : f6n2huuf8s7hdk3vb33gy;



  assign ar7ss7g0h7o9d58_adekeyg  = bmvfssucdy0r3n27ax8n0lk & bh0_09jdv_nabkpizd8n;
  assign nb3914w6z5nmnlsmou     = dsix6p9ipz7r85mja3fr; 



  wire pcfm3_o_60ze1zpucjl;
  assign hln5byq3t_zxwy8c51dq = vcmhu_hc1hyry96oi3iy & bh0_09jdv_nabkpizd8n;
  assign y5ramxcxkrqsz12gk      = pcfm3_o_60ze1zpucjl ? (

                                         ulyzdpaocwknytnebndi 
                                     ): dsix6p9ipz7r85mja3fr;



  assign kw11y7fxacdlitoe4r8m = pg1c74tginny3v957a;
  assign ry8d7x33kgj4n14g      = ojf5u64xjqjjuk3p;



  assign jen_u9yotkl41mh0z6i_ = soksz54m8dbj9im9wsptt & jetszpnn_3n3x0k4d;
  assign bmoq17r3wc66qf26      = uk1oi33ntqrycsuxu;



  assign bx88i6bwlcax77b86ju78j9 = rs9cr43eb36gq815zlxyw & jetszpnn_3n3x0k4d; 
  assign xhsqvfdidt5pi73vflj      = uk1oi33ntqrycsuxu;


  assign z34lqkyodsolv0ogf = 
            bx88i6bwlcax77b86ju78j9 | 
            wfoen161d4r42bkqp34lj | ar7ss7g0h7o9d58_adekeyg |
            hln5byq3t_zxwy8c51dq | kw11y7fxacdlitoe4r8m | jen_u9yotkl41mh0z6i_;


  assign bv6l6emrtk2jtqlt = 
              ({psxtg_0xr2lkj4049fu{wfoen161d4r42bkqp34lj}} & u99tnldu986760c5)
            | ({psxtg_0xr2lkj4049fu{ar7ss7g0h7o9d58_adekeyg}} & nb3914w6z5nmnlsmou)
            | ({psxtg_0xr2lkj4049fu{hln5byq3t_zxwy8c51dq}} & y5ramxcxkrqsz12gk)
            | ({psxtg_0xr2lkj4049fu{kw11y7fxacdlitoe4r8m}} & ry8d7x33kgj4n14g)
            | ({psxtg_0xr2lkj4049fu{jen_u9yotkl41mh0z6i_}} & bmoq17r3wc66qf26)
            | ({psxtg_0xr2lkj4049fu{bx88i6bwlcax77b86ju78j9}} & xhsqvfdidt5pi73vflj)
              ;

  ux607_gnrl_dfflr #(psxtg_0xr2lkj4049fu) q6b8flgtd20mns11fqijy0 (z34lqkyodsolv0ogf, bv6l6emrtk2jtqlt, kjlcok4umxxx55_7a, gf33atgy, ru_wi);


  wire zqa26f3l044pht447ti8x_r8rmh = bh0_09jdv_nabkpizd8n & pcfm3_o_60ze1zpucjl & (~rs9cr43eb36gq815zlxyw);


  wire rxdv_strr1zu5v3089;

  wire azquruhbc8yno4oiyxp3 = bh0_09jdv_nabkpizd8n & dm5b92mx0redfbuhs1u3d;

  wire w8g9twm7ppcb3d_8vph7tuhb = (rxdv_strr1zu5v3089 & zqa26f3l044pht447ti8x_r8rmh & (~rs9cr43eb36gq815zlxyw)) | (rs9cr43eb36gq815zlxyw) | jen_u9yotkl41mh0z6i_;
  wire jagkgo9nth3fi4klq_oq = azquruhbc8yno4oiyxp3 |   w8g9twm7ppcb3d_8vph7tuhb;
  wire y028n58upnp4w9hwyjwqs = azquruhbc8yno4oiyxp3 & (~w8g9twm7ppcb3d_8vph7tuhb);
  ux607_gnrl_dfflr #(1) d0cwbbaw7vf012nya43lz1ze4y (jagkgo9nth3fi4klq_oq, y028n58upnp4w9hwyjwqs, rxdv_strr1zu5v3089, gf33atgy, ru_wi);


  wire s78ikg9hquflzdsoa50 = rxdv_strr1zu5v3089 | dm5b92mx0redfbuhs1u3d;

  localparam dxx8rixryrt7szii2ccmya6wpv0siby6 = (4-1);


  wire [2-1:0] kwbmlmwj_ec;

  wire d2jsegrkoa154kuy = s9hgy6syn2arl9fxs8kb0;

  wire bxc0qc1hr_cb1a4x1zadth = (kwbmlmwj_ec == 2'b0);
  wire nlfdn3rz3118m7vvwo = (kwbmlmwj_ec == dxx8rixryrt7szii2ccmya6wpv0siby6[2-1:0]);
  wire jxpj6_9tx5iktrgs = (s9hgy6syn2arl9fxs8kb0 & nlfdn3rz3118m7vvwo & (~s2cclwenb)) | (s9hgy6syn2arl9fxs8kb0 & s2cclwenb);
  wire v0t2k69nbehh = d2jsegrkoa154kuy | jxpj6_9tx5iktrgs;
  wire [2-1:0] ox18q467wzh8vsuj = 
                                   jxpj6_9tx5iktrgs ? {2{1'b0}}
                                 : d2jsegrkoa154kuy ? (kwbmlmwj_ec + {{2-1{1'b0}},1'b1})
                                 : kwbmlmwj_ec;

  ux607_gnrl_dfflr #(2) opyi12br8u9_35k_ni (v0t2k69nbehh, ox18q467wzh8vsuj, kwbmlmwj_ec, gf33atgy, ru_wi);



  wire srsur0x8i_d2khxf83xzyc0;
  
  wire lgt21324tq1wwwu167_ec2;
      
  wire wab0wlezupg8xip1e_f3y4 = zqa26f3l044pht447ti8x_r8rmh;
  wire cmyozk4r25iwfy7f3ed5kq = ~y7_io5z_hoy7o_sd1g7q[1];
  ux607_gnrl_dfflr #(1) x9tkawrtfc58mp1fsvb32 (wab0wlezupg8xip1e_f3y4, cmyozk4r25iwfy7f3ed5kq, lgt21324tq1wwwu167_ec2, gf33atgy, ru_wi);


      
  wire rvqd_f3xavh2sant2_yfgtyzk =   wfoen161d4r42bkqp34lj
                               & (~vcalsdo6q)       
                               ;
       
  
  
  
  
  wire yohv8w1bq84fhs5y__rl62uil = (~xvnxfgnlx05) ? 1'b0 : (~h6yap55ubdbc2) ? 1'b1 : smqoz2oj8ww5don ? 1'b1 : dh_clbn0o20fgf4 ? 1'b0 : lgt21324tq1wwwu167_ec2; 
  ux607_gnrl_dfflr #(1) tigdtt8h6mfvro2f41idum07j5 (rvqd_f3xavh2sant2_yfgtyzk, yohv8w1bq84fhs5y__rl62uil, srsur0x8i_d2khxf83xzyc0, gf33atgy, ru_wi);
  assign y7_io5z_hoy7o_sd1g7q = {srsur0x8i_d2khxf83xzyc0,~srsur0x8i_d2khxf83xzyc0};








  
  
  
  
  



      
  wire lrfp7w5wbqmdbgg =   jetszpnn_3n3x0k4d & (~lkjqs6kiuyj) 
                    & (~vcalsdo6q)    
                    & (~y75xeozj0wna88fi2) 
                    & (~(~t3tudcq0j & aknbc4862andzqg1530a & ylm6yo9kkk2s745bw1ay)) 
                    & (~ub__mzukp2wlfwg)  
                    & (~peo2y31x_joi)    
                    ; 
      
  wire i9bwopch0ryfz = afyql3m7n_e_ &        
                    (  vldo6rbn 
                     | rofqn5vmqgj3
                     | vcalsdo6q      
                     | y75xeozj0wna88fi2   
                     | (~t3tudcq0j & aknbc4862andzqg1530a & ylm6yo9kkk2s745bw1ay)   
                     | ub__mzukp2wlfwg 
                     | peo2y31x_joi      
                    );
  wire ybr_23ro0z = lrfp7w5wbqmdbgg |   i9bwopch0ryfz;
  wire f7jj894j70g5aoz = lrfp7w5wbqmdbgg | (~i9bwopch0ryfz);
  ux607_gnrl_dfflr #(1) odr241tuo1wb1bf5w (ybr_23ro0z, f7jj894j70g5aoz, afyql3m7n_e_, gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1) cf9xoiepa_wr5eja06whun (lrfp7w5wbqmdbgg, ffd_fx0uggmz_c, bvs0w3jafe5oum96j06, gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1) pth9eymd51tgse0c4h8b (lrfp7w5wbqmdbgg, r2zjd7aqmv0bk_c4, swrbe70hp3wsvkt04, gf33atgy, ru_wi);





  wire tqiycgs52p5ubxsuyib_v1zt7;


  wire xb8j0rrc_88sw9m1_7ximu1sj = (vldo6rbn | s2cclwenb)
                               & (~(ub__mzukp2wlfwg & b0nb3z34fjl))  
                               ;

  wire ydasmvx5h2ezeqd8nzjocww = tqiycgs52p5ubxsuyib_v1zt7 & jxpj6_9tx5iktrgs;
  wire u27qjkb5zqe12szsltsn84e = xb8j0rrc_88sw9m1_7ximu1sj |   ydasmvx5h2ezeqd8nzjocww;
  wire oy67t8p1b1as7_r4qp4hek3jt = xb8j0rrc_88sw9m1_7ximu1sj & (~ydasmvx5h2ezeqd8nzjocww);
  ux607_gnrl_dfflr #(1) v3tueeign88vdxdo7qvw12ytrgj (u27qjkb5zqe12szsltsn84e, oy67t8p1b1as7_r4qp4hek3jt, tqiycgs52p5ubxsuyib_v1zt7, gf33atgy, ru_wi);

  assign  rinamilgle00i5xmx_vt = tqiycgs52p5ubxsuyib_v1zt7; 
  wire  [64-1:0] wtk3umqu7dl52syp47vyeq99nc = {nf7a14kdh46q_gb4d27t5o,kwbmlmwj_ec,{5-2{1'b0}}};   
  assign  z64bwdr23steb7s9y9j  = s2cclwenb ? axng6pw6x_ngow1o7_7e[64-1:0] : wtk3umqu7dl52syp47vyeq99nc[64-1:0];
  assign  cneu8a119tg3vmie6zr2h_  = z5oodn6lsltcchb6;
  assign  jw2dzv9gi7gygudyqql6fz  = w_45r8lsw7umpt;
  assign  ybcilssdlw64sqj1jf2uuk  = mu_grj5_po0a4ek;
  assign  bg1spy6_v2kbo75pz1d6  = 1'b1;
  assign  b7aet1zp_fcfxn8h7rw0u1 = s2cclwenb ? 3'b0 : 3'b001; 
  wire  q7k1vzcndghghxtpbf = bxc0qc1hr_cb1a4x1zadth;
  wire  cu9wchz0hcex50o2m_yx   = nlfdn3rz3118m7vvwo;
  assign  t3szwnvfo2nj3wk6r5kvt = s2cclwenb ? 2'b0 : {cu9wchz0hcex50o2m_yx,q7k1vzcndghghxtpbf};

  assign  o_7kpry6inkqpqi1bf1nd  = ik4xc_1hh4vb;

  assign bngbyv57e7juc0vkk2y8i = 2'b11;
  assign znotwr53pu47f5m1agm = vcalsdo6q; 

  assign  c86b14qr2qo45_qw2ns = 1'b1;





  wire [2-1:0] m8e4y5p5zfei0w;

  wire rzjjndlw_np7otl63 = bh0_09jdv_nabkpizd8n;

  wire xp_8ug3xaxvs1hzjo4ime = (m8e4y5p5zfei0w == 2'b0);
  assign pcfm3_o_60ze1zpucjl = (m8e4y5p5zfei0w == dxx8rixryrt7szii2ccmya6wpv0siby6[2-1:0]);
  wire xzheht9iavqj32dq7zx = bh0_09jdv_nabkpizd8n & (pcfm3_o_60ze1zpucjl | rs9cr43eb36gq815zlxyw);
  wire ddht2k_7yytr_fa5yogp = rzjjndlw_np7otl63 | xzheht9iavqj32dq7zx;
  wire [2-1:0] csy24t9fh7gacp9f = 
                                   xzheht9iavqj32dq7zx ? {2{1'b0}}
                                 : rzjjndlw_np7otl63 ? (m8e4y5p5zfei0w + {{2-1{1'b0}},1'b1})
                                 : m8e4y5p5zfei0w;

  ux607_gnrl_dfflr #(2) ui0nyss5vsvizbzfh0s (ddht2k_7yytr_fa5yogp, csy24t9fh7gacp9f, m8e4y5p5zfei0w, gf33atgy, ru_wi);


  
  

  wire [7-1:0] oidscd0mdfv76z6y5i2;
  wire [54-1:0] t3xigewvakukwi5op5n;

  wire cyr03zozo15rbmqfsz = zqa26f3l044pht447ti8x_r8rmh;
  assign oidscd0mdfv76z6y5i2 =  pkmbkt_zq0yhlemrgi;
  wire smyk8ej9_zno4ljmfy31z27 = (~jy8uskaamz5hsuj8mmvvc) & (~s78ikg9hquflzdsoa50); 
  assign t3xigewvakukwi5op5n = {smyk8ej9_zno4ljmfy31z27,(~s78ikg9hquflzdsoa50),jcbv86t6ccbny9um2sm};

  wire   op8ambdz_hjfyg81uq = cyr03zozo15rbmqfsz;
  assign gsf_5l61c1nvvp_  = 1'b1;
  assign akg6apmoz04bjkagrh = oidscd0mdfv76z6y5i2;
  assign fxu0h92n3g4evsus = t3xigewvakukwi5op5n;
  
  
  

  assign l7sauvhwo7orvwq0tz6tql = op8ambdz_hjfyg81uq & (y7_io5z_hoy7o_sd1g7q[0]);
  assign d3j_g8wp81xd22uqe66u = op8ambdz_hjfyg81uq & (y7_io5z_hoy7o_sd1g7q[1]);
  

  wire [64-1:0] fdmi7fg9f6ept_m29;
  wire [9-1:0] l01f_bx4m_wbuk6qjo;

  wire n82reuy_65gf4spkcsb;

  assign l01f_bx4m_wbuk6qjo = {pkmbkt_zq0yhlemrgi,m8e4y5p5zfei0w[2-1:0]};
  assign n82reuy_65gf4spkcsb = bh0_09jdv_nabkpizd8n
                            & (~rs9cr43eb36gq815zlxyw)
                            ;
  assign fdmi7fg9f6ept_m29 = c3vtv1izxu7rm5646jsmmke;

  wire [9-1:0] a8hig8_6g8dji5gkavyf5x9;
  wire [64-1:0] ql3qkkln3havus2mn;

  wire s0czoufc7wwoykscl3ay = pg1c74tginny3v957a;
  assign a8hig8_6g8dji5gkavyf5x9 = {pkmbkt_zq0yhlemrgi,m603xpg5m7bwf6h1d[5-1:3]};
  assign ql3qkkln3havus2mn = 64'b0;

  wire   cfi2cflhc_lax1a0 = s0czoufc7wwoykscl3ay | n82reuy_65gf4spkcsb;
  assign r5947sq0alkh4q  = ~s0czoufc7wwoykscl3ay;  
  assign g7c1415q8kv_x6ed0 = s0czoufc7wwoykscl3ay ? a8hig8_6g8dji5gkavyf5x9 : l01f_bx4m_wbuk6qjo;
  assign dkn8bvcvpdmu34 = fdmi7fg9f6ept_m29;
  

  assign rj69sa3044rb1cz6lvd6 = cfi2cflhc_lax1a0 & (y7_io5z_hoy7o_sd1g7q[0]);
  assign atpyq4kwa38ur5a1v4jxl = cfi2cflhc_lax1a0 & (y7_io5z_hoy7o_sd1g7q[1]);











  assign h7f6k_ims_9p3 = 

      (gdc31z_ah0g & dd8s8azwnmm78) ? 64'b0 :

      (s2cclwenb & dd8s8azwnmm78) ? 64'b0 :
      (gjkof2a42or0w) ? c3vtv1izxu7rm5646jsmmke :
      ikf61_i17b0iv;

  assign b24yx4ictsbkcpj =  soksz54m8dbj9im9wsptt;


  localparam s3xvyho = 1
                    +1
                    +1
                    ;
  localparam ldebclccia0aslswkob = 64 + s3xvyho +1;
  assign iaaolhc_afh_9est07sqv = 1'b1;
  wire ygjpyr2srt2fpb7a;
  wire k0p07wax7i8qs4irfw = klkflmsyyf5w7ar;

  assign wy36iirxspfw56864 = ygjpyr2srt2fpb7a;
  wire [s3xvyho-1:0] iwxu78sftoab_xrp = { sxxoah7zbvh8noti 
                                  ,wgls7kw8r0vwnfoaa5 
                                  ,ub__mzukp2wlfwg 
                                  };

  wire [ldebclccia0aslswkob-1:0] r194g36kplm5e5jwt = { h7f6k_ims_9p3
                                              ,lkjqs6kiuyj 
                                              ,iwxu78sftoab_xrp };

  wire [ldebclccia0aslswkob-1:0] d7jq9fe2dpeqo396iig;
  wire [64-1:0] k2vp4nzypxpjqeoddj5a;
  wire u6w9b_jfa7l3hw7mrgi;
  wire [s3xvyho-1:0] q1oyh77hy0fh3o_gc7l4p;

  assign {  k2vp4nzypxpjqeoddj5a, 
            u6w9b_jfa7l3hw7mrgi,
            q1oyh77hy0fh3o_gc7l4p} = d7jq9fe2dpeqo396iig;





 ux607_gnrl_pipe_stage # (
  .CUT_READY(0),
  .DP(1),
  .DW(ldebclccia0aslswkob)
 ) qoccbsp276dce0kljty6520ey1 (
   .i_vld(k0p07wax7i8qs4irfw),
   .i_rdy(ygjpyr2srt2fpb7a), 
   .i_dat(r194g36kplm5e5jwt),
   .o_vld(zs89k7qgupd1xlvx63l2r), 
   .o_rdy(iaaolhc_afh_9est07sqv), 
   .o_dat(d7jq9fe2dpeqo396iig),
 
   .clk  (gf33atgy  ),
   .rst_n(ru_wi)  
  );

  wire lgp85z8w1yr70nji5eu7s;

  assign {
            ba1ucnyekcm68i9wuqwmn,
            bpyef3a0dnkkyqdpymy,
            wv442dsr_nxty0qoldk7qmqg
            ,b2loifdzo9b2smec06r0t
            ,lgp85z8w1yr70nji5eu7s
                                    } = d7jq9fe2dpeqo396iig; 

  assign phzkntckzzbndu4wevf1o6 =   zs89k7qgupd1xlvx63l2r
                                & (~lgp85z8w1yr70nji5eu7s)  
                                ; 

  wire p8i6r5vz69gazn0pr;
  wire cxou18bigclxcjkbnjml = op8ambdz_hjfyg81uq;  
  wire rzpb_jtv4nmn84vmfqq = s78ikg9hquflzdsoa50;
  ux607_gnrl_dfflr #(1) x3j5r33aste6_n1_oz28_ (cxou18bigclxcjkbnjml, rzpb_jtv4nmn84vmfqq, p8i6r5vz69gazn0pr, gf33atgy, ru_wi);

  assign vh2j7b0kt7n2s59 = p8i6r5vz69gazn0pr;

  assign tx07brh7_ullbwlubonaqwg2 = 1'b0;






  

  
  wire vqky7j0dc35ibhbc5wg = cyjoizk175tz59s73g1; 
  assign v94hbvyskjuea4n7wsw4d = pkmbkt_zq0yhlemrgi; 
  assign wfvfwnnky0p7at5zp07vtk = jcbv86t6ccbny9um2sm; 
  ux607_gnrl_dfflr #(                      1)  gcz4yve1rlu_vw5611          (vqky7j0dc35ibhbc5wg, gdc31z_ah0g,           egsj_v4pl_4,           gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(                      1)  ternu54dvn4sosl1ye         (vqky7j0dc35ibhbc5wg, vldo6rbn,          wo2xz_n9y7nkzka,          gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(                      1)  efjs13ek0oj8afashz90       (vqky7j0dc35ibhbc5wg, vcalsdo6q,        vkhotkpp9yeqfbubp,        gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(                      1)  yyvt0w6igryqos5r97hfv      (vqky7j0dc35ibhbc5wg, dd8s8azwnmm78,       mhd_d53mz4u2o78ojq,       gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(                      1)  bfj_uo4nyv0a8hbbtbpmofmb     (vqky7j0dc35ibhbc5wg, b0nb3z34fjl,      tqd1xxmvx9svwxcdh32,      gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(                      1)  k9hlwsjcmz3xs3b3un2cr7     (vqky7j0dc35ibhbc5wg, u7ja7msr33bxl,      fdjtu3kedjy4crxuyi,      gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(                      1)  k1rbzcuqcppq_ud_1z081gn       (vqky7j0dc35ibhbc5wg, b293miy3ig80jz,        nd_hcfia24v6mp0zx,        gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(                      1)  x9nt12zywu39zp1bogffrc_3z  (vqky7j0dc35ibhbc5wg, l_razgaao587019p,   z1gnqpih0tzo73j7opinl,   gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(                      1)  ub4nbhqwq6mtg6rwr4en2_x8r       (vqky7j0dc35ibhbc5wg, yz14ncxfv0,        va1c1blelsdo93uz,        gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(                      1)  rfwuhyd7j4kd1pbp1r7rfg3kye12  (vqky7j0dc35ibhbc5wg, iq0t6kp6qfri0qe61w,   cwxkjxgleg8vuggc_nh2xt8c,   gf33atgy, ru_wi);



  
  
  
  

  assign peo2y31x_joi = 1'b0; 
  assign jm9hjt3oqbob590sdfe = 7'b0;
  assign wb4vwdrejqmlx7swh7a_0b  = 54'b0;

   assign rjy1mb7tnflt7ea = 1'b0;  
   assign hxztlrjkqickn6urw = 1'b0;

  
  assign zug6nwomkc29qfxbzdpocn = v94hbvyskjuea4n7wsw4d        ; 
  assign d9hprjtpa534yd5p17wt33b9h = wfvfwnnky0p7at5zp07vtk        ; 
  assign rng0m4_qo_00          = egsj_v4pl_4            ;
  assign zbshs61j683bajzde         = wo2xz_n9y7nkzka           ;
  assign zej0zy3isij_80da       = vkhotkpp9yeqfbubp         ;
  assign tr3x6j926x74p00e      = mhd_d53mz4u2o78ojq        ;
  assign luex4fm_4zh4bo58e1b4l     = tqd1xxmvx9svwxcdh32       ;
  assign wtbx6tgxz2r4ze7xt     = fdjtu3kedjy4crxuyi       ;
  assign c3pqxq1ukkc352nk       = nd_hcfia24v6mp0zx         ;
  assign kw97mqedpw8dwl56q6_zx5  = z1gnqpih0tzo73j7opinl    ;
  assign hkvmg02232a2c9zb       = va1c1blelsdo93uz         ;
  assign duy9wppkj4is5xqmehcjyu6  = cwxkjxgleg8vuggc_nh2xt8c    ;

  
  assign ig7796duzb8wqodp = ~wz_if_2q_23jhl2;


endmodule


















module pgil4p_zywsz2lytb (
  input  s7eq8f6z1uyi2in,

  input  hab9b2zcdgrlbutx5,
  input  uub2rxsi1qvmca,
  input  p_xqcszydp2j5d821j,
  input  hwpkcsh2atrq  ,
  input  v3e6l1k7eo9k3 ,
  input  hxrmt706n071lic0f7,
  input  [4*8-1:0] horqgj1y_r_5aplro,
  output [4*8-1:0] iqaziwvuq5463k3, 
  output [4*8-1:0] hs5w0q7r19myj9eezz, 
  output [7:0] rhrr146mr7lt9h,
  output [7:0] io1uhjqtpgin_,
  output [2:0] gohm8ye7tw32so,
  input  [2:0] d0q_15ed0hmwqygja,
  input  vp5_qftup10p3v7_jw8,
  input  [7:0] q1zci4ybfd7ftj8qxl2,
  input  v7rzl8qveorn2jg6659m69,
  input  v_k8ohy_e2e9vlp6az04,
  input [2-1:0] gtvau5cygdmb10dr_makqf,
  input  [9-1:0] p54semfzu2zyfb,
  output [9-1:0] m2_t547jr8crh6jgy4c,
  input  [64-1:0] y_vw514j6xmphhfhc,



  input  [64-1:0] pz6cvxcjpgv,
  input  [64-1:0] haezj87elp_,
  input  [64-1:0] z1p1oekb0pd,
  input  [64-1:0] js_7wqgsstbnxcjr29, 
  input  [64-1:0] eajem3pnezl,
  input  vmfcanu2o,
  input  v5uyqoe,
  input  agjzm78wm,


  input lln3b7iev7jpvogh964ro_9bc_3y,
  input q97rqfy8n7ixfm2a5wev4nd5sylpcq3j,
  input hujgg6hjnhtbspbkekuz5_u,
  input v3pnt81kfrgbaanm1mhh51w,
  input [64-1:0] i08eq60d_snxeq8si_ezod,

  input y8wz7aud_fd6dfiakjtx2i0g,
  input dgnjyd9xs8efyxm0tdlsvfq4eop,
  input a3xib90kwk4_hm1,
  input nfzexr8q9g893gi,
  input [64-1:0] opkkwp3eg8g3448t,


  input  bnjz04i86zhxx6,
  input  qpotfvbjdo6qtsy1,
  input  ua8gydukonfboz,
  input  vkfewi0rkx,
  input  iq5y0wse0y2,
  input  [64-1:0] ueimo2s8tf29_f,
  input  jzcjplpewzvpowh,

  input  jvcw7os6duv6_6,
  input  k0q5465tih57fj,
  input  sfgacjvxnybsqrx_,
  input  z9lf1gw3iz9e,
  input  m_pst8fyu48q6i4,
  input  [64-1:0] xl0lr2g890tskf74yu8,
  input  jvt4ma57k62vz,


  output jrkjeqdo7hhdsjna,  
  output cmvxg4cmkkrry,  
  output r9arh0s0wxc_0,
  output vgno0maw8a,
  output gj95joew8j70jj4,  
  output [64-1:0] cs_6ujj3b74,
  output v0u85q8u16_pwgz7h17cl4,
  output yov0d70301nwd4bbqbyv,
  output [2-1:0] dwz7mnj7ox5,
  output g1iutrfs,




  input  tbs7se44h1m47t,
  input  ct8_j4rs_zvw4xjl_ncf,
  input  ovuaqnjxywro47yxbn20wg3m,
  output v4gayo0h8l6na,
  output [64-1:0] nmy2nw74r7gg,

  input  gf33atgy,
  input  ru_wi
);

localparam n8duywjqdzotwzmrk9_pvp = 4 - 1;





assign r9arh0s0wxc_0 = 1'b1;
assign vgno0maw8a = ~jrkjeqdo7hhdsjna;
wire rgktjw6f9n9zt88ljy = (iq5y0wse0y2 | bnjz04i86zhxx6);
wire qe_4occxaraqc2ts = (m_pst8fyu48q6i4 | jvcw7os6duv6_6);
wire vgaethe0agg = (iq5y0wse0y2 | bnjz04i86zhxx6 | qpotfvbjdo6qtsy1);
wire zqoqj6wzo4ba = (m_pst8fyu48q6i4 | jvcw7os6duv6_6 | k0q5465tih57fj);
wire ld01d40_n3 = vgaethe0agg ? 1'b1 : zqoqj6wzo4ba;
wire k3epsun0zhok7c = bnjz04i86zhxx6 | qpotfvbjdo6qtsy1;
wire w5ijrcxx7v_ = jvcw7os6duv6_6 | k0q5465tih57fj;
wire c52s23xseom3eeuj7rv1p6c = hab9b2zcdgrlbutx5 & (~ct8_j4rs_zvw4xjl_ncf)
                            & (~ovuaqnjxywro47yxbn20wg3m)
                            ;
wire cd3xfhf_7i5g014tqu9 = ld01d40_n3 & c52s23xseom3eeuj7rv1p6c;
wire v13larpmyvauxb09yna = (ua8gydukonfboz & (~vkfewi0rkx));
wire embwyxsrpkcrh8lpx5n = (~jrkjeqdo7hhdsjna) & (sfgacjvxnybsqrx_ & (~z9lf1gw3iz9e));
wire a1ga0w9x_xs14kysw = (~ua8gydukonfboz) & vkfewi0rkx;
wire vyyjlm5cyybbpwqm = (~jrkjeqdo7hhdsjna) & (~sfgacjvxnybsqrx_) & z9lf1gw3iz9e;
wire ywsaub3r999h9pyn = v13larpmyvauxb09yna | embwyxsrpkcrh8lpx5n; 
wire r12cr5tap6v  = a1ga0w9x_xs14kysw  | vyyjlm5cyybbpwqm; 

wire [64-1:0] xe0fwqp049g43;
wire qvjzfqc6tqntswnail = cd3xfhf_7i5g014tqu9 & ywsaub3r999h9pyn;
wire wqior_n5rxvoa3677tk = cd3xfhf_7i5g014tqu9 & r12cr5tap6v;
wire [64-1:0] cfl5vsneikbk178yg = v13larpmyvauxb09yna ? haezj87elp_ : eajem3pnezl;

wire [4-1:0] hz7o7599ynpzl85u_;
wire [4-1:0] uzf98ssxae_2yyluij2_;
wire [64*4-1:0] b9nie3as2itq9uwhb;
wire [4-1:0] ezszbkw3zin7538qds1fl;
wire [64*4-1:0] pucwp8ukjgqsm8k2pk71;
wire [4-1:0] d5w1v6m8iup9wx4yilq_tfw1wu;
wire [4-1:0] mwmqribws2g9iv7qhjdvg1fmff;
wire [64*4-1:0] qguwwpo1_cvf5xrfx51bfwx;
wire [64*4-1:0] ip7o8y9uhp6ghrk;
wire [4-1:0] ko5r9koxflyi2;
wire [4-1:0] nz37pr5kdbvvivl;

wire pwdhc0a__bijmzio7gex_9drs8as9_tcm75hz;
wire aj_vxfegy_shy6wejfx7h030ac;
wire nzr8b08z878kkyjporqv8l4z9tesua1_tm;
wire zxvy4k9s3wmbt4828om4 = dgnjyd9xs8efyxm0tdlsvfq4eop & aj_vxfegy_shy6wejfx7h030ac;
wire vlg_ydu5zngc34fl0zi1n94g3w = (q97rqfy8n7ixfm2a5wev4nd5sylpcq3j & (~dgnjyd9xs8efyxm0tdlsvfq4eop)) & pwdhc0a__bijmzio7gex_9drs8as9_tcm75hz;
wire n85msjeqs4hcws4eadp7i =  zxvy4k9s3wmbt4828om4 | vlg_ydu5zngc34fl0zi1n94g3w; 

wire ipg89cfwypzx93hyc2c9n  = dgnjyd9xs8efyxm0tdlsvfq4eop & nzr8b08z878kkyjporqv8l4z9tesua1_tm;
wire j3hvi4xu8v_1e184xsbn2yg = y8wz7aud_fd6dfiakjtx2i0g & a3xib90kwk4_hm1;
wire gs0ylhknmfa43yp5pdreui9iga3o8 = lln3b7iev7jpvogh964ro_9bc_3y & hujgg6hjnhtbspbkekuz5_u;

genvar i;
generate
    for (i=0; i<4; i=i+1) begin:uc80ngop2mcb
assign b9nie3as2itq9uwhb[64*(i+1)-1:64*i] = zxvy4k9s3wmbt4828om4 ? 
                                                                (
                                                                    (j3hvi4xu8v_1e184xsbn2yg & ko5r9koxflyi2[i]) ?
                                                                                          opkkwp3eg8g3448t : 
                                                                                          ip7o8y9uhp6ghrk[64*(i+1)-1:64*i]
                                                                )
                                                                : (
                                                                    (gs0ylhknmfa43yp5pdreui9iga3o8 & ezszbkw3zin7538qds1fl[i]) ? 
                                                                                           i08eq60d_snxeq8si_ezod : 
                                                                                           pucwp8ukjgqsm8k2pk71[64*(i+1)-1:64*i]
                                                                  );

assign qguwwpo1_cvf5xrfx51bfwx[64*(i+1)-1:64*i] = (
                                                                       y8wz7aud_fd6dfiakjtx2i0g & 
                                                                       a3xib90kwk4_hm1 &
                                                                       ko5r9koxflyi2[i]
                                                                                     ) ?  opkkwp3eg8g3448t
                                                                                       :  ip7o8y9uhp6ghrk[64*(i+1)-1:64*i];  
    end
endgenerate

assign uzf98ssxae_2yyluij2_ =  zxvy4k9s3wmbt4828om4 ? (y8wz7aud_fd6dfiakjtx2i0g ? nz37pr5kdbvvivl 
                                                                          : ko5r9koxflyi2
                                                                          )
                                                 : (lln3b7iev7jpvogh964ro_9bc_3y ? d5w1v6m8iup9wx4yilq_tfw1wu 
                                                                                : ezszbkw3zin7538qds1fl
                                                                                )
                                                 ;
assign mwmqribws2g9iv7qhjdvg1fmff = y8wz7aud_fd6dfiakjtx2i0g ? nz37pr5kdbvvivl : ko5r9koxflyi2;

wire [5:0] av1knj27e6usz4u73;
wire [5:0] lrlesb91b476d44aqsj9ij8;
wire [5:0] acw0h9s07558hb5vs3;
wire [5:0] wcwsqyyganwv3c0akygn;
wire [5:0] nk19sm_cd4kwt126vaoe0u4rl;
wire [5:0] t8dr6tuoip7dpev2t5;
wire [5:0] sk27p61gpcedx_dx552 = av1knj27e6usz4u73 + 1'b1; 
wire [5:0] f7ty9qo488rjon9u9aqc3c = lrlesb91b476d44aqsj9ij8 + 1'b1; 
wire [5:0] ibzncuj29jn0t_a533 = acw0h9s07558hb5vs3 + 1'b1; 

assign wcwsqyyganwv3c0akygn =
                                (y8wz7aud_fd6dfiakjtx2i0g & a3xib90kwk4_hm1) ? t8dr6tuoip7dpev2t5 : 
                                                   dgnjyd9xs8efyxm0tdlsvfq4eop ? acw0h9s07558hb5vs3 : 
                    (lln3b7iev7jpvogh964ro_9bc_3y & hujgg6hjnhtbspbkekuz5_u) ? f7ty9qo488rjon9u9aqc3c : 
                                             q97rqfy8n7ixfm2a5wev4nd5sylpcq3j ? lrlesb91b476d44aqsj9ij8 : 
                                                                            sk27p61gpcedx_dx552;

wire ptxajgmm3swyp9ye = qvjzfqc6tqntswnail | q97rqfy8n7ixfm2a5wev4nd5sylpcq3j | dgnjyd9xs8efyxm0tdlsvfq4eop;
ux607_gnrl_dfflr #(6) asltng8nljtaq7bjwdeg3r8hxo(ptxajgmm3swyp9ye, wcwsqyyganwv3c0akygn, av1knj27e6usz4u73, gf33atgy, ru_wi);


assign nk19sm_cd4kwt126vaoe0u4rl =  (y8wz7aud_fd6dfiakjtx2i0g & a3xib90kwk4_hm1) ? t8dr6tuoip7dpev2t5 :
                                                   dgnjyd9xs8efyxm0tdlsvfq4eop ? acw0h9s07558hb5vs3 : 
                                                                            f7ty9qo488rjon9u9aqc3c;

wire uyms1h3s_s3u38su64o0vh_93 = hujgg6hjnhtbspbkekuz5_u | dgnjyd9xs8efyxm0tdlsvfq4eop;
ux607_gnrl_dfflr #(6) hytwxzqox21zvw1zm4md0ziazn7vt_kvhh2(uyms1h3s_s3u38su64o0vh_93, nk19sm_cd4kwt126vaoe0u4rl, lrlesb91b476d44aqsj9ij8, gf33atgy, ru_wi);


assign t8dr6tuoip7dpev2t5 =  ibzncuj29jn0t_a533;
wire eunxx9kthob_lj = a3xib90kwk4_hm1;
ux607_gnrl_dfflr #(6) brw3gv33083z85uzckuxw3dr9m(eunxx9kthob_lj, t8dr6tuoip7dpev2t5, acw0h9s07558hb5vs3, gf33atgy, ru_wi);

assign pwdhc0a__bijmzio7gex_9drs8as9_tcm75hz = (~(av1knj27e6usz4u73 == lrlesb91b476d44aqsj9ij8)) | (~(hz7o7599ynpzl85u_ == ezszbkw3zin7538qds1fl));
assign aj_vxfegy_shy6wejfx7h030ac       = (~(av1knj27e6usz4u73 == acw0h9s07558hb5vs3))       | (~(hz7o7599ynpzl85u_ == ko5r9koxflyi2));
assign nzr8b08z878kkyjporqv8l4z9tesua1_tm   = (~(lrlesb91b476d44aqsj9ij8 == acw0h9s07558hb5vs3))   | (~(ezszbkw3zin7538qds1fl == ko5r9koxflyi2));


p651q_8n0fzsut5za #(
    .onr7l(64),
    .mhdlk(4)
) l4k0j6krogkpjwzqvn23l21qd(
    .u22pp          (qvjzfqc6tqntswnail & s7eq8f6z1uyi2in),
    .irka0          (wqior_n5rxvoa3677tk & s7eq8f6z1uyi2in),
    .qbjvs30wtb          (cfl5vsneikbk178yg),
    .dqgck5s          (xe0fwqp049g43),
    .pc6rgvhuc_wry1q     (),
    .ks96miyn2gm4     (hz7o7599ynpzl85u_),
    .lexmfixlro03vle63iq (),
    .mhilu6fd3fe       (n85msjeqs4hcws4eadp7i & s7eq8f6z1uyi2in),
    .u60e_km0nn      (uzf98ssxae_2yyluij2_),
    .vjgphsh5tfo      (b9nie3as2itq9uwhb),
    .gf33atgy            (gf33atgy),
    .ru_wi          (ru_wi)
);

p651q_8n0fzsut5za #(
    .onr7l(64),
    .mhdlk(4)
) g2ozpw2q3rt7_2ss8qlzy(
    .u22pp          (hujgg6hjnhtbspbkekuz5_u & s7eq8f6z1uyi2in),
    .irka0          (v3pnt81kfrgbaanm1mhh51w & s7eq8f6z1uyi2in),
    .qbjvs30wtb          (i08eq60d_snxeq8si_ezod),
    .dqgck5s          (),
    .pc6rgvhuc_wry1q     (pucwp8ukjgqsm8k2pk71),
    .ks96miyn2gm4     (ezszbkw3zin7538qds1fl),
    .lexmfixlro03vle63iq (d5w1v6m8iup9wx4yilq_tfw1wu),
    .mhilu6fd3fe       (ipg89cfwypzx93hyc2c9n & s7eq8f6z1uyi2in),
    .u60e_km0nn      (mwmqribws2g9iv7qhjdvg1fmff),
    .vjgphsh5tfo      (qguwwpo1_cvf5xrfx51bfwx),
    .gf33atgy            (gf33atgy),
    .ru_wi          (ru_wi)
);

p651q_8n0fzsut5za #(
    .onr7l(64),
    .mhdlk(4)
) tk6q26mk3ftm14xnel1m(
    .u22pp          (a3xib90kwk4_hm1 & s7eq8f6z1uyi2in),
    .irka0          (nfzexr8q9g893gi & s7eq8f6z1uyi2in),
    .qbjvs30wtb          (opkkwp3eg8g3448t),
    .dqgck5s          (),
    .pc6rgvhuc_wry1q     (ip7o8y9uhp6ghrk),
    .ks96miyn2gm4     (ko5r9koxflyi2),
    .lexmfixlro03vle63iq (nz37pr5kdbvvivl),
    .mhilu6fd3fe       (1'b0),
    .u60e_km0nn      ({4{1'b0}}),
    .vjgphsh5tfo      ({64*4{1'b0}}),
    .gf33atgy            (gf33atgy),
    .ru_wi          (ru_wi)
);






wire [8-1:0] h1wgjzny5b2pljqb7ri;
wire [8-1:0] s1t3yek2syb4ot1hg0e_57qn9l;
wire                       l0ys343o73vqgkhn0dr0;
wire [8-1:0] a4rpu4iz_3odwqz;

wire wt74a9t1bcclq_xftx2 = v3e6l1k7eo9k3 & s7eq8f6z1uyi2in;
wire [8-1:0] qtzwuy827n9qcqls278 = {a4rpu4iz_3odwqz[8-2:0] ,hxrmt706n071lic0f7}; 

ux607_gnrl_dfflr #(8)  hc1h97jg2avrou(wt74a9t1bcclq_xftx2, qtzwuy827n9qcqls278, a4rpu4iz_3odwqz, gf33atgy, ru_wi);

assign l0ys343o73vqgkhn0dr0 = (wt74a9t1bcclq_xftx2 && hwpkcsh2atrq) || ((iq5y0wse0y2 | (vgno0maw8a & m_pst8fyu48q6i4)) && c52s23xseom3eeuj7rv1p6c);
assign s1t3yek2syb4ot1hg0e_57qn9l  = (hwpkcsh2atrq && wt74a9t1bcclq_xftx2) ? qtzwuy827n9qcqls278 : {h1wgjzny5b2pljqb7ri[8-2:0] ,gj95joew8j70jj4};

ux607_gnrl_dfflr #(8)  o4j1yb5u2uyaxt05_(l0ys343o73vqgkhn0dr0, s1t3yek2syb4ot1hg0e_57qn9l, h1wgjzny5b2pljqb7ri, gf33atgy, ru_wi);

wire  [8-1:0] i770uc76y777jzpfptztemfl;
wire  [8-1:0] q44ggnacf3_7f825zvirlm0owgd0;
wire  [1:0]                 jxcs4f4npbmy89g7pu0dwd680;
wire  [1:0]                 u5ls7fh44rneoy5rbkg0fjwarn;
wire                        xcuko0jmist_fz_ssr0gb4raa2has;
wire                        a1rgppa6mdbatjs4nhapuatya;
wire  [8-1:0] wcbtej7qnyi8h9j58z7vr134ulj;
wire  [8-1:0] s8o7h0k4g9_xuy00hgcfm4d0;
wire  [1:0]                 k4w5f9hywpks8xc21mnzjr;
wire  [1:0]                 pz4yvi8rtvnyll9wc_sl8aja8;
wire                        pizin3jqw9dy383sys4vfakj579;
wire                        eigqul3fdk4hzvxbs_b52aw63;
wire  [8-1:0] o2hausg38teon3_2f7g00su02;
wire  [8-1:0] ax7gdpn6yehlgk0b4bcdap_nvs2;
wire  [1:0]                 ppu_9xb8cwtqbebcovtfl6;
wire  [1:0]                 vtpt106_9th9gncs9klumvuhb8m;
wire                        f2k2cih_4nxcx3c0_a4s15af5d58;
wire                        mqzjxfzpvomdory6rh2y_v8l8wk;
wire  [8-1:0] m2kzu5wsbvwjfwip3zfvssodc;
wire  [8-1:0] x3y5kyk8pk33679m9na1o500m0;
wire  [1:0]                 qxlwggw4wsgzonfuseo_pxc0;
wire  [1:0]                 wouml_54ky8eqv944y579n_qxq;
wire                        ozxqwwwzp4tdkef1udq1k9io69;
wire                        iyzrt9begsn1vu57u29myyut79n_g;
wire                        vc9gmmgtdr7kzh38v5j8gi;
wire                        fm8pi4mpn8uavs13t1u7j7we5d;
wire                        csxakpuvys2li42lnx683; 
wire                        q1vioa1dabxncrn32vbvv237e; 

assign   gohm8ye7tw32so = {csxakpuvys2li42lnx683, fm8pi4mpn8uavs13t1u7j7we5d, vc9gmmgtdr7kzh38v5j8gi};
assign   rhrr146mr7lt9h   = {qxlwggw4wsgzonfuseo_pxc0, ppu_9xb8cwtqbebcovtfl6, k4w5f9hywpks8xc21mnzjr, jxcs4f4npbmy89g7pu0dwd680};
assign   io1uhjqtpgin_   = {wouml_54ky8eqv944y579n_qxq, vtpt106_9th9gncs9klumvuhb8m, pz4yvi8rtvnyll9wc_sl8aja8, u5ls7fh44rneoy5rbkg0fjwarn};
assign   iqaziwvuq5463k3 = {m2kzu5wsbvwjfwip3zfvssodc, o2hausg38teon3_2f7g00su02, wcbtej7qnyi8h9j58z7vr134ulj, i770uc76y777jzpfptztemfl};
assign   hs5w0q7r19myj9eezz = {x3y5kyk8pk33679m9na1o500m0, ax7gdpn6yehlgk0b4bcdap_nvs2, s8o7h0k4g9_xuy00hgcfm4d0, q44ggnacf3_7f825zvirlm0owgd0};

wire     j9o8oc6yq3_fysgtjobnt01uqzwx = (d0q_15ed0hmwqygja[2:0] > 3'b010) && (d0q_15ed0hmwqygja[2:0] != 3'b100);
wire     nzf2317tccqob2z6h9ikbg9fh = d0q_15ed0hmwqygja[2];
wire     bl6t_9ry6h3igt9wm = j9o8oc6yq3_fysgtjobnt01uqzwx ^ nzf2317tccqob2z6h9ikbg9fh;
wire     oa_kgnl_1mm8dm1ys = !(nzf2317tccqob2z6h9ikbg9fh ^ hxrmt706n071lic0f7); 

wire     o48_mos4a4ob9xa_kagb    =  (gohm8ye7tw32so > 3'b010) && (gohm8ye7tw32so != 3'b100);
wire     g9di1w52q5woe8u919tn71   = csxakpuvys2li42lnx683;
wire     hzkgfxff7gsdkbrpx3r_x =  (o48_mos4a4ob9xa_kagb == vc9gmmgtdr7kzh38v5j8gi ) ? xcuko0jmist_fz_ssr0gb4raa2has :
                                 (o48_mos4a4ob9xa_kagb == fm8pi4mpn8uavs13t1u7j7we5d ) ? pizin3jqw9dy383sys4vfakj579 :
                                 (o48_mos4a4ob9xa_kagb == csxakpuvys2li42lnx683 ) ? f2k2cih_4nxcx3c0_a4s15af5d58 : 1'b0;

wire     lvdr9knr1d5l1e3ij_gr =  (o48_mos4a4ob9xa_kagb == vc9gmmgtdr7kzh38v5j8gi ) ? a1rgppa6mdbatjs4nhapuatya :
                                 (o48_mos4a4ob9xa_kagb == fm8pi4mpn8uavs13t1u7j7we5d ) ? eigqul3fdk4hzvxbs_b52aw63 :
                                 (o48_mos4a4ob9xa_kagb == csxakpuvys2li42lnx683 ) ? mqzjxfzpvomdory6rh2y_v8l8wk : 1'b0;


assign   gj95joew8j70jj4 =  (q1vioa1dabxncrn32vbvv237e ? g9di1w52q5woe8u919tn71 : o48_mos4a4ob9xa_kagb) & s7eq8f6z1uyi2in; 
assign   jrkjeqdo7hhdsjna =  (q1vioa1dabxncrn32vbvv237e ? f2k2cih_4nxcx3c0_a4s15af5d58 : hzkgfxff7gsdkbrpx3r_x) & s7eq8f6z1uyi2in;
assign   cmvxg4cmkkrry =  (q1vioa1dabxncrn32vbvv237e ? mqzjxfzpvomdory6rh2y_v8l8wk : lvdr9knr1d5l1e3ij_gr) & s7eq8f6z1uyi2in;



j2erzc_owhcewvkb_q1j #(
  .iomfaylbnp5kdw(0), 
  .y3p_4z5zrymxb1pgv(0)
)h0vj4kq_xobtca75w3bld1ga_q7cxccp(
 .pz6cvxcjpgv        (pz6cvxcjpgv), 
 .z1p1oekb0pd        (js_7wqgsstbnxcjr29), 
 .iq5y0wse0y2       (iq5y0wse0y2),
 .bnjz04i86zhxx6       (bnjz04i86zhxx6),
 .qpotfvbjdo6qtsy1      (qpotfvbjdo6qtsy1),
 .m_pst8fyu48q6i4       (m_pst8fyu48q6i4),
 .jvcw7os6duv6_6       (jvcw7os6duv6_6),
 .k0q5465tih57fj      (k0q5465tih57fj),
 .bl6t_9ry6h3igt9wm    (1'b1),
 .d0q_15ed0hmwqygja  (d0q_15ed0hmwqygja[0]),
 .q1zci4ybfd7ftj8qxl2   (q1zci4ybfd7ftj8qxl2[1:0]),
 .horqgj1y_r_5aplro     (horqgj1y_r_5aplro[8-1:0]),
 .h1wgjzny5b2pljqb7ri(h1wgjzny5b2pljqb7ri),
 .hxrmt706n071lic0f7    (hxrmt706n071lic0f7),
 .v3e6l1k7eo9k3     (wt74a9t1bcclq_xftx2),
 .hwpkcsh2atrq      (hwpkcsh2atrq),
 .iqaziwvuq5463k3    (i770uc76y777jzpfptztemfl),
 .hs5w0q7r19myj9eezz    (q44ggnacf3_7f825zvirlm0owgd0),
 .rhrr146mr7lt9h      (jxcs4f4npbmy89g7pu0dwd680),
 .io1uhjqtpgin_      (u5ls7fh44rneoy5rbkg0fjwarn),
 .jrkjeqdo7hhdsjna    (xcuko0jmist_fz_ssr0gb4raa2has),
 .cmvxg4cmkkrry    (a1rgppa6mdbatjs4nhapuatya),
 .gj95joew8j70jj4       (vc9gmmgtdr7kzh38v5j8gi),
 .gf33atgy              (gf33atgy),
 .ru_wi            (ru_wi)
);


j2erzc_owhcewvkb_q1j #(
  .iomfaylbnp5kdw(1), 
  .y3p_4z5zrymxb1pgv(1)
)q91cpb2g5h6uc3nhxt2qm9xm54ti0faxs(
 .pz6cvxcjpgv        (pz6cvxcjpgv), 
 .z1p1oekb0pd        (js_7wqgsstbnxcjr29), 
 .iq5y0wse0y2       (iq5y0wse0y2),
 .bnjz04i86zhxx6       (bnjz04i86zhxx6),
 .qpotfvbjdo6qtsy1      (qpotfvbjdo6qtsy1),
 .m_pst8fyu48q6i4       (m_pst8fyu48q6i4),
 .jvcw7os6duv6_6       (jvcw7os6duv6_6),
 .k0q5465tih57fj      (k0q5465tih57fj),
 .bl6t_9ry6h3igt9wm    (1'b1),
 .d0q_15ed0hmwqygja  (d0q_15ed0hmwqygja[1]),
 .q1zci4ybfd7ftj8qxl2   (q1zci4ybfd7ftj8qxl2[3:2]),
 .horqgj1y_r_5aplro     (horqgj1y_r_5aplro[2*8-1:8]),
 .h1wgjzny5b2pljqb7ri(h1wgjzny5b2pljqb7ri),
 .hxrmt706n071lic0f7    (hxrmt706n071lic0f7),
 .v3e6l1k7eo9k3     (wt74a9t1bcclq_xftx2),
 .hwpkcsh2atrq      (hwpkcsh2atrq),
 .iqaziwvuq5463k3    (wcbtej7qnyi8h9j58z7vr134ulj),
 .hs5w0q7r19myj9eezz    (s8o7h0k4g9_xuy00hgcfm4d0),
 .rhrr146mr7lt9h      (k4w5f9hywpks8xc21mnzjr),
 .io1uhjqtpgin_      (pz4yvi8rtvnyll9wc_sl8aja8),
 .jrkjeqdo7hhdsjna    (pizin3jqw9dy383sys4vfakj579),
 .cmvxg4cmkkrry    (eigqul3fdk4hzvxbs_b52aw63),
 .gj95joew8j70jj4       (fm8pi4mpn8uavs13t1u7j7we5d),
 .gf33atgy              (gf33atgy),
 .ru_wi            (ru_wi)
);

j2erzc_owhcewvkb_q1j #(
  .iomfaylbnp5kdw(2),  
  .y3p_4z5zrymxb1pgv(0)
)s9igz2x3_tayp6wifps0xk3_6zv49da3t9(
 .pz6cvxcjpgv        (pz6cvxcjpgv), 
 .z1p1oekb0pd        (js_7wqgsstbnxcjr29), 
 .iq5y0wse0y2       (iq5y0wse0y2),
 .bnjz04i86zhxx6       (bnjz04i86zhxx6),
 .qpotfvbjdo6qtsy1      (qpotfvbjdo6qtsy1),
 .m_pst8fyu48q6i4       (m_pst8fyu48q6i4),
 .jvcw7os6duv6_6       (jvcw7os6duv6_6),
 .k0q5465tih57fj      (k0q5465tih57fj),
 .bl6t_9ry6h3igt9wm    (1'b1),
 .d0q_15ed0hmwqygja  (d0q_15ed0hmwqygja[2]),
 .q1zci4ybfd7ftj8qxl2   (q1zci4ybfd7ftj8qxl2[5:4]),
 .horqgj1y_r_5aplro     (horqgj1y_r_5aplro[3*8-1:2*8]),
 .h1wgjzny5b2pljqb7ri(h1wgjzny5b2pljqb7ri),
 .hxrmt706n071lic0f7    (hxrmt706n071lic0f7),
 .v3e6l1k7eo9k3     (wt74a9t1bcclq_xftx2),
 .hwpkcsh2atrq      (hwpkcsh2atrq),
 .iqaziwvuq5463k3    (o2hausg38teon3_2f7g00su02),
 .hs5w0q7r19myj9eezz    (ax7gdpn6yehlgk0b4bcdap_nvs2),
 .rhrr146mr7lt9h      (ppu_9xb8cwtqbebcovtfl6),
 .io1uhjqtpgin_      (vtpt106_9th9gncs9klumvuhb8m),
 .jrkjeqdo7hhdsjna    (f2k2cih_4nxcx3c0_a4s15af5d58),
 .cmvxg4cmkkrry    (mqzjxfzpvomdory6rh2y_v8l8wk),
 .gj95joew8j70jj4       (csxakpuvys2li42lnx683),
 .gf33atgy(gf33atgy),
 .ru_wi(ru_wi)
);


j2erzc_owhcewvkb_q1j #(
  .iomfaylbnp5kdw(3), 
  .y3p_4z5zrymxb1pgv(1)
)rmk9si1hgbpd1tq42vyvxbj_4f_o9y3(
 .pz6cvxcjpgv        (pz6cvxcjpgv), 
 .z1p1oekb0pd        (js_7wqgsstbnxcjr29), 
 .iq5y0wse0y2       (iq5y0wse0y2),
 .bnjz04i86zhxx6       (bnjz04i86zhxx6),
 .qpotfvbjdo6qtsy1      (qpotfvbjdo6qtsy1),
 .m_pst8fyu48q6i4       (m_pst8fyu48q6i4),
 .jvcw7os6duv6_6       (jvcw7os6duv6_6),
 .k0q5465tih57fj      (k0q5465tih57fj),
 .bl6t_9ry6h3igt9wm    (bl6t_9ry6h3igt9wm),
 .d0q_15ed0hmwqygja  (1'b0),
 .q1zci4ybfd7ftj8qxl2   (q1zci4ybfd7ftj8qxl2[7:6]),
 .horqgj1y_r_5aplro     (horqgj1y_r_5aplro[4*8-1:3*8]),
 .h1wgjzny5b2pljqb7ri(h1wgjzny5b2pljqb7ri),
 .hxrmt706n071lic0f7    (oa_kgnl_1mm8dm1ys),
 .v3e6l1k7eo9k3     (wt74a9t1bcclq_xftx2),
 .hwpkcsh2atrq      (hwpkcsh2atrq),
 .iqaziwvuq5463k3    (m2kzu5wsbvwjfwip3zfvssodc),
 .hs5w0q7r19myj9eezz    (x3y5kyk8pk33679m9na1o500m0),
 .rhrr146mr7lt9h      (qxlwggw4wsgzonfuseo_pxc0),
 .io1uhjqtpgin_      (wouml_54ky8eqv944y579n_qxq),
 .jrkjeqdo7hhdsjna    (ozxqwwwzp4tdkef1udq1k9io69),
 .cmvxg4cmkkrry    (iyzrt9begsn1vu57u29myyut79n_g),
 .gj95joew8j70jj4       (q1vioa1dabxncrn32vbvv237e),
 .gf33atgy(gf33atgy),
 .ru_wi(ru_wi)
);





localparam uiscsj0ggxny4qsi = 1+64+9; 

wire [64-1:0] kwvtupo;
wire [9-1:0] p7catsccgqg9wuhtqc;
wire [9-1:0] c695qtwp4kj548m;
l04yr52g7m6wt2i7hqm2aw  wmyalu09heh_88b_2qh9wdpaej1(pz6cvxcjpgv, p7catsccgqg9wuhtqc);
l04yr52g7m6wt2i7hqm2aw  qulw4t9i5ka2huu9e3nkq8a__n(z1p1oekb0pd, c695qtwp4kj548m);
assign m2_t547jr8crh6jgy4c = qpotfvbjdo6qtsy1 ? p7catsccgqg9wuhtqc : c695qtwp4kj548m;
wire g0ypjo0t4_n2wq = v_k8ohy_e2e9vlp6az04; 
wire pa3159orjs0c7fzs = v7rzl8qveorn2jg6659m69;


wire [4-1:0] rh8uk7p_ab7;
wire [uiscsj0ggxny4qsi-1:0] s5z2_2_bh_kf = (g0ypjo0t4_n2wq | pa3159orjs0c7fzs)  ? {1'b1,p54semfzu2zyfb,y_vw514j6xmphhfhc} : {uiscsj0ggxny4qsi{1'b0}};

wire [4-1:0] yx4azp2s7xg9gwb;
wire [4-1:0] gbgwpg279vpb0lar;
wire [uiscsj0ggxny4qsi-1:0] nym1mjycr7iaotj[0:4-1];
generate
    for(i=0;i<4;i=i+1) begin:kac2z2lmdgv3hyzvdl48j 
        assign yx4azp2s7xg9gwb[i] = (nym1mjycr7iaotj[i][uiscsj0ggxny4qsi-2 -: 9] == m2_t547jr8crh6jgy4c) & nym1mjycr7iaotj[i][uiscsj0ggxny4qsi-1];
        assign gbgwpg279vpb0lar[i] =  nym1mjycr7iaotj[i][uiscsj0ggxny4qsi-1]; 
    end
endgenerate

integer nzd5e;
reg [uiscsj0ggxny4qsi-1:0] dfrvd_zgwdya0g_;
reg [2-1:0] nfzsawv303q959_9i9;
always @(*) begin
        dfrvd_zgwdya0g_ = {uiscsj0ggxny4qsi{1'b0}};
        nfzsawv303q959_9i9 = 2'b0;
    for(nzd5e=0;nzd5e<4;nzd5e=nzd5e+1) begin:xungopik1hk90uze3yyc 
        dfrvd_zgwdya0g_ = dfrvd_zgwdya0g_ | ({uiscsj0ggxny4qsi{yx4azp2s7xg9gwb[nzd5e]}} & nym1mjycr7iaotj[nzd5e]);
        nfzsawv303q959_9i9 = nfzsawv303q959_9i9 | ({2{yx4azp2s7xg9gwb[nzd5e]}} & $unsigned(nzd5e[2-1:0]));
    end
end

assign g1iutrfs = |yx4azp2s7xg9gwb;
assign dwz7mnj7ox5 = nfzsawv303q959_9i9;

wire [64-1:0] emumg2cintt8ejip = dfrvd_zgwdya0g_[0 +: 64];





wire [n8duywjqdzotwzmrk9_pvp-1:0] gn6izsi_0245qw_;
wire szzun48kzh6tzdu = &gbgwpg279vpb0lar; 
wire [n8duywjqdzotwzmrk9_pvp-1:0] c1yipthvqif8bij;
wire [4-1:0] oai_mut7mosalu;
wire [4-1:0] woeys9p57z7rn51v1;
wire [4-1:0] y8xt0av09z_y5vt8v3hiizwwmdw; 

generate
if(4 ==16) begin:bicdcir425


















































    assign y8xt0av09z_y5vt8v3hiizwwmdw =  ( 16'b1 << gtvau5cygdmb10dr_makqf);

    assign oai_mut7mosalu[0]  = ~gn6izsi_0245qw_[7]  &  ~gn6izsi_0245qw_[3] & ~gn6izsi_0245qw_[1] &  ~gn6izsi_0245qw_[0] & szzun48kzh6tzdu;
    assign oai_mut7mosalu[1]  =  gn6izsi_0245qw_[7]  &  ~gn6izsi_0245qw_[3] & ~gn6izsi_0245qw_[1] &  ~gn6izsi_0245qw_[0] & szzun48kzh6tzdu;
    assign oai_mut7mosalu[2]  = ~gn6izsi_0245qw_[8]  &   gn6izsi_0245qw_[3] & ~gn6izsi_0245qw_[1] &  ~gn6izsi_0245qw_[0] & szzun48kzh6tzdu;
    assign oai_mut7mosalu[3]  =  gn6izsi_0245qw_[8]  &   gn6izsi_0245qw_[3] & ~gn6izsi_0245qw_[1] &  ~gn6izsi_0245qw_[0] & szzun48kzh6tzdu;
    assign oai_mut7mosalu[4]  = ~gn6izsi_0245qw_[9]  &  ~gn6izsi_0245qw_[4] &  gn6izsi_0245qw_[1] &  ~gn6izsi_0245qw_[0] & szzun48kzh6tzdu;
    assign oai_mut7mosalu[5]  =  gn6izsi_0245qw_[9]  &  ~gn6izsi_0245qw_[4] &  gn6izsi_0245qw_[1] &  ~gn6izsi_0245qw_[0] & szzun48kzh6tzdu;
    assign oai_mut7mosalu[6]  = ~gn6izsi_0245qw_[10] &   gn6izsi_0245qw_[4] &  gn6izsi_0245qw_[1] &  ~gn6izsi_0245qw_[0] & szzun48kzh6tzdu;
    assign oai_mut7mosalu[7]  =  gn6izsi_0245qw_[10] &   gn6izsi_0245qw_[4] &  gn6izsi_0245qw_[1] &  ~gn6izsi_0245qw_[0] & szzun48kzh6tzdu;
    assign oai_mut7mosalu[8]  = ~gn6izsi_0245qw_[11] &  ~gn6izsi_0245qw_[5] & ~gn6izsi_0245qw_[2] &   gn6izsi_0245qw_[0] & szzun48kzh6tzdu;
    assign oai_mut7mosalu[9]  =  gn6izsi_0245qw_[11] &  ~gn6izsi_0245qw_[5] & ~gn6izsi_0245qw_[2] &   gn6izsi_0245qw_[0] & szzun48kzh6tzdu;
    assign oai_mut7mosalu[10] = ~gn6izsi_0245qw_[12] &   gn6izsi_0245qw_[5] & ~gn6izsi_0245qw_[2] &   gn6izsi_0245qw_[0] & szzun48kzh6tzdu;
    assign oai_mut7mosalu[11] =  gn6izsi_0245qw_[12] &   gn6izsi_0245qw_[5] & ~gn6izsi_0245qw_[2] &   gn6izsi_0245qw_[0] & szzun48kzh6tzdu;
    assign oai_mut7mosalu[12] = ~gn6izsi_0245qw_[13] &  ~gn6izsi_0245qw_[6] &  gn6izsi_0245qw_[2] &   gn6izsi_0245qw_[0] & szzun48kzh6tzdu;
    assign oai_mut7mosalu[13] =  gn6izsi_0245qw_[13] &  ~gn6izsi_0245qw_[6] &  gn6izsi_0245qw_[2] &   gn6izsi_0245qw_[0] & szzun48kzh6tzdu;
    assign oai_mut7mosalu[14] = ~gn6izsi_0245qw_[14] &   gn6izsi_0245qw_[6] &  gn6izsi_0245qw_[2] &   gn6izsi_0245qw_[0] & szzun48kzh6tzdu;
    assign oai_mut7mosalu[15] =  gn6izsi_0245qw_[14] &   gn6izsi_0245qw_[6] &  gn6izsi_0245qw_[2] &   gn6izsi_0245qw_[0] & szzun48kzh6tzdu;

    assign c1yipthvqif8bij = ({15{woeys9p57z7rn51v1[0]}} & {gn6izsi_0245qw_[14:8],1'b1,gn6izsi_0245qw_[6:4],1'b1,gn6izsi_0245qw_[2], 2'b11}) |
                             ({15{woeys9p57z7rn51v1[1]}} & {gn6izsi_0245qw_[14:8],1'b0,gn6izsi_0245qw_[6:4],1'b1,gn6izsi_0245qw_[2], 2'b11}) |
                             ({15{woeys9p57z7rn51v1[2]}} & {gn6izsi_0245qw_[14:9],1'b1,gn6izsi_0245qw_[7:4],1'b0,gn6izsi_0245qw_[2], 2'b11}) |
                             ({15{woeys9p57z7rn51v1[3]}} & {gn6izsi_0245qw_[14:9],1'b0,gn6izsi_0245qw_[7:4],1'b0,gn6izsi_0245qw_[2], 2'b11}) |
                             ({15{woeys9p57z7rn51v1[4]}} & {gn6izsi_0245qw_[14:10],1'b1,gn6izsi_0245qw_[8:5],1'b1,gn6izsi_0245qw_[3:2], 2'b01}) |
                             ({15{woeys9p57z7rn51v1[5]}} & {gn6izsi_0245qw_[14:10],1'b0,gn6izsi_0245qw_[8:5],1'b1,gn6izsi_0245qw_[3:2], 2'b01}) |
                             ({15{woeys9p57z7rn51v1[6]}} & {gn6izsi_0245qw_[14:11],1'b1,gn6izsi_0245qw_[9:5],1'b0,gn6izsi_0245qw_[3:2], 2'b01}) |
                             ({15{woeys9p57z7rn51v1[7]}} & {gn6izsi_0245qw_[14:11],1'b0,gn6izsi_0245qw_[9:5],1'b0,gn6izsi_0245qw_[3:2], 2'b01}) |
                             ({15{woeys9p57z7rn51v1[8]}} & {gn6izsi_0245qw_[14:12],1'b1,gn6izsi_0245qw_[10:6],1'b1,gn6izsi_0245qw_[4:3],  1'b1,gn6izsi_0245qw_[1],1'b0}) |
                             ({15{woeys9p57z7rn51v1[9]}} & {gn6izsi_0245qw_[14:12],1'b0,gn6izsi_0245qw_[10:6],1'b1,gn6izsi_0245qw_[4:3],  1'b1,gn6izsi_0245qw_[1],1'b0}) |
                             ({15{woeys9p57z7rn51v1[10]}} & {gn6izsi_0245qw_[14:13],1'b1,gn6izsi_0245qw_[11:6],1'b0,gn6izsi_0245qw_[4:3], 1'b1,gn6izsi_0245qw_[1],1'b0}) |
                             ({15{woeys9p57z7rn51v1[11]}} & {gn6izsi_0245qw_[14:13],1'b0,gn6izsi_0245qw_[11:6],1'b0,gn6izsi_0245qw_[4:3], 1'b1,gn6izsi_0245qw_[1],1'b0}) |
                             ({15{woeys9p57z7rn51v1[12]}} & {gn6izsi_0245qw_[14],1'b1,gn6izsi_0245qw_[12:7],1'b1,gn6izsi_0245qw_[5:3],  1'b0,gn6izsi_0245qw_[1],1'b0}) |
                             ({15{woeys9p57z7rn51v1[13]}} & {gn6izsi_0245qw_[14],1'b0,gn6izsi_0245qw_[12:7],1'b1,gn6izsi_0245qw_[5:3],  1'b0,gn6izsi_0245qw_[1],1'b0}) |
                             ({15{woeys9p57z7rn51v1[14]}} & {1'b1,gn6izsi_0245qw_[13:7],1'b0,gn6izsi_0245qw_[5:3], 1'b0,gn6izsi_0245qw_[1],1'b0}) |
                             ({15{woeys9p57z7rn51v1[15]}} & {1'b0,gn6izsi_0245qw_[13:7],1'b0,gn6izsi_0245qw_[5:3], 1'b0,gn6izsi_0245qw_[1],1'b0});
end
else if(4 ==8) begin:bk561






































    assign y8xt0av09z_y5vt8v3hiizwwmdw =  ( 8'b1 << gtvau5cygdmb10dr_makqf);

    assign oai_mut7mosalu[0]  = ~gn6izsi_0245qw_[3] & ~gn6izsi_0245qw_[1] &  ~gn6izsi_0245qw_[0] & szzun48kzh6tzdu;
    assign oai_mut7mosalu[1]  =  gn6izsi_0245qw_[3] & ~gn6izsi_0245qw_[1] &  ~gn6izsi_0245qw_[0] & szzun48kzh6tzdu;
    assign oai_mut7mosalu[2]  = ~gn6izsi_0245qw_[4] &  gn6izsi_0245qw_[1] &  ~gn6izsi_0245qw_[0] & szzun48kzh6tzdu;
    assign oai_mut7mosalu[3]  =  gn6izsi_0245qw_[4] &  gn6izsi_0245qw_[1] &  ~gn6izsi_0245qw_[0] & szzun48kzh6tzdu;
    assign oai_mut7mosalu[4]  = ~gn6izsi_0245qw_[5] & ~gn6izsi_0245qw_[2] &   gn6izsi_0245qw_[0] & szzun48kzh6tzdu;
    assign oai_mut7mosalu[5]  =  gn6izsi_0245qw_[5] & ~gn6izsi_0245qw_[2] &   gn6izsi_0245qw_[0] & szzun48kzh6tzdu;
    assign oai_mut7mosalu[6]  = ~gn6izsi_0245qw_[6] &  gn6izsi_0245qw_[2] &   gn6izsi_0245qw_[0] & szzun48kzh6tzdu;
    assign oai_mut7mosalu[7]  =  gn6izsi_0245qw_[6] &  gn6izsi_0245qw_[2] &   gn6izsi_0245qw_[0] & szzun48kzh6tzdu;



    assign c1yipthvqif8bij = ({7{woeys9p57z7rn51v1[0]}} & {gn6izsi_0245qw_[6:4],1'b1,gn6izsi_0245qw_[2],2'b11})
                           | ({7{woeys9p57z7rn51v1[1]}} & {gn6izsi_0245qw_[6:4],1'b0,gn6izsi_0245qw_[2],2'b11})
                           | ({7{woeys9p57z7rn51v1[2]}} & {gn6izsi_0245qw_[6:5],1'b1,gn6izsi_0245qw_[3:2],2'b01})
                           | ({7{woeys9p57z7rn51v1[3]}} & {gn6izsi_0245qw_[6:5],1'b0,gn6izsi_0245qw_[3:2],2'b01})
                           | ({7{woeys9p57z7rn51v1[4]}} & {gn6izsi_0245qw_[6],1'b1,gn6izsi_0245qw_[4:3],1'b1,gn6izsi_0245qw_[1],1'b0})
                           | ({7{woeys9p57z7rn51v1[5]}} & {gn6izsi_0245qw_[6],1'b0,gn6izsi_0245qw_[4:3],1'b1,gn6izsi_0245qw_[1],1'b0})
                           | ({7{woeys9p57z7rn51v1[6]}} & {1'b1,gn6izsi_0245qw_[5:3],1'b0,gn6izsi_0245qw_[1],1'b0})
                           | ({7{woeys9p57z7rn51v1[7]}} & {1'b0,gn6izsi_0245qw_[5:3],1'b0,gn6izsi_0245qw_[1],1'b0})
                           ;
end
else begin:nha0mie






























    assign y8xt0av09z_y5vt8v3hiizwwmdw =  ( 4'b1 << gtvau5cygdmb10dr_makqf);

    assign oai_mut7mosalu[0]  =  ~gn6izsi_0245qw_[1] &  ~gn6izsi_0245qw_[0] & szzun48kzh6tzdu;
    assign oai_mut7mosalu[1]  =   gn6izsi_0245qw_[1] &  ~gn6izsi_0245qw_[0] & szzun48kzh6tzdu;
    assign oai_mut7mosalu[2]  =  ~gn6izsi_0245qw_[2] &   gn6izsi_0245qw_[0] & szzun48kzh6tzdu;
    assign oai_mut7mosalu[3]  =   gn6izsi_0245qw_[2] &   gn6izsi_0245qw_[0] & szzun48kzh6tzdu;



    assign c1yipthvqif8bij = ({3{woeys9p57z7rn51v1[0]}} & {gn6izsi_0245qw_[2],2'b11})
                           | ({3{woeys9p57z7rn51v1[1]}} & {gn6izsi_0245qw_[2],2'b01})
                           | ({3{woeys9p57z7rn51v1[2]}} & {1'b1,gn6izsi_0245qw_[1],1'b0})
                           | ({3{woeys9p57z7rn51v1[3]}} & {1'b0,gn6izsi_0245qw_[1],1'b0})
                           ;
end
endgenerate

assign woeys9p57z7rn51v1 = vp5_qftup10p3v7_jw8 ? y8xt0av09z_y5vt8v3hiizwwmdw : oai_mut7mosalu;

wire hi62hgv_y1z;
wire kcfm0dqoofinxx90dud = szzun48kzh6tzdu & (g0ypjo0t4_n2wq | vp5_qftup10p3v7_jw8);
ux607_gnrl_dfflr #(n8duywjqdzotwzmrk9_pvp) jr6gmj9vw9yj74bur11(kcfm0dqoofinxx90dud,c1yipthvqif8bij,gn6izsi_0245qw_,gf33atgy,ru_wi); 

wire [4-1:0] herugzgzjy5zca2e80uy2 =  {gbgwpg279vpb0lar[4-2:0],1'b1} ^ gbgwpg279vpb0lar;
wire [4-1:0] tm1p18nx0x1ww3w6zb4y;

generate
for(i=0;i<4;i=i+1) begin:sxq_amt5geudw_mtdr8g2d41y2
    if(i==0) begin:t9w81cc3ejd_
        assign tm1p18nx0x1ww3w6zb4y[i] = herugzgzjy5zca2e80uy2[0];
    end
    else begin:cghdgmfjwlvv
        assign tm1p18nx0x1ww3w6zb4y[i] = |herugzgzjy5zca2e80uy2[i:0];
    end
end
endgenerate

wire [4-1:0] qt5mfy2zxpo0tt21z17ivvy7 = {tm1p18nx0x1ww3w6zb4y[4-2:0],1'b0} ^ tm1p18nx0x1ww3w6zb4y;

wire [4-1:0] euhhrqai6b;

  assign euhhrqai6b =  g0ypjo0t4_n2wq ? (szzun48kzh6tzdu ? oai_mut7mosalu : qt5mfy2zxpo0tt21z17ivvy7)
                                      :  y8xt0av09z_y5vt8v3hiizwwmdw;

wire idyndq1pypwlt = qpotfvbjdo6qtsy1  & (~vkfewi0rkx);
wire tqbfdjlxiac1c = k0q5465tih57fj  & (~z9lf1gw3iz9e);
wire cicg1i1w91s5_ = idyndq1pypwlt ? 1'b1 : (vgno0maw8a & tqbfdjlxiac1c);
assign hi62hgv_y1z =  (g0ypjo0t4_n2wq | pa3159orjs0c7fzs) & s7eq8f6z1uyi2in; 

generate
for(i=0;i<4;i=i+1) begin:gfexls9l1l2nl
    if(4 ==16) begin:axalui_g7g3y
        assign rh8uk7p_ab7[i] = (euhhrqai6b == (16'b1<<i)) & hi62hgv_y1z;
    end
    else if(4 ==8) begin:u0iw0z1nfu9wh4c
        assign rh8uk7p_ab7[i] = (euhhrqai6b == (8'b1<<i)) & hi62hgv_y1z;
    end
    else begin:hckskius5po7
        assign rh8uk7p_ab7[i] = (euhhrqai6b == (4'b1<<i)) & hi62hgv_y1z;
    end
        ux607_gnrl_dfflr #(uiscsj0ggxny4qsi) cu7ld1ljb980w1wblz(rh8uk7p_ab7[i], s5z2_2_bh_kf, nym1mjycr7iaotj[i],gf33atgy, ru_wi);
    end
endgenerate



wire [64-1:0] ygbc6czf = jrkjeqdo7hhdsjna ? pz6cvxcjpgv : z1p1oekb0pd;
wire [64-1:0] bdhv0j4zhtx9nxmz = jrkjeqdo7hhdsjna ? ueimo2s8tf29_f : xl0lr2g890tskf74yu8;
wire l78_ius4cmnzogx4p;
wire lskus_x793x4;
wire aviywg23jao_ad4f = cd3xfhf_7i5g014tqu9;
wire krjcsiswo73ice = lskus_x793x4;
wire b8s56xam46vfi = aviywg23jao_ad4f | krjcsiswo73ice;
wire h5p6lfvmmjno2q = aviywg23jao_ad4f | (~krjcsiswo73ice); 
ux607_gnrl_dfflr #(1) hp60hynux10oen7(b8s56xam46vfi, h5p6lfvmmjno2q, lskus_x793x4, gf33atgy, ru_wi);

localparam u4yrh3l613ygudlvvn54xf = 64 + 2*64 + 2; 
wire a4hsmvk7b78o;
wire [u4yrh3l613ygudlvvn54xf-1:0] szfrddcfc54;
wire [u4yrh3l613ygudlvvn54xf-1:0] zsybyys3zaz;
wire [64-1:0] k4zhwibysy1g0wdq2;
wire [64-1:0] sl4ljoqdgrgf5xq;
wire rj8vqubs4fbhoqdmdbutku;
assign  zsybyys3zaz = { ygbc6czf,
                       cs_6ujj3b74,
                       l78_ius4cmnzogx4p, 
                       gj95joew8j70jj4,
                       bdhv0j4zhtx9nxmz
                       };
assign { kwvtupo,
         sl4ljoqdgrgf5xq,
         rj8vqubs4fbhoqdmdbutku, 
         a4hsmvk7b78o,
         k4zhwibysy1g0wdq2
        }         = szfrddcfc54;

ux607_gnrl_dfflr #(u4yrh3l613ygudlvvn54xf) kxts4ldrv5nb8v(aviywg23jao_ad4f, zsybyys3zaz, szfrddcfc54, gf33atgy, ru_wi);
wire nh1ik6l45z8raeul = (r12cr5tap6v & (~ywsaub3r999h9pyn)) & s7eq8f6z1uyi2in;
wire tvm48wkm3j3 = g1iutrfs & cicg1i1w91s5_ & s7eq8f6z1uyi2in;

assign v4gayo0h8l6na = a4hsmvk7b78o & lskus_x793x4;
wire [64-1:0] ohu0bjo6f234 = (kwvtupo + k4zhwibysy1g0wdq2[64-1:0]);
assign nmy2nw74r7gg = rj8vqubs4fbhoqdmdbutku ? sl4ljoqdgrgf5xq : ohu0bjo6f234;

localparam p_2qaaa2_ubd6_u6xhek0jbxu751qdv = 8 + 2;
wire [64-1:0] iwo1igeb = jrkjeqdo7hhdsjna ? haezj87elp_ : eajem3pnezl;

assign cs_6ujj3b74 = nh1ik6l45z8raeul ? xe0fwqp049g43
                   : tvm48wkm3j3 ? emumg2cintt8ejip
                   : iwo1igeb
                   ;
assign v0u85q8u16_pwgz7h17cl4 = qpotfvbjdo6qtsy1; 
assign yov0d70301nwd4bbqbyv =  (~jrkjeqdo7hhdsjna) & k0q5465tih57fj;
assign l78_ius4cmnzogx4p =  v0u85q8u16_pwgz7h17cl4 | yov0d70301nwd4bbqbyv;

endmodule


module j2erzc_owhcewvkb_q1j #(
    parameter iomfaylbnp5kdw = 0,
    parameter y3p_4z5zrymxb1pgv = 0

) (
  input  [64-1:0]   pz6cvxcjpgv, 
  input  [64-1:0]   z1p1oekb0pd, 
  input                        iq5y0wse0y2,
  input                        bnjz04i86zhxx6,
  input                        qpotfvbjdo6qtsy1,
  input                        m_pst8fyu48q6i4,
  input                        jvcw7os6duv6_6,
  input                        k0q5465tih57fj,
  input                        bl6t_9ry6h3igt9wm,
  input                        d0q_15ed0hmwqygja,
  input  [1:0]                 q1zci4ybfd7ftj8qxl2,
  input  [8-1:0] horqgj1y_r_5aplro,
  input  [8-1:0] h1wgjzny5b2pljqb7ri,
  input                        hxrmt706n071lic0f7,
  input                        v3e6l1k7eo9k3,
  input                        hwpkcsh2atrq,
  output [8-1:0] iqaziwvuq5463k3,
  output [8-1:0] hs5w0q7r19myj9eezz,
  output [1:0]                 rhrr146mr7lt9h,
  output [1:0]                 io1uhjqtpgin_,
  output                       jrkjeqdo7hhdsjna,
  output                       cmvxg4cmkkrry,
  output                       gj95joew8j70jj4,

  input                        gf33atgy,
  input                        ru_wi
);

localparam ji61pdozd8f3gq4938iy = 256 >> y3p_4z5zrymxb1pgv;
wire [ji61pdozd8f3gq4938iy-1:0] ak93fzwbz6_y4l;
wire [ji61pdozd8f3gq4938iy-1:0] wsgwrutpw75o4;
wire [ji61pdozd8f3gq4938iy-1:0] gghojhrb3mb4hz28i;
wire [ji61pdozd8f3gq4938iy-1:0] bfkih8wqvcqfmw;
wire [1:0] txnz6o1bihuu4ottib9r [0:ji61pdozd8f3gq4938iy-1];

b83pl9mk1y2z58pcocbgh #(iomfaylbnp5kdw) ppbwccpy6z6bnq8mrtup5j47(pz6cvxcjpgv, h1wgjzny5b2pljqb7ri, iqaziwvuq5463k3);
b83pl9mk1y2z58pcocbgh #(iomfaylbnp5kdw) jlnl665nxxawv8ra2xlhg2o(z1p1oekb0pd, h1wgjzny5b2pljqb7ri, hs5w0q7r19myj9eezz);

wire [1:0] i4q4ffjklbhi6fad;
generate 
 if (iomfaylbnp5kdw == 3) begin: ysowyz834__amh1w
   assign i4q4ffjklbhi6fad[1] = (q1zci4ybfd7ftj8qxl2[1] & q1zci4ybfd7ftj8qxl2[0]) | (q1zci4ybfd7ftj8qxl2[0] & hxrmt706n071lic0f7) | (q1zci4ybfd7ftj8qxl2[1] & hxrmt706n071lic0f7); 
   assign i4q4ffjklbhi6fad[0] = !hxrmt706n071lic0f7;
 end
 else begin: xf2lctmwm266j7v69zpq
   assign i4q4ffjklbhi6fad[1] = (q1zci4ybfd7ftj8qxl2[1] & q1zci4ybfd7ftj8qxl2[0]) | (!q1zci4ybfd7ftj8qxl2[0] & hxrmt706n071lic0f7); 
   assign i4q4ffjklbhi6fad[0] = (q1zci4ybfd7ftj8qxl2[1] & hxrmt706n071lic0f7) | (!q1zci4ybfd7ftj8qxl2[1] & !hxrmt706n071lic0f7);
  end
endgenerate 

genvar i;
wire [1:0] qwlu67h3_7y2a = i4q4ffjklbhi6fad;
wire       jl2zgroagizditrkrcflw75 = ~hwpkcsh2atrq & (hxrmt706n071lic0f7 == d0q_15ed0hmwqygja);
 generate

      for (i=0; i<ji61pdozd8f3gq4938iy;i=i+1) begin: dxij2dw1p5i52hoalv
          assign ak93fzwbz6_y4l[i] = (horqgj1y_r_5aplro == $unsigned(i[8-1:0]));
          if ( iomfaylbnp5kdw == 3) begin: ouowg6gft0ema8wb
            assign wsgwrutpw75o4[i] = bl6t_9ry6h3igt9wm & v3e6l1k7eo9k3 & ak93fzwbz6_y4l[i]; 
          end 
          else begin : g4lh30hfs2ssquhvnrh
            assign wsgwrutpw75o4[i] = (hwpkcsh2atrq | jl2zgroagizditrkrcflw75) & v3e6l1k7eo9k3 & ak93fzwbz6_y4l[i] & bl6t_9ry6h3igt9wm; 
          end

         ux607_gnrl_dfflr #(2) mwdl1qmtvn_ui667lv (wsgwrutpw75o4[i], qwlu67h3_7y2a, txnz6o1bihuu4ottib9r[i], gf33atgy, ru_wi);

         assign gghojhrb3mb4hz28i[i] = (iqaziwvuq5463k3 == $unsigned(i[8-1:0]));
         assign bfkih8wqvcqfmw[i] = (hs5w0q7r19myj9eezz == $unsigned(i[8-1:0]));
      end
  endgenerate

   reg [1:0] mfkrfmi7cybk2nw97;
   reg [1:0] gpxbyslsrqxa763fqh;

   integer nzd5e;

   always @* begin:cp2t3voyssrtlzqh
       mfkrfmi7cybk2nw97 = 2'b0;
       gpxbyslsrqxa763fqh = 2'b0;

       for(nzd5e=0; nzd5e<ji61pdozd8f3gq4938iy; nzd5e=nzd5e+1) begin: l7thhsn6_f3p
         mfkrfmi7cybk2nw97 = mfkrfmi7cybk2nw97 | ({2{gghojhrb3mb4hz28i[nzd5e]}} & txnz6o1bihuu4ottib9r[nzd5e]);
         gpxbyslsrqxa763fqh = gpxbyslsrqxa763fqh | ({2{bfkih8wqvcqfmw[nzd5e]}} & txnz6o1bihuu4ottib9r[nzd5e]);
       end
   end

assign rhrr146mr7lt9h = mfkrfmi7cybk2nw97;
assign io1uhjqtpgin_ = gpxbyslsrqxa763fqh;

generate 
  if (iomfaylbnp5kdw == 3) begin: s6t_3_solj27klz
    assign jrkjeqdo7hhdsjna = rhrr146mr7lt9h[1];
    assign cmvxg4cmkkrry = io1uhjqtpgin_[1];
  end 
  else begin: o48_mos4a4ob9xa_kagb
    assign jrkjeqdo7hhdsjna = ((rhrr146mr7lt9h[1] & iq5y0wse0y2) | bnjz04i86zhxx6 | qpotfvbjdo6qtsy1);
    assign cmvxg4cmkkrry = ((io1uhjqtpgin_[1] & m_pst8fyu48q6i4) | jvcw7os6duv6_6 | k0q5465tih57fj);
  end
endgenerate

assign gj95joew8j70jj4 = jrkjeqdo7hhdsjna | cmvxg4cmkkrry; 

endmodule 




module b83pl9mk1y2z58pcocbgh #(
    parameter iomfaylbnp5kdw = 0
) (
    input [64-1:0] k4p2,
    input [8-1:0] ghpk,
    output [8-1:0] wo008jpoe
);

 generate 
   if (iomfaylbnp5kdw == 0 || iomfaylbnp5kdw == 3) begin: bjnces_oe_
     wire [8:0] rirj80qeof_vbhu = k4p2[18:10] ^ k4p2[10:2];
     wire [1:0] ua8b3abbvcxpux2o = ghpk[7:6] ^ ghpk[4:3] ^ ghpk[1:0]; 
     assign wo008jpoe = {ua8b3abbvcxpux2o^rirj80qeof_vbhu[7:6],rirj80qeof_vbhu[5:0]}; 
   end
   else if (iomfaylbnp5kdw == 1) begin : shsrzcx82vo
     wire [8:0] rirj80qeof_vbhu = k4p2[18:10] ^ k4p2[10:2];
     assign wo008jpoe =  ghpk ^ rirj80qeof_vbhu[7:0]; 
   end 
   else begin : zfcj4ba
       assign wo008jpoe = k4p2[8:2];
   end
 endgenerate 


endmodule

module l04yr52g7m6wt2i7hqm2aw (
    input [64-1:0] k4p2,
    output [9-1:0] wo008jpoe
);

assign wo008jpoe = k4p2[9*2 - 1 : 9] ^
              k4p2[9:1];
endmodule









module tr81ezgbvz5391e_kkgo4g3lvka05 # (
  parameter tcebpmbl7g = 0,
  parameter mhdlk   = 8,
  parameter onr7l   = 32
) (

  input           veibgbyke,

  input           bw6ftrau0, 
  output          eef2g8, 
  input  [onr7l-1:0] qbjvs30wtb,
  output          wqljp, 
  input           h9378, 
  output [onr7l-1:0] dqgck5s,
  output          p3mxtqc2ivbcmm0,

  input           gf33atgy,
  input           ru_wi
);



    wire [onr7l-1:0] w2z87rfaf8 [mhdlk-1:0];
    wire [mhdlk-1:0] k8cq9veedzws;


    wire kxaplzy = (bw6ftrau0 & eef2g8);
    wire fumg8 = (wqljp & h9378);



    wire [mhdlk-1:0] tzr9_pu0gkgq459gy; 
    wire [mhdlk-1:0] dz1thuu43r;
    wire [mhdlk-1:0] kv5lv5mhl4m9_kh; 
    wire [mhdlk-1:0] wxlsjrqo2a;

    assign tzr9_pu0gkgq459gy = 
          veibgbyke ? { {mhdlk-1{1'b0}}, 1'b1 } :
          dz1thuu43r[mhdlk-1] ? {{mhdlk-1{1'b0}}, 1'b1} :
                          (dz1thuu43r << 1);

    assign kv5lv5mhl4m9_kh =
          veibgbyke ? { {mhdlk-1{1'b0}}, 1'b1 } :
          wxlsjrqo2a[mhdlk-1] ? {{mhdlk-1{1'b0}}, 1'b1} :
                          (wxlsjrqo2a << 1);

    ux607_gnrl_dfflrs #(1)    qnwogo1l036nyvzk_i  ((fumg8 | veibgbyke), tzr9_pu0gkgq459gy[0]     , dz1thuu43r[0]     , gf33atgy, ru_wi);
    ux607_gnrl_dfflrs #(1)    mn4pzjreki9yvykae  ((kxaplzy | veibgbyke), kv5lv5mhl4m9_kh[0]     , wxlsjrqo2a[0]     , gf33atgy, ru_wi);
    ux607_gnrl_dfflr  #(mhdlk-1) fipb6zpafcl9yge96au  ((fumg8 | veibgbyke), tzr9_pu0gkgq459gy[mhdlk-1:1], dz1thuu43r[mhdlk-1:1], gf33atgy, ru_wi);
    ux607_gnrl_dfflr  #(mhdlk-1) hh9891_eoeau0wkyll5  ((kxaplzy | veibgbyke), kv5lv5mhl4m9_kh[mhdlk-1:1], wxlsjrqo2a[mhdlk-1:1], gf33atgy, ru_wi);



    wire [mhdlk:0] uipdtjs;
    wire [mhdlk:0] acm0zbhvam;
    wire [mhdlk:0] oi40qurrxr; 
    wire [mhdlk:0] n89fv;

    wire jlo7_b_z = (fumg8 ^ kxaplzy ) | veibgbyke;
    assign oi40qurrxr = veibgbyke ? { {mhdlk{1'b0}}, 1'b1 } : kxaplzy ? {n89fv[mhdlk-1:0], 1'b1} : (n89fv >> 1);  

    ux607_gnrl_dfflrs #(1)  svv3sz17bdpp     (jlo7_b_z, oi40qurrxr[0]     , n89fv[0]     ,     gf33atgy, ru_wi);
    ux607_gnrl_dfflr  #(mhdlk) j3hui4o9q5lg     (jlo7_b_z, oi40qurrxr[mhdlk:1], n89fv[mhdlk:1],     gf33atgy, ru_wi);

    assign uipdtjs = {1'b0,n89fv[mhdlk:1]};
    assign acm0zbhvam = {1'b0,n89fv[mhdlk:1]};



    genvar i;
    generate 


    if(tcebpmbl7g==1) begin: lvfon_zgkwp229
    assign eef2g8 = (~uipdtjs[mhdlk-1]);

    assign p3mxtqc2ivbcmm0 = (~uipdtjs[1]);
    end
    else begin:ugkahrezmhzxybh191t
    assign eef2g8 = (~uipdtjs[mhdlk-1]) | fumg8;

    assign p3mxtqc2ivbcmm0 = (~uipdtjs[1]) | (fumg8 & (~kxaplzy) & ~uipdtjs[2]);

    end

      for (i=0; i<mhdlk; i=i+1) begin:m_wwntxzhohqg5
        assign k8cq9veedzws[i] = kxaplzy & wxlsjrqo2a[i];

        ux607_gnrl_dfflr  #(onr7l) c9h7cqhau6oedhp (k8cq9veedzws[i], qbjvs30wtb, w2z87rfaf8[i], gf33atgy, ru_wi);
      end

    endgenerate


    integer j;
    reg [onr7l-1:0] ui9y38d1t;
    always @*
    begin : e82692n5bc4eh
      ui9y38d1t = {onr7l{1'b0}};
      for(j=0; j<mhdlk; j=j+1) begin
        ui9y38d1t = ui9y38d1t | ({onr7l{dz1thuu43r[j]}} & w2z87rfaf8[j]);
      end
    end



    assign dqgck5s = ui9y38d1t;


    assign wqljp = (acm0zbhvam[0]);


endmodule 


module bh912j8o17nne6z_zsk9c #(
  parameter tcebpmbl7g= 0,
  parameter mhdlk = 8,
  parameter onr7l = 32
) (
  input           veibgbyke,
  input           bw6ftrau0,
  output          eef2g8,
  output          p3mxtqc2ivbcmm0,
  input  [onr7l-1:0] qbjvs30wtb,

  output          wqljp,
  input           h9378,
  output [onr7l-1:0] dqgck5s,

  input           gf33atgy,
  input           ru_wi
);
  wire          bskljx6b_bvnqj4h;
  wire          zvyiwdpyvt;
  wire          o0ozobxf1oc2t5;
  wire [onr7l-1:0] jf92hqkj0cxz;

  wire          mgjqsgpiza1dr;
  wire          qos62pcur8;
  wire [onr7l-1:0] jae1i1kz83d2c;
  wire          pzbrn1v8f4udbk0tm;



  generate 
  if(mhdlk == 1) begin: oo11sjc9w
    ac6zxmzb4w0hgrfychpxv_xj # (
         .tcebpmbl7g(tcebpmbl7g),
         .mhdlk(mhdlk),
         .onr7l(onr7l)
    ) bds_ov5rlhhtc6aixp8cra013a(
      .veibgbyke (bskljx6b_bvnqj4h),
      .bw6ftrau0   (zvyiwdpyvt),
      .eef2g8   (o0ozobxf1oc2t5),
      .qbjvs30wtb   (jf92hqkj0cxz),
      .wqljp   (mgjqsgpiza1dr),
      .h9378   (qos62pcur8),
      .dqgck5s   (jae1i1kz83d2c),
      .gf33atgy     (gf33atgy  ),
      .ru_wi   (ru_wi)
    );
    assign pzbrn1v8f4udbk0tm = 1'b0;

  end
  else begin: rwwqt_zj36eixlt3

    tr81ezgbvz5391e_kkgo4g3lvka05 # (
         .tcebpmbl7g(tcebpmbl7g),
         .mhdlk(mhdlk),
         .onr7l(onr7l)
    ) bds_ov5rlhhtc6aixp8cra013a(
      .veibgbyke (bskljx6b_bvnqj4h),
      .bw6ftrau0   (zvyiwdpyvt),
      .eef2g8   (o0ozobxf1oc2t5),
      .qbjvs30wtb   (jf92hqkj0cxz),
      .wqljp   (mgjqsgpiza1dr),
      .h9378   (qos62pcur8),
      .dqgck5s   (jae1i1kz83d2c),
      .p3mxtqc2ivbcmm0(pzbrn1v8f4udbk0tm),
      .gf33atgy     (gf33atgy  ),
      .ru_wi   (ru_wi)
    );
  end
  endgenerate




  assign bskljx6b_bvnqj4h = veibgbyke;
  assign eef2g8 = o0ozobxf1oc2t5;
  assign p3mxtqc2ivbcmm0 = pzbrn1v8f4udbk0tm;



  wire fzf_yfd = bw6ftrau0 & h9378 & (~mgjqsgpiza1dr);


  assign qos62pcur8 = h9378;


  assign wqljp = mgjqsgpiza1dr | bw6ftrau0;


  assign dqgck5s = mgjqsgpiza1dr ? jae1i1kz83d2c : qbjvs30wtb;

  assign jf92hqkj0cxz  = qbjvs30wtb; 


  assign zvyiwdpyvt = bw6ftrau0 & (~fzf_yfd);

endmodule 

module ixyqarhsqal9rouebde # (
  parameter mhdlk   = 8,
  parameter onr7l   = 32
) (

  input           veibgbyke,

  input           bw6ftrau0, 
  output          eef2g8, 
  input  [onr7l-1:0] qplwyaz47s,
  input  [onr7l-1:0] qdbq74,
  output          wqljp, 
  input           h9378, 
  output [onr7l-1:0] dqgck5s,

  input           gf33atgy,
  input           ru_wi
);



    wire [onr7l-1:0] w2z87rfaf8 [mhdlk-1:0];
    wire [mhdlk-1:0] k8cq9veedzws;
    wire [mhdlk-1:0] fjclvexm6y5j8i;
    wire [mhdlk-1:0] nb3l28dm4ze1u3at;
    wire [onr7l-1:0] z1u1ts_k1h5jrd[mhdlk-1:0];


    wire fk0i0zw0m7z = (bw6ftrau0 & eef2g8);
    wire fumg8 = (wqljp & h9378);
    wire n1kgjxrls = fk0i0zw0m7z & qplwyaz47s[onr7l-1];
    wire d0yt9d65 = fk0i0zw0m7z & qdbq74[onr7l-1];
    wire kxg2usnf2g = n1kgjxrls & d0yt9d65;
    wire kxaplzy = n1kgjxrls | d0yt9d65;



    wire [mhdlk-1:0] tzr9_pu0gkgq459gy; 
    wire [mhdlk-1:0] dz1thuu43r;
    wire [mhdlk-1:0] kv5lv5mhl4m9_kh; 
    wire [mhdlk-1:0] wxlsjrqo2a;
    wire [mhdlk-1:0] wgnqmwnpaqxd3yvuxe_qr0 = wxlsjrqo2a << 1;

    wire [mhdlk-1:0] g9j6_wgc1qjli77u = wxlsjrqo2a;
    wire [mhdlk-1:0] lw3x2mny6rj = wxlsjrqo2a[mhdlk-1] ? {{mhdlk-1{1'b0}}, 1'b1} : wgnqmwnpaqxd3yvuxe_qr0;

    assign tzr9_pu0gkgq459gy = 
          veibgbyke ? { {mhdlk-1{1'b0}}, 1'b1 } :
          dz1thuu43r[mhdlk-1] ? {{mhdlk-1{1'b0}}, 1'b1} :
                          (dz1thuu43r << 1);

    assign kv5lv5mhl4m9_kh =
          veibgbyke ? { {mhdlk-1{1'b0}}, 1'b1 } :
          wxlsjrqo2a[mhdlk-1] ? (kxg2usnf2g ? {{mhdlk-2{1'b0}}, 2'b10} : {{mhdlk-1{1'b0}}, 1'b1}):
          wxlsjrqo2a[mhdlk-2] ? (kxg2usnf2g ? {{mhdlk-1{1'b0}}, 1'b1}  : wgnqmwnpaqxd3yvuxe_qr0):
                              (kxg2usnf2g ? (wxlsjrqo2a << 2)    : wgnqmwnpaqxd3yvuxe_qr0);

    ux607_gnrl_dfflrs #(1)    qnwogo1l036nyvzk_i  ((fumg8 | veibgbyke), tzr9_pu0gkgq459gy[0]     , dz1thuu43r[0]     , gf33atgy, ru_wi);
    ux607_gnrl_dfflrs #(1)    mn4pzjreki9yvykae ((kxaplzy | veibgbyke), kv5lv5mhl4m9_kh[0]     , wxlsjrqo2a[0]     , gf33atgy, ru_wi);

    ux607_gnrl_dfflr  #(mhdlk-1) fipb6zpafcl9yge96au  ((fumg8 | veibgbyke), tzr9_pu0gkgq459gy[mhdlk-1:1], dz1thuu43r[mhdlk-1:1], gf33atgy, ru_wi);
    ux607_gnrl_dfflr  #(mhdlk-1) hh9891_eoeau0wkyll5 ((kxaplzy | veibgbyke), kv5lv5mhl4m9_kh[mhdlk-1:1], wxlsjrqo2a[mhdlk-1:1], gf33atgy, ru_wi);




    wire [mhdlk:0] uipdtjs;
    wire [mhdlk:0] acm0zbhvam;
    wire [mhdlk:0] oi40qurrxr; 
    wire [mhdlk:0] n89fv;

    wire jlo7_b_z = veibgbyke
                | (~(   (~(fumg8 | n1kgjxrls | d0yt9d65)) 
                      | (fumg8 & (n1kgjxrls ^ d0yt9d65))  
                    ))
                ;
    assign oi40qurrxr =                    veibgbyke ? {{mhdlk{1'b0}}, 1'b1 } : 
                        ((~fumg8) & n1kgjxrls & d0yt9d65)  ? {n89fv[mhdlk-2:0], 2'b11} :
                      (fumg8 & (~n1kgjxrls) & (~d0yt9d65)) ? (n89fv >> 1) 
                                                : {n89fv[mhdlk-1:0], 1'b1}
                                                ;

    ux607_gnrl_dfflrs #(1)  svv3sz17bdpp     (jlo7_b_z, oi40qurrxr[0]   , n89fv[0]   ,     gf33atgy, ru_wi);
    ux607_gnrl_dfflr  #(mhdlk) j3hui4o9q5lg     (jlo7_b_z, oi40qurrxr[mhdlk:1], n89fv[mhdlk:1],     gf33atgy, ru_wi);

    assign uipdtjs = {1'b0,n89fv[mhdlk:1]};
    assign acm0zbhvam = {1'b0,n89fv[mhdlk:1]};



    genvar i;
    generate 





    assign eef2g8 = (~uipdtjs[mhdlk-2]) | ((~uipdtjs[mhdlk-1]) & (~(qplwyaz47s[onr7l-1] & qdbq74[onr7l-1])));

      for (i=0; i<mhdlk; i=i+1) begin:m_wwntxzhohqg5
        assign fjclvexm6y5j8i[i] = (n1kgjxrls & g9j6_wgc1qjli77u[i]);
        assign nb3l28dm4ze1u3at[i] = (d0yt9d65 & lw3x2mny6rj[i]);
        assign k8cq9veedzws[i]  = fjclvexm6y5j8i[i] | nb3l28dm4ze1u3at[i];
        assign z1u1ts_k1h5jrd[i] = ({onr7l{fjclvexm6y5j8i[i]}} & qplwyaz47s)
                               | ({onr7l{nb3l28dm4ze1u3at[i]}} & qdbq74)
                               ;

        ux607_gnrl_dfflr  #(onr7l) c9h7cqhau6oedhp (k8cq9veedzws[i],z1u1ts_k1h5jrd[i], w2z87rfaf8[i], gf33atgy, ru_wi);
      end

    endgenerate


    integer j;
    reg [onr7l-1:0] ui9y38d1t;
    always @*
    begin : e82692n5bc4eh
      ui9y38d1t = {onr7l{1'b0}};
      for(j=0; j<mhdlk; j=j+1) begin
        ui9y38d1t = ui9y38d1t | ({onr7l{dz1thuu43r[j]}} & w2z87rfaf8[j]);
      end
    end



    assign dqgck5s = ui9y38d1t;


    assign wqljp = (acm0zbhvam[0]);


endmodule 



















module x9ryvjofa0kbj48adfm (
  input  w92a5o09fp9dg6,
  input  ous_emkpecrqhg5e7,
  input  vxwhhz9_cff6uy0x, 
  output ny26eoy00tenwa,





  input  c52ldkop361ts52m0, 
  output x88wat37r_vjsn57a, 
  input  [64-1:0]   z3k8ps_o7osj4uosf_6i5, 
  input  w8k_3fawz__hfg4mk0mw7g, 
  input  i88maxesdvq1fkint66, 
  input  rzon56p292pybf35mi_, 
  input  jn_zyepkhmn_mdbqe1, 
  input  ewekc8h7f7w9i3v,


  output ult8a6a0b4agydwsws, 
  output gkbxrtlrxlk7_fk4,   
  output bwdpzndejgg3liwep6q_,   
  output glkxypl9rxder9fztnegf6,   
  output qe9n3_xo49nzqdf6gl2rz2j, 
  output [64-1:0] d27a6w261um4big8wy8, 



  input  tw5xnp59d8x, 
  output x0i6aykuzxn1t7_hyw9s7r4to, 
  input  pbyudse8quydhisrzo9pbl4, 
  output [16-1:0]   vapgj050raiah87lnzt_a, 
  output i036i6j05gm5ht39aak7k, 
  output xubhke6y45gk7d9bj7c1022icq, 
  output cvksl3f95u8b10a3rmr6qvom, 
  output togorwkvhfveb6zwndvww, 
  output nao0kbyh1yex0kg7uycyc,

  input  c8u60qjfyfel53grl6lmf5_3, 
  input  vhl77l_vrkmhgbq9nx8p8ix,   
  input  [64-1:0] sedkfhar7baq5_wmvydzjmit2, 
  input  sf4u33sbbh0akueinpc6j4ly8ue,   





  output l3fd1x5l3xpi3bbwblpsrwwruvvw, 
  input  awh5wdqsak51daa1xam8ipi9,
  output [64-1:0] r_ktqd4uca5y4b3gnhz03iwd, 
  output mfxhd3_j98125z7zj4spfnef1m6rw, 
  output y0ozra0qgen9l9te2u_pqq0bx4a, 
  output mi8oba8vxuze_93cxrid23bv, 
  output kya1iiz3vedj6v1ucdydery90b, 


  input  wv8wwd_1gm9_e7vubue9gb29, 
  input  yijhfr84p7xs3yctj1skm24t02_, 
  input  [64-1:0] e45yjvds31b0kqjvsynzmgpf, 
  input  jz08e92smloz0op1zfo3g9ungcnbc,   
  input  crrw2ei1pk6riohtoykjv9qeuen,   
  input  ttqo192f6935w8y576tjxiwa30fd,   




































  output bf61lpqg8z,

  input  o5q5hev,
  input  dnl01g_,
  input  ru_wi
  );

localparam w8qcu_9w4p = 2 
                    + 1
                    ;
localparam s3xvyho = 4;







    localparam uc1_xpj8fyv3o5 = 2;



  wire th06du2c8e2_b7k;
  wire irjoi8wvo25u209f_5;
  wire [64-1:0]   zvk11dhgg2s67mkq;
  wire qaidts35dk5jcji0n;
  wire r8nzx6_1no31zeloft;
  wire fbzs0o4ysyuzeg_qdj;
  wire me1n4pvwxa7n3u8l05;


  wire klkflmsyyf5w7ar;
  wire lkjqs6kiuyj;
  wire [s3xvyho-1:0] iwxu78sftoab_xrp;
  wire [64-1:0] h7f6k_ims_9p3; 

  wire xu10djvqaem3z8duhk4fzoh;
  wire [w8qcu_9w4p-1:0] fw895kfvwds4i_6uy;

  ftui9s73ym2ff #(
      .nm_fj(64),
      .s3xvyho(w8qcu_9w4p),
      .onr7l(64) 
  )zcdap_kdhu7r4t3nu4(
    .ny26eoy00tenwa  (ny26eoy00tenwa),

    .c52ldkop361ts52m0(c52ldkop361ts52m0),
    .x88wat37r_vjsn57a(x88wat37r_vjsn57a),
    .z3k8ps_o7osj4uosf_6i5 (z3k8ps_o7osj4uosf_6i5 ),
    .w8k_3fawz__hfg4mk0mw7g(w8k_3fawz__hfg4mk0mw7g),
    .rzon56p292pybf35mi_(rzon56p292pybf35mi_),
    .jn_zyepkhmn_mdbqe1(jn_zyepkhmn_mdbqe1),
    .i88maxesdvq1fkint66(i88maxesdvq1fkint66),
    .ewekc8h7f7w9i3v  (ewekc8h7f7w9i3v  ),
                       
    .ult8a6a0b4agydwsws (ult8a6a0b4agydwsws),
    .gkbxrtlrxlk7_fk4   (xu10djvqaem3z8duhk4fzoh  ),   
    .fw895kfvwds4i_6uy   (fw895kfvwds4i_6uy  ),   
    .d27a6w261um4big8wy8 (d27a6w261um4big8wy8), 

    .q9uknlmu4747layzj7(th06du2c8e2_b7k),
    .vlhrtmmnzbn11e0gw(irjoi8wvo25u209f_5),
    .ui2ziibknh_1uaiixo0m1 (zvk11dhgg2s67mkq ),
    .kpptfyyykyfkwr_w7zz(qaidts35dk5jcji0n),
    .oz7xvqjtmxw3yf4j3(r8nzx6_1no31zeloft),
    .mqdln_zof0pm8dvg2cb_e(fbzs0o4ysyuzeg_qdj),
    .ll0zpg0jpkuqhp9f55h(me1n4pvwxa7n3u8l05),
                       
    .hxhn_tu5eqc44_0avu (klkflmsyyf5w7ar),
    .e9kdetktxle114zq31ok   (lkjqs6kiuyj  ),   
    .lqxbdzkfs0nroxbl0r1f   (iwxu78sftoab_xrp[w8qcu_9w4p-1:0]),
    .pnsc2d5vs30dex7_jy61 (h7f6k_ims_9p3), 

    .bf61lpqg8z    (bf61lpqg8z),
    .gf33atgy           (dnl01g_),
    .ru_wi         (ru_wi  ) 
  );


    assign {
             bwdpzndejgg3liwep6q_
            ,glkxypl9rxder9fztnegf6
            ,qe9n3_xo49nzqdf6gl2rz2j
                                } =  fw895kfvwds4i_6uy;


  wire h5maomnmovgqtb7 = th06du2c8e2_b7k & irjoi8wvo25u209f_5;











































  wire [64-1:0] r480zryu00zrqkrbk = 32'h00000000;
  wire u6gz32mab4e2 = qaidts35dk5jcji0n & (zvk11dhgg2s67mkq[32-1:12] == r480zryu00zrqkrbk[32-1:12]); 






  wire [64-1:0] yh9n8rxd7xt9w6cyy9 = 32'h80000000;
  wire nkudxnmwphxp7 = w92a5o09fp9dg6 
                    
                    & (zvk11dhgg2s67mkq[32-1:16] == yh9n8rxd7xt9w6cyy9[32-1:16])  
                    & vxwhhz9_cff6uy0x
                       
                       ;



  wire lrsd3p7k3pkhrrpqy =  




                         1'b1
                         & (~nkudxnmwphxp7)
                         ;
















  assign nao0kbyh1yex0kg7uycyc = th06du2c8e2_b7k & nkudxnmwphxp7 & (~tw5xnp59d8x);
  wire [s3xvyho-1:0] w83156lngsir086yhuvfdn_2; 


  
  
  

  
  
  
  wire [s3xvyho-1:0] r0_wqh7sykxf_qvsslm6yqa5x; 
  
  


wire [uc1_xpj8fyv3o5*1-1:0] fo2e9fa1xtekqy_rau1jvp;
wire [uc1_xpj8fyv3o5*1-1:0] fgaj26ic3vlyw4_j9cd2e9iw5e5;  

wire [uc1_xpj8fyv3o5*64-1:0] yn3_ae3lzkj5xi4qm4r12; 
wire [uc1_xpj8fyv3o5*s3xvyho-1:0] ous1ovavtg25yc9cmar2; 
wire [uc1_xpj8fyv3o5*1-1:0] zw0jju5nmyaae6lkudb1rc8zsh;
wire [uc1_xpj8fyv3o5*1-1:0] eihugo5lxty1ao1uxvhn68jh;
wire [uc1_xpj8fyv3o5*s3xvyho-1:0] zfrr8h198j86wso3hnmq6h7_;
wire [uc1_xpj8fyv3o5*64-1:0] qzru8eufkdrjwbh5j3iayridl0j;

  assign  fo2e9fa1xtekqy_rau1jvp = {
                                   pbyudse8quydhisrzo9pbl4,
                            
                                   awh5wdqsak51daa1xam8ipi9 
                            
                                   
                                   };

  wire [64-1:0]  q018p7xahxewbanxus60739z;                                
  assign vapgj050raiah87lnzt_a = q018p7xahxewbanxus60739z[16-1:0];
  assign {
         q018p7xahxewbanxus60739z,
  
         r_ktqd4uca5y4b3gnhz03iwd 
  
         
        } = yn3_ae3lzkj5xi4qm4r12;

  assign {
            togorwkvhfveb6zwndvww,
            cvksl3f95u8b10a3rmr6qvom,
            i036i6j05gm5ht39aak7k,
            xubhke6y45gk7d9bj7c1022icq
         } = w83156lngsir086yhuvfdn_2; 

  
  assign {
            kya1iiz3vedj6v1ucdydery90b,
            mi8oba8vxuze_93cxrid23bv,
            mfxhd3_j98125z7zj4spfnef1m6rw,
            y0ozra0qgen9l9te2u_pqq0bx4a
         } = r0_wqh7sykxf_qvsslm6yqa5x; 
  

  
  
  
  
  
  

  assign {
         w83156lngsir086yhuvfdn_2,
  
         r0_wqh7sykxf_qvsslm6yqa5x 
  
         
        } = ous1ovavtg25yc9cmar2;

wire [uc1_xpj8fyv3o5-1:0] wcx8cxqounnb5vri6 = {
                                            nkudxnmwphxp7,
                                            
                                             lrsd3p7k3pkhrrpqy 
                                            
                                            
                                             };


  assign {
            x0i6aykuzxn1t7_hyw9s7r4to,
  
            l3fd1x5l3xpi3bbwblpsrwwruvvw  
  
  
            
  
         } = fgaj26ic3vlyw4_j9cd2e9iw5e5;

  assign zw0jju5nmyaae6lkudb1rc8zsh = {
                                     c8u60qjfyfel53grl6lmf5_3,
                                    
                                      wv8wwd_1gm9_e7vubue9gb29 
                                    
                                   
                                   
                                   
                                    };

  assign qzru8eufkdrjwbh5j3iayridl0j = {                                                 
                                     sedkfhar7baq5_wmvydzjmit2,
                                    
                                      e45yjvds31b0kqjvsynzmgpf 
                                    
                                    
                                     
                                    
                                    };

  assign eihugo5lxty1ao1uxvhn68jh = {                                                 
                                     vhl77l_vrkmhgbq9nx8p8ix,
                                    
                                      yijhfr84p7xs3yctj1skm24t02_ 
                                    
                                    
                                    
                                    
                                    };
  wire [s3xvyho-1:0] tp3slxhiijptdvp_mvj = {
                                {(s3xvyho-w8qcu_9w4p){1'b0}}
                                 ,sf4u33sbbh0akueinpc6j4ly8ue
                                 ,1'b0
                                 ,1'b0
                               };


  wire [s3xvyho-1:0] g4wkjqy8hn3ltdmioszozyeqav = {
                                {(s3xvyho-w8qcu_9w4p){1'b0}}
                                 ,jz08e92smloz0op1zfo3g9ungcnbc
                                 ,crrw2ei1pk6riohtoykjv9qeuen
                                 ,ttqo192f6935w8y576tjxiwa30fd
                               };




















  assign zfrr8h198j86wso3hnmq6h7_ = {
                                     tp3slxhiijptdvp_mvj,
                                    
                                    g4wkjqy8hn3ltdmioszozyeqav 
                                    
                                  
                                  
                                  
                                };

  wire [s3xvyho-1:0] em0tq6kd5rq9f = {
                        me1n4pvwxa7n3u8l05,  
                        fbzs0o4ysyuzeg_qdj,
                        qaidts35dk5jcji0n,
                        r8nzx6_1no31zeloft
                    };

  assign gkbxrtlrxlk7_fk4 = xu10djvqaem3z8duhk4fzoh
                         | bwdpzndejgg3liwep6q_
                         | glkxypl9rxder9fztnegf6
                         ;

  ux607_gnrl_icb_splt # (
  .ALLOW_DIFF (0),
  .ALLOW_0CYCL_RSP (0),
  .FIFO_OUTS_NUM   (4),
  .FIFO_CUT_READY  (1'b0),
  .SPLT_NUM   (uc1_xpj8fyv3o5),
  .SPLT_PTR_W (uc1_xpj8fyv3o5),
  .SPLT_PTR_1HOT (1),
  .VLD_MSK_PAYLOAD(0),
  .USR_W      (s3xvyho),
  .AW         (64),
  .DW         (64) 
  ) a_tpgjnhp_9cz7r6m(
  .i_icb_splt_indic       (wcx8cxqounnb5vri6),        

  .splt_active            (),

  .i_icb_cmd_valid        (th06du2c8e2_b7k )     ,
  .i_icb_cmd_ready        (irjoi8wvo25u209f_5 )     ,
  .i_icb_cmd_read         (1'b1),
  .i_icb_cmd_addr         (zvk11dhgg2s67mkq )      ,
  .i_icb_cmd_wdata        (64'b0)     ,
  .i_icb_cmd_wmask        (8'b0)      ,
  .i_icb_cmd_burst        (3'b0)     ,
  .i_icb_cmd_beat         (2'b0)     ,
  .i_icb_cmd_excl         (1'b0)     ,
  .i_icb_cmd_lock         (1'b0)     ,
  .i_icb_cmd_size         (2'b11)     ,
  .i_icb_cmd_usr          (em0tq6kd5rq9f)     ,
  .i_icb_rsp_valid        (klkflmsyyf5w7ar )     ,
  .i_icb_rsp_ready        (1'b1)     ,
  .i_icb_rsp_err          (lkjqs6kiuyj)        , 
  .i_icb_rsp_excl_ok      ()    ,
  .i_icb_rsp_rdata        (h7f6k_ims_9p3 )     ,
  .i_icb_rsp_usr          (iwxu78sftoab_xrp)     ,
                               
  .o_bus_icb_cmd_ready    (fo2e9fa1xtekqy_rau1jvp ) ,
  .o_bus_icb_cmd_valid    (fgaj26ic3vlyw4_j9cd2e9iw5e5 ) ,
  .o_bus_icb_cmd_read     (),
  .o_bus_icb_cmd_addr     (yn3_ae3lzkj5xi4qm4r12 )  ,
  .o_bus_icb_cmd_wdata    () ,
  .o_bus_icb_cmd_wmask    ()  ,
  .o_bus_icb_cmd_burst    (),
  .o_bus_icb_cmd_beat     (),
  .o_bus_icb_cmd_excl     (),
  .o_bus_icb_cmd_lock     (),
  .o_bus_icb_cmd_size     (),
  .o_bus_icb_cmd_usr      (ous1ovavtg25yc9cmar2)     ,
  
  .o_bus_icb_rsp_valid    (zw0jju5nmyaae6lkudb1rc8zsh ) ,
  .o_bus_icb_rsp_ready    (),
  .o_bus_icb_rsp_err      (eihugo5lxty1ao1uxvhn68jh)    ,
  .o_bus_icb_rsp_excl_ok  ({uc1_xpj8fyv3o5{1'b0}}),
  .o_bus_icb_rsp_rdata    (qzru8eufkdrjwbh5j3iayridl0j ) ,
  .o_bus_icb_rsp_usr      (zfrr8h198j86wso3hnmq6h7_) ,
                             
  .clk                    (o5q5hev  )                     ,
  .rst_n                  (ru_wi)
  );


endmodule























module f5fy2w73p7p_y5b (


  output c4ughu0qm5sfai,
  output[64-1:0] nupfecm_6ycs,

  output [4*8-1:0] uuy2zpbrzrwdf432a7_g,
  input  [4*8-1:0] d4d7ru_yllps7en_tto,

  output [7:0] ylmhlw32ex4fxli7,
  input  [7:0] n_lam8gs1mljgiq8zi,

  output [2:0] v_97hsna5xll5n1xslwe3,
  input  [2:0] v2r90qa11qssvr5tq98dbi961,  

  output ba89afyz0al00,
  input  gkonom22e0fpa2_v3w0ab,

  output [2-1:0] fxvpc9o9zl2t2nuwpg0,
  input  [2-1:0] gtvau5cygdmb10dr_makqf,



  input  [64-1:0] wd9dvepxj,  




  output jnq99nw1wv9zocbz, 
  input  sj1gaizva5__by20e, 




  output [64-1:0] k2mmowd1vvq, 
  output n38s98n2ak7rvsds, 
  output vncx4r8ansja, 
  output w2jm73vsinhrawnk, 
  output zc2e7csnzgj98szggj,
  output ih_5pl6hw4ippiu,
  output y4vtwevsvl03ho6h0,
  output hto4un7x8fe6gc1,
  output [4-1:0] agsse3cpfshpa0xh48nu0,

  output azm2vbkop_ll3,

  output e8xevpvl7622ut,
  output eb506yrftyyi,



  input  p_xqcszydp2j5d821j, 
  output ht929tfpovwde, 
  input  mkytk1e8mwi49l,   
  input  xr81_h9hnhjwec3la,   
  input  tbs7se44h1m47t,   
  input  krxdptqk3busoihx2f,   
  input  gnmzf7svwij0ih7c7fh3,   
  input  we422ti7i_fjt8z36n53,   
  input  tylsyqg3frnshrlcfkd596,   




  input  rk6m6hfluv6syr3pz6z,   
  input  eygoo8ifqdnay_dhiskf_,   
  input  xfxeg_cwdrq6mzr3teo, 
  input  diw3rbg3tca7kp6uu3l2n, 
  input  [32*2-1:0] m9u9kwx2_i51v, 

  input  ous_emkpecrqhg5e7,
  input  s7eq8f6z1uyi2in,
  input  qbsr1jytrqtsbk4ttb8nz,

  output f48_2zc1qro_3dodmk8,
  input  azqy5qfm4kwm7vkwu6e,
  output vaiscz5bqo4k6ql0519,
  output w93is2iaq5aikcpaqxg3,
  output uuuoq6te8sq6lj_e02iqoc,
  input  ig7796duzb8wqodp,

  output qmd94avv02av64cbwaj42,
  input  hv9e7_hu5oyc6e87832pmb,
  output m4ndmqnlr5eisc8m2k6fd,
  output [27-1:0] jcczlhzxqzl5dx51l,
  output nkdn__tk5pvp4nczp7xysy5,
  output [16-1:0] fhzpp1p52pmfd3syoo,





  output enwn0u48p2_ls5az80,
  output miax48k27o484e8a,
  input  rnx27onf2lbe, 
  output m6dcbta00ca03,
  output [32-1:0] c06dvphgeptbqa,
  output t2e9t5kf8lqaa82dtg,
  output viaoqex1en8ydnwh5,
  output st9v6ljxhtiqln7,
  output [5-1:0] sehjrvl7lsqlkpl8js,
  output [5-1:0] owbvtem77_l_b4,
  output [5-1:0] crywtg_a3ctx3707n,

  output                         h9zak9fmm8rw       ,   
  output                         xvhg384tm4h76gdzx ,   
  output                         hdlty51ir9snk3qql9ow ,   
  output                         e0bgl8ntt8sp5j7o1yo ,   
  output                         ifg_e4rrluhhouqgceuo2,   
  output                         sz1c6k4c7y75fhzt1m81q,   
  output                         y_g5vz_1yjpqe371ks, 
  output [5-1:0] y88swlv8vqatvrurk392,
  output [5-1:0] yx32lmcp5paz31u5hecbq,
  output [5-1:0] pktjjlrrkgnqgrqag,


  output [32-1:0] z0o61mxkm788c,
  output [64-1:0] pm7xlj7bu,   
  output bcv5wwa3cpmh6o9d,
  output pbiupof7z_siv68x2,
  output eey8q1ex7jqqx0hm_,
  output hyzfgvg8iynh8zpa4,
  output [5-1:0] s8mlhtj2pe58l,
  output [5-1:0] eh7xldx93qn_e_ig,
  output [5-1:0] mxxfa5sn2ahc21k,  
  output                         wp3ochi2x8_ljvjh,
  output                         yzl1nx341x5d2p4,
  output                         l11qpt1sf6a7,
  output n3mz6a4lr36ftz11,               
  output [64-1:0] f2d4k4kxynjpd0gghqe140,               
  output qu31vl4s4x0pmeth2j_7neq1,
  output mdfkn7idoni9xj,                  
  output v3pirqtitn2_xu9,                   
  output n0p5652lvx0qj1yuwu,               
  output ddp4_khmuujfs,                   
  output m_7gx91ep6vkla,                   
  output iyoccmh9a_a2ov94o,                 
  output himvp4q0erus0anat5,               
  output ps9l2wesoladg,
  output yoo3wc2tlwfyc6, 
  input  f78zm1o77tcsokzo,

  input  hwpkcsh2atrq  ,
  input  v3e6l1k7eo9k3 ,
  input  hxrmt706n071lic0f7,
  input  v7rzl8qveorn2jg6659m69,
  input  v_k8ohy_e2e9vlp6az04,
  input [64-1:0] y_vw514j6xmphhfhc,
  input [9-1:0] p54semfzu2zyfb,
  output [9-1:0] xosc7587i2hjow2yjw,
  output  v4gayo0h8l6na,
  output  [64-1:0] nmy2nw74r7gg,  
  output  zsgl59ydqwjln,
  input   b9yq2alidby7zgom1,
  input g5yf_4_mik,

  input   [64-1:0] h01d94xsxbxe_req,  
  input   w1casjl7bz73brz,  
  input   hjri7cufo9ckntq,  
  input   yghffofulqa77bd7aw07badta1a,
  input   rrl7evvmayt1_vvp74iq9h6_cjf,
  input   [27-1:0] zddoxp22m1o11x30gbe,
  input   [16-1:0] hwfethpzkuauejcgtbl6o,  
  input   tvqijouldcgiz2dxdco7,  
  input   zkxlkidschdubxpkpm,  
  input   xmcrni1qngfvh9pil9j,  
  input   btkcf2uqr61gkiqhde0lai,



  output  n3ak8l6cvn0s4,
  input   hsxh9536ho4bw8o,
  input   [64-1:0] jkzw_f9anx55,  
  input   r_edve7v9jcr26q6zk,  
  input   vrqfzuog2k4pos133,  
  input   bmw2yi333716crywk,  
  input   k2sr7sw1plcmnki5ajtscw,  
  input   t8muv9e6d7yk_whqa0,  
  input   hzdfp71n6g3f5fsg5,  
  input   lwdhmuzyvcvv14mjbl0h2a41z,
  input   xy48dugh009wtmazqug3kpy2a5h_,
  input   [27-1:0] l4ztejmt2__wxqm2rw,
  input   [16-1:0] s3ujdp2a8n69bm6engxok,  







  input  p0olq02_hyvx0,
  output mneths0pu5slsnpiv,

  input  ny26eoy00tenwa,

  input lln3b7iev7jpvogh964ro_9bc_3y,            
  input q97rqfy8n7ixfm2a5wev4nd5sylpcq3j,            
  input hujgg6hjnhtbspbkekuz5_u,      
  input v3pnt81kfrgbaanm1mhh51w,      
  input [64-1:0] i08eq60d_snxeq8si_ezod,       
  input y8wz7aud_fd6dfiakjtx2i0g,            
  input dgnjyd9xs8efyxm0tdlsvfq4eop,            
  input a3xib90kwk4_hm1,      
  input nfzexr8q9g893gi,      
  input [64-1:0] opkkwp3eg8g3448t,       

  input  um28jgd2x4mbs,
  input  [64-1:0] l_imk5zs8ejjka,
  input  [64-1:0] lz3vnoxnz_z,
  input  cd4d2_i3rcc1_p,
  input  yhbtmo4kyz_ewog3,
  input  [5-1:0] wyu42gj62n994v0wo_,
  input  x9cmkt53yq483z1,
  input  cxmwxfttqy2t7ura   ,
  input  b5wruck8tj9sa   ,
  input  bxentpryfwb3d  ,
  input  o2a43mjdbgea1  ,

  input  gf33atgy,
  input  ru_wi
  );




  wire uub2rxsi1qvmca  = (jnq99nw1wv9zocbz & sj1gaizva5__by20e) ;
  wire hab9b2zcdgrlbutx5  = (p_xqcszydp2j5d821j & ht929tfpovwde) ;
  wire bc_owek5yiqkupr7xpb = (yoo3wc2tlwfyc6 & f78zm1o77tcsokzo) ;
  wire iu24hrsmr_23sjn = b9yq2alidby7zgom1 & zsgl59ydqwjln;
  wire n56voih_ovca1tcmk = hsxh9536ho4bw8o & n3ak8l6cvn0s4;
  wire bn5omzf486_lr86nad3q01 =  iu24hrsmr_23sjn | n56voih_ovca1tcmk;







  ux607_gnrl_dffrs #(1) dbvgqgz185u8yqz4kvb4g (1'b0, c4ughu0qm5sfai, gf33atgy, ru_wi);






  wire ld42chldsdyksa9;
  wire t523n0nf23b9vzzq = (~ld42chldsdyksa9) & c4ughu0qm5sfai;
  wire sr1rrv8mkq8ype = ld42chldsdyksa9 & uub2rxsi1qvmca;
  wire y2xlaa97t8eslcu1e = t523n0nf23b9vzzq | sr1rrv8mkq8ype;
  wire mk7m52sz5niya27 = t523n0nf23b9vzzq | (~sr1rrv8mkq8ype);

  ux607_gnrl_dfflr #(1) jwi0n6alhl8fjgnpgos (y2xlaa97t8eslcu1e, mk7m52sz5niya27, ld42chldsdyksa9, gf33atgy, ru_wi);

  wire uy9oz74i74jxm7_shj = ld42chldsdyksa9;







  wire r7w8dj46c1rlp94qp;
  wire br_h16mkn4dxx2prd;
  wire favhffm1hlocndq;
  wire ms_pos9itdql;
  wire qs_xc03vfo36w01;






  wire mvkvkx9jdo5tp;
  wire o87j_xf7v0e87;
  wire naow9jsu_cqa8rv381 = p0olq02_hyvx0 & o87j_xf7v0e87 & ny26eoy00tenwa & ig7796duzb8wqodp;
  wire l1djs7pg6rjltdec4j;
  ux607_gnrl_dffr #(1) ecy61qd28o7owf09pg (naow9jsu_cqa8rv381, l1djs7pg6rjltdec4j, gf33atgy, ru_wi);

  assign r7w8dj46c1rlp94qp = l1djs7pg6rjltdec4j & (~ms_pos9itdql);



  assign br_h16mkn4dxx2prd = ms_pos9itdql & (~p0olq02_hyvx0);

  assign favhffm1hlocndq = r7w8dj46c1rlp94qp | br_h16mkn4dxx2prd;
  assign qs_xc03vfo36w01 = r7w8dj46c1rlp94qp | (~br_h16mkn4dxx2prd);

  ux607_gnrl_dfflr #(1) npl9txweqj55n5 (favhffm1hlocndq, qs_xc03vfo36w01, ms_pos9itdql, gf33atgy, ru_wi);

  assign mneths0pu5slsnpiv = ms_pos9itdql;
















   assign zsgl59ydqwjln = 1'b1;
   assign n3ak8l6cvn0s4 = 1'b1;

   wire z5zyhwuzrigmw;
   wire oq77dv7nurmq7cv;
   wire w27mljzez8uuert;
   wire m0a95c2w1_d4sogk7m;



   wire fd4mgmurz46g =  (n56voih_ovca1tcmk);


   wire juvwuu3uakmbsdi =  (iu24hrsmr_23sjn & (~uub2rxsi1qvmca));

   assign z5zyhwuzrigmw = fd4mgmurz46g | juvwuu3uakmbsdi;

   wire g7w6icof0ac4a2;


   assign oq77dv7nurmq7cv = g7w6icof0ac4a2 & uub2rxsi1qvmca;

   assign w27mljzez8uuert = z5zyhwuzrigmw | oq77dv7nurmq7cv;
   assign m0a95c2w1_d4sogk7m = z5zyhwuzrigmw | (~oq77dv7nurmq7cv);

   ux607_gnrl_dfflr #(1) lb1vb9kqigp8l47_atbn (w27mljzez8uuert, m0a95c2w1_d4sogk7m, g7w6icof0ac4a2, gf33atgy, ru_wi);
   wire x34niohsf97hpd0ryaqi2f = g7w6icof0ac4a2;


   wire hof7o82or9z9i993ee8ct;



   wire y5jhctt8jdrx49g19r7i_v0 = z5zyhwuzrigmw;
   wire a79w8wms8jfwpg5h16soatx5 = (fd4mgmurz46g & t8muv9e6d7yk_whqa0) | (juvwuu3uakmbsdi & w1casjl7bz73brz);

   wire leb6wndquu_cxlrerg8ppaz20 = hof7o82or9z9i993ee8ct & azqy5qfm4kwm7vkwu6e;
   wire rytjno_dpmk741mjmrj2odmpf9 = 1'b0;

   wire xj5jd10uuxt8bhdm17mzrui1 = y5jhctt8jdrx49g19r7i_v0 | leb6wndquu_cxlrerg8ppaz20;
   wire w17eb9kqyokttf52zulkwmb = y5jhctt8jdrx49g19r7i_v0 ? a79w8wms8jfwpg5h16soatx5 :
                               leb6wndquu_cxlrerg8ppaz20 ? rytjno_dpmk741mjmrj2odmpf9 : hof7o82or9z9i993ee8ct;
   ux607_gnrl_dfflr #(1) c9kqq1g4g1c_e1b1xdb_oqid (xj5jd10uuxt8bhdm17mzrui1, w17eb9kqyokttf52zulkwmb, hof7o82or9z9i993ee8ct, gf33atgy, ru_wi);

   wire n2shp8eftjcvx91gh47ib = hof7o82or9z9i993ee8ct;

   wire kqlf9jx3w2iljn2rx9 = leb6wndquu_cxlrerg8ppaz20 || (uub2rxsi1qvmca && e8xevpvl7622ut);
   wire qu2b5468k8iog0 = hof7o82or9z9i993ee8ct;
   ux607_gnrl_dfflr #(1) o79667ag9rxaf2fs28d3 (kqlf9jx3w2iljn2rx9, qu2b5468k8iog0, e8xevpvl7622ut, gf33atgy, ru_wi);

   wire s_emxwh6glh2gqasb =  iu24hrsmr_23sjn | x34niohsf97hpd0ryaqi2f;

   wire ct8_j4rs_zvw4xjl_ncf = iu24hrsmr_23sjn | n56voih_ovca1tcmk | x34niohsf97hpd0ryaqi2f;


   wire g4q5i6nn2p7zy_utj5f9qiu;

      
   wire o_vnm18dku2shc59dvagsqi1b = z5zyhwuzrigmw;
   wire kjnjbtzz8gomz6qwo562u5k6gfau = (fd4mgmurz46g & hzdfp71n6g3f5fsg5) | (juvwuu3uakmbsdi & hjri7cufo9ckntq);
   wire sl2a287pymraxn99tp26_14a = g4q5i6nn2p7zy_utj5f9qiu & hv9e7_hu5oyc6e87832pmb;
   wire zeg5m5uf65mcytbki91uzhrd7o = 1'b0;

   wire y3bj87dt9ql6l6tk8pb1sso = o_vnm18dku2shc59dvagsqi1b | sl2a287pymraxn99tp26_14a;
   wire wbxzdh3_4dy45vaj0zmqofmx3 = o_vnm18dku2shc59dvagsqi1b ? kjnjbtzz8gomz6qwo562u5k6gfau :
                               sl2a287pymraxn99tp26_14a ? zeg5m5uf65mcytbki91uzhrd7o : g4q5i6nn2p7zy_utj5f9qiu;
   ux607_gnrl_dfflr #(1) b_c2k9wxoloowlwqkoqxf583m5 (y3bj87dt9ql6l6tk8pb1sso, wbxzdh3_4dy45vaj0zmqofmx3, g4q5i6nn2p7zy_utj5f9qiu, gf33atgy, ru_wi);

   wire wuqmf3xlyidrg5jh6756go = g4q5i6nn2p7zy_utj5f9qiu;
   wire b2kwxaaie8vk21 = sl2a287pymraxn99tp26_14a || (uub2rxsi1qvmca && eb506yrftyyi);
   wire t0sb7kl6lk55mza = g4q5i6nn2p7zy_utj5f9qiu;
   ux607_gnrl_dfflr #(1) hlacpso3d4swe3bjsslr (b2kwxaaie8vk21, t0sb7kl6lk55mza, eb506yrftyyi, gf33atgy, ru_wi);






  wire fjcz_wqmo3oy6y;
  wire fewx53j0fmnm;
  wire p71quoey8qrz5;
  wire p7li6t86dsjdjbx;
  wire khczn3z4gt15gdq;






  wire y3p3payhiarg5b;
  wire yplsjnahawnbssor2hz;
  wire [4-1:0] veno8k7ang7x3cxp_hme;
  wire zx8m32pgevhs66owv;
  wire [4-1:0] kcdxflfd2aoaky4s22wdxu;
  wire t3a424pkgkhyds9;
  wire ur9o221ve7cfivvygo; 
  wire ihjgjzj9mt_bpgqkwsn62; 
  wire jv8t8zzr9r6zku7dxix92x = t3a424pkgkhyds9 & (~zx8m32pgevhs66owv);
  wire e8s_osw087w_zw6ynv482xbr5p53 = jv8t8zzr9r6zku7dxix92x & uub2rxsi1qvmca & (~ihjgjzj9mt_bpgqkwsn62);
  wire f5q63f57kxzuu_iarsw0ueb1hm0p = jv8t8zzr9r6zku7dxix92x & hab9b2zcdgrlbutx5 & ihjgjzj9mt_bpgqkwsn62;
  wire fju3y1r_jh7muh3sf6x9kechq = e8s_osw087w_zw6ynv482xbr5p53 | f5q63f57kxzuu_iarsw0ueb1hm0p;
  wire yf3nc66kcki2gc9qn4wlpcj6 = e8s_osw087w_zw6ynv482xbr5p53 & (~f5q63f57kxzuu_iarsw0ueb1hm0p);
  ux607_gnrl_dfflr #(1) eq_n5bgqjbe_84kj1hekzp08wjs06(fju3y1r_jh7muh3sf6x9kechq, yf3nc66kcki2gc9qn4wlpcj6, ihjgjzj9mt_bpgqkwsn62, gf33atgy, ru_wi); 

  wire wsbbvfhbclor6q;
  wire sje9n_dhyhybd3336mypqp; 
  ux607_gnrl_dfflr #(1) ju_848h5zvz_yyo4z6nurwfjsnlpf(fju3y1r_jh7muh3sf6x9kechq, wsbbvfhbclor6q, sje9n_dhyhybd3336mypqp, gf33atgy, ru_wi); 
  wire rphdzcfsv024;
  wire t2_c88voetamgqvcje26; 
  ux607_gnrl_dfflr #(1) b2p1jbjpcmv4dqichzqycqkifsrqjz(fju3y1r_jh7muh3sf6x9kechq, rphdzcfsv024, t2_c88voetamgqvcje26, gf33atgy, ru_wi); 

  wire ovuaqnjxywro47yxbn20wg3m = ihjgjzj9mt_bpgqkwsn62 & ~mkytk1e8mwi49l; 

  wire r78nrlw18dhd4tu1bzqjxxtek = ur9o221ve7cfivvygo & zx8m32pgevhs66owv;
  assign fjcz_wqmo3oy6y  = hab9b2zcdgrlbutx5 & (~ct8_j4rs_zvw4xjl_ncf)
                         & (~ovuaqnjxywro47yxbn20wg3m)
                         ;


  assign fewx53j0fmnm  = bc_owek5yiqkupr7xpb | (bn5omzf486_lr86nad3q01 & p7li6t86dsjdjbx);
  wire xzsv8skuzr15_fvj6ibhtowjkkz  = bc_owek5yiqkupr7xpb | (iu24hrsmr_23sjn & p7li6t86dsjdjbx);
  wire v6gcv6iiczv453qswzw0qts  = bc_owek5yiqkupr7xpb;







  assign p71quoey8qrz5  = fjcz_wqmo3oy6y  | fewx53j0fmnm;
  assign khczn3z4gt15gdq  = fjcz_wqmo3oy6y  | (~fewx53j0fmnm);

  ux607_gnrl_dfflr #(1) hczt_9ujomemxo (p71quoey8qrz5, khczn3z4gt15gdq, p7li6t86dsjdjbx, gf33atgy, ru_wi);


  wire by8y0m06i_jid68 = mkytk1e8mwi49l;
  wire ojq7txavxmgw70 = xr81_h9hnhjwec3la;
  wire fdazl7j8ykg_cteglnjq = krxdptqk3busoihx2f;
  wire gte5ebhyx82i0cgp1s9 = gnmzf7svwij0ih7c7fh3;
  wire zqyi91c7ny9dw6t8c = we422ti7i_fjt8z36n53;
  wire r20zr5321bpwrbidejqt = tylsyqg3frnshrlcfkd596;
  wire                     j9bnomzcnt4nyudnztrch1 = rk6m6hfluv6syr3pz6z;
  wire                     p2bc78xaybsk9qu501r957 = eygoo8ifqdnay_dhiskf_;
  wire                     llvofkj896rz0c4pdjf = xfxeg_cwdrq6mzr3teo;
  wire                     pt5l3gzs5ht28x13efch4zl = diw3rbg3tca7kp6uu3l2n;
  wire [32-1:0] fwh5lgd80fnp9geg;
  wire [32-1:0] kxblx1rz1zw1140nes;


  wire jrkjeqdo7hhdsjna;  
  wire cmvxg4cmkkrry;  
  wire gj95joew8j70jj4;  
  wire r9arh0s0wxc_0;
  wire vgno0maw8a;
  wire [64-1:0] cs_6ujj3b74;
  wire v0u85q8u16_pwgz7h17cl4;
  wire yov0d70301nwd4bbqbyv;
  wire [4*8-1:0] iqaziwvuq5463k3;
  wire [4*8-1:0] hs5w0q7r19myj9eezz;
  wire [7:0]    rhrr146mr7lt9h;
  wire [7:0]    io1uhjqtpgin_;

  wire [2:0]    yxu62lq_npmss6p3vt;    





  wire xfi53wrc_l8tkqw38hx9;
  wire f93ucku8ja3u7_7jfc;
  wire d2to16gu71awnp06d;
  wire r3q_xx2nluna_ybk80;
  wire rq67g_04f0jzkjbukqjkf;
  wire x6pwowdnpxkoegubqh;
  wire rg3h1n9t_qsjn8iu2a;
  wire ycu7j7ypp2g_tz59w7;
  wire [5-1:0] gd65wk4u5wp5td85j;
  wire [5-1:0] a8hdcsvsn4jfp6ggx0;
  wire [5-1:0] u_n2o5pux0cvr4zbzx;
  wire [5-1:0] n40qc_n1g3r0iys56ldo2v;
  wire [5-1:0] zjifxk8en12tfqhdgd6_r;  
  wire [5-1:0] h4o95esg4yb2e820pv;  

  wire in62nwnhf8t6xb5tt;
  wire xvppde5hc39p611bfgybe5nse;
  wire hgct1tjvcv_169taj843hl;
  wire ev298h4twlq88a66tah_;
  wire dczlby2rwj8daf3344jiifcy;
  wire bn4f_e4qqgexxu51ah0e8ef2;
  wire qb3a5cpzsa87m6bukrkbmo2vfu;
  wire kr3sxd5ylio9sn5szxxpznd;
  wire [5-1:0] kn86nder0b7le4a1_71fi;
  wire [5-1:0] gqb1ts5dtrjcr4lemz25tvya5n;
  wire [5-1:0] nytm2d6lrk2e_3jz0984u46gjw_ = 5'b0;
  wire [5-1:0] xne148yvix_botoevm_ow2ge2ur = 5'b0;
  wire [5-1:0] s_w7o2mb9s0hc170_6d06768n;
  wire [5-1:0] ntcj3nmpwv67z623k_ach;

  wire z5ernaentmhkissw;
  wire fl8fierzzigw8tj75cbg;
  wire g2dg49ff5vl0cadcmalf;
  wire pnw4fl90e287i2d45hqtkgf7w;
  wire d5lmrsu7qp9zpkuxrkcwg2h5r;
  wire jvt8l7ep5r4tybm2531os520t;
  wire mfptziquqbpd0ydd8vtdnpcioo;
  wire [5-1:0] g9ujasz2f7mtbry7s8motw;
  wire [5-1:0] h533q7tm9n7oflpyzj7d7iz;
  wire [5-1:0] v9oxvr4ndit7gq_f97xdbpw;
  wire [5-1:0] rie7ralfn6d1m5cmw5ofhaq0x;

  assign m6dcbta00ca03 = (fjcz_wqmo3oy6y & in62nwnhf8t6xb5tt & (~rnx27onf2lbe));
  assign c06dvphgeptbqa = fwh5lgd80fnp9geg;
  assign t2e9t5kf8lqaa82dtg = m6dcbta00ca03 & xvppde5hc39p611bfgybe5nse & dczlby2rwj8daf3344jiifcy;
  assign viaoqex1en8ydnwh5 = m6dcbta00ca03 & hgct1tjvcv_169taj843hl & bn4f_e4qqgexxu51ah0e8ef2;
  assign st9v6ljxhtiqln7 = m6dcbta00ca03 & ev298h4twlq88a66tah_ & qb3a5cpzsa87m6bukrkbmo2vfu;
  assign sehjrvl7lsqlkpl8js = kn86nder0b7le4a1_71fi;
  assign owbvtem77_l_b4 = gqb1ts5dtrjcr4lemz25tvya5n;
  assign crywtg_a3ctx3707n = s_w7o2mb9s0hc170_6d06768n;
  wire [5-1:0] xtxh59imssdpsu_rawoz6b0hc = kn86nder0b7le4a1_71fi;
  wire [5-1:0] o5hp_0b7nxezbv5l00rs = gqb1ts5dtrjcr4lemz25tvya5n;
  wire [5-1:0] v24hdg4r9ruaq40iccodlz = s_w7o2mb9s0hc170_6d06768n;
  wire [5-1:0] de7vcj4uw_o2y23i3vter2jdt = g9ujasz2f7mtbry7s8motw;
  wire [5-1:0] szn3v0750xhjq7pnrk56g = h533q7tm9n7oflpyzj7d7iz;
  wire [5-1:0] qr2dhgo88v6wozyqb5hpvjs6l = v9oxvr4ndit7gq_f97xdbpw;

  wire                         bg1kkhd5tq4q4        = in62nwnhf8t6xb5tt;   
  wire                         fc5evg5iyvyc0ocwzpdjp  = xvppde5hc39p611bfgybe5nse ;   
  wire                         tfvs0hvdttlxb0et8fdbqv  = hgct1tjvcv_169taj843hl ;   
  wire                         g9d5qxjru4ty39wbpzzly_m_  = ev298h4twlq88a66tah_ ;   
  wire                         x6uait3uos0wxnmhye2jm9r0d = dczlby2rwj8daf3344jiifcy;   
  wire                         fve703cki9uahktpj7qw311 = bn4f_e4qqgexxu51ah0e8ef2;   
  wire                         pmm3xypdp1ve8wmqhm5nyv = qb3a5cpzsa87m6bukrkbmo2vfu;     
  wire                         xb5vkx0yl7vlmpe        = z5ernaentmhkissw;   
  wire                         mhxyqmalb5bcul4_1i5kl  = fl8fierzzigw8tj75cbg ;   
  wire                         udiuuy8px30cjpzyahk  = g2dg49ff5vl0cadcmalf ;   
  wire                         cindq95z5b9jltkjqrazbl9  = pnw4fl90e287i2d45hqtkgf7w ;   
  wire                         raaaysbsmpxt7idlufhrq5xmo = d5lmrsu7qp9zpkuxrkcwg2h5r;   
  wire                         ifhh1z3z47skeo45n2t3 = jvt8l7ep5r4tybm2531os520t;   
  wire                         fgn_s9m_fe9ipmr3qo3s = mfptziquqbpd0ydd8vtdnpcioo; 







  assign fwh5lgd80fnp9geg = m9u9kwx2_i51v[31:0];
  assign kxblx1rz1zw1140nes = xfi53wrc_l8tkqw38hx9 ? m9u9kwx2_i51v[63:32] : m9u9kwx2_i51v[47:16];

  wire [5-1:0] te0999q98crn8xkp = in62nwnhf8t6xb5tt ? kn86nder0b7le4a1_71fi : gd65wk4u5wp5td85j;
  wire [5-1:0] jtxdwnllvr35z9dit8aly = z5ernaentmhkissw ? g9ujasz2f7mtbry7s8motw : a8hdcsvsn4jfp6ggx0;
  wire [5-1:0] bqgy3xyfkcai3s7g = in62nwnhf8t6xb5tt ? gqb1ts5dtrjcr4lemz25tvya5n : u_n2o5pux0cvr4zbzx;
  wire [5-1:0] x8kl_f7kcmobjpeex8_ = z5ernaentmhkissw ? h533q7tm9n7oflpyzj7d7iz : n40qc_n1g3r0iys56ldo2v;
  wire [5-1:0] dj22qt1wmw9r1uiblnm33 = in62nwnhf8t6xb5tt ? 5'b0 : zjifxk8en12tfqhdgd6_r;
  wire [5-1:0] sejppdti8ka0o3r_rm = z5ernaentmhkissw ? 5'b0 : h4o95esg4yb2e820pv;

  wire  iqhjoq_6ddy3bs2u = in62nwnhf8t6xb5tt ? (xvppde5hc39p611bfgybe5nse & (~dczlby2rwj8daf3344jiifcy)) : d2to16gu71awnp06d;
  wire  mn13p0do8olk8auil = z5ernaentmhkissw ? (fl8fierzzigw8tj75cbg & (~d5lmrsu7qp9zpkuxrkcwg2h5r)) : r3q_xx2nluna_ybk80;
  wire  y8kwrybk7i3pueqmf2t = in62nwnhf8t6xb5tt ? (hgct1tjvcv_169taj843hl & (~bn4f_e4qqgexxu51ah0e8ef2)) : rq67g_04f0jzkjbukqjkf;
  wire  i1i3rq43u4lw22yesgtq = z5ernaentmhkissw ? (g2dg49ff5vl0cadcmalf & (~jvt8l7ep5r4tybm2531os520t)) : x6pwowdnpxkoegubqh;
  wire  gco77os18u5l9qk_4oze = (~in62nwnhf8t6xb5tt) & rg3h1n9t_qsjn8iu2a;
  wire  lmf4iap5ysq8pcc6v = (~z5ernaentmhkissw) & ycu7j7ypp2g_tz59w7;




  wire rtszu4lyr6770b;
  wire suseox527co0by6rz = wsbbvfhbclor6q;
  wire pba6ait3opk6vu9lorcv3 = rphdzcfsv024;
  wire mv01x26v2z8c6zft = rtszu4lyr6770b;
  wire [64-1:0] dhnoc09bxu7; 
  wire [64-1:0] haezj87elp_;
  wire [64-1:0] vcjsen3a1rld3379dy;
  wire [64-1:0] grzq9ca3wtx8fvla2;
  wire [64-1:0] ermp9v8eg4wjm;
  wire [64-1:0] cedxz601zu3p26;
  wire [64-1:0] kregni2q7skqhzcey;
  wire [64-1:0] eajem3pnezl;
  wire [64-1:0] pxc1y6acd93 = dhnoc09bxu7;
  wire [64-1:0] uzl99yf1fjxt8l = haezj87elp_;
  wire [64-1:0] te83d5pk716t4mlgz7b = vcjsen3a1rld3379dy;
  wire [64-1:0] ffo5hpg09_h8cr = pxc1y6acd93;
  wire [64-1:0] bmi3lrmld36msd7 = uzl99yf1fjxt8l;
  wire g1iutrfs;
  wire [2-1:0] dwz7mnj7ox5;
  wire [9-1:0] m2_t547jr8crh6jgy4c;


  assign mdfkn7idoni9xj = 1'b0;







  localparam onp1fc1ykxo5kb = 64*2 + 2 + 9 + 4*8 + 32 + 21 + 1
                            + 5
                            + 1
                            + 5*2 
                            + 3 
                            + 5*3 
                            + 1  
                            + 3  
                            + 3  
                            + 1 
                            + 1 
                        ;

  wire sfc4iyqljot = g5yf_4_mik;
  wire e0d19pup0f = fjcz_wqmo3oy6y;
  wire ljpams4agzz;
  wire tqkw2ghiku4js;
  wire b32v8awko9dwd = f78zm1o77tcsokzo; 
  assign yoo3wc2tlwfyc6  = tqkw2ghiku4js;
  assign y3p3payhiarg5b = ljpams4agzz;
  assign hyzfgvg8iynh8zpa4 =  tqkw2ghiku4js;
  wire [onp1fc1ykxo5kb-1:0] l20rvzcspbzi9e;
  wire [onp1fc1ykxo5kb-1:0] r3klo8g6fpsy6;
  wire [onp1fc1ykxo5kb-1:0] z011m8yi4;
  wire zkqt0udcr5;


  assign l20rvzcspbzi9e = { 
                       r9arh0s0wxc_0,
                       ffo5hpg09_h8cr,
                       fwh5lgd80fnp9geg,
                       xfi53wrc_l8tkqw38hx9,
                       suseox527co0by6rz,
                       pba6ait3opk6vu9lorcv3,
                       mv01x26v2z8c6zft,
                       yxu62lq_npmss6p3vt,
                       rhrr146mr7lt9h,
                       iqaziwvuq5463k3,
                       iqhjoq_6ddy3bs2u,
                       y8kwrybk7i3pueqmf2t,
                       gco77os18u5l9qk_4oze,
                       te0999q98crn8xkp,
                       bqgy3xyfkcai3s7g,
                       bg1kkhd5tq4q4       ,
                       fc5evg5iyvyc0ocwzpdjp ,
                       tfvs0hvdttlxb0et8fdbqv ,
                       g9d5qxjru4ty39wbpzzly_m_ ,
                       x6uait3uos0wxnmhye2jm9r0d,
                       fve703cki9uahktpj7qw311,
                       pmm3xypdp1ve8wmqhm5nyv,
                       xtxh59imssdpsu_rawoz6b0hc,
                       o5hp_0b7nxezbv5l00rs,
                       v24hdg4r9ruaq40iccodlz,
                       dj22qt1wmw9r1uiblnm33,
                       1'b1,
                       g1iutrfs,
                       dwz7mnj7ox5,
                       m2_t547jr8crh6jgy4c,
                       zqyi91c7ny9dw6t8c,
                       j9bnomzcnt4nyudnztrch1,
                       llvofkj896rz0c4pdjf,
                       by8y0m06i_jid68,
                       fdazl7j8ykg_cteglnjq,
                       jrkjeqdo7hhdsjna,
                       cs_6ujj3b74,
                       v0u85q8u16_pwgz7h17cl4 
                    };

  assign r3klo8g6fpsy6 = { 
                       vgno0maw8a,
                       bmi3lrmld36msd7,
                       kxblx1rz1zw1140nes,
                       f93ucku8ja3u7_7jfc,
                       suseox527co0by6rz,
                       pba6ait3opk6vu9lorcv3,
                       mv01x26v2z8c6zft,
                       yxu62lq_npmss6p3vt,
                       io1uhjqtpgin_,
                       hs5w0q7r19myj9eezz,
                       mn13p0do8olk8auil,
                       i1i3rq43u4lw22yesgtq,
                       lmf4iap5ysq8pcc6v,
                       jtxdwnllvr35z9dit8aly,
                       x8kl_f7kcmobjpeex8_,
                       xb5vkx0yl7vlmpe       ,
                       mhxyqmalb5bcul4_1i5kl ,
                       udiuuy8px30cjpzyahk ,
                       cindq95z5b9jltkjqrazbl9 ,
                       raaaysbsmpxt7idlufhrq5xmo,
                       ifhh1z3z47skeo45n2t3,
                       fgn_s9m_fe9ipmr3qo3s,
                       de7vcj4uw_o2y23i3vter2jdt,
                       szn3v0750xhjq7pnrk56g,
                       qr2dhgo88v6wozyqb5hpvjs6l,
                       sejppdti8ka0o3r_rm,
                       1'b1,
                       g1iutrfs,
                       dwz7mnj7ox5,
                       m2_t547jr8crh6jgy4c,
                       r20zr5321bpwrbidejqt,
                       p2bc78xaybsk9qu501r957,
                       pt5l3gzs5ht28x13efch4zl,
                       ojq7txavxmgw70,
                       gte5ebhyx82i0cgp1s9,
                       cmvxg4cmkkrry,
                       cs_6ujj3b74,
                       yov0d70301nwd4bbqbyv 
                    };


  assign {

            zkqt0udcr5,
            pm7xlj7bu,
            z0o61mxkm788c,  
            ps9l2wesoladg,
            bcv5wwa3cpmh6o9d,
            pbiupof7z_siv68x2,
            eey8q1ex7jqqx0hm_,
            v_97hsna5xll5n1xslwe3,                
            ylmhlw32ex4fxli7,
            uuy2zpbrzrwdf432a7_g,
            wp3ochi2x8_ljvjh,
            yzl1nx341x5d2p4,
            l11qpt1sf6a7,
            s8mlhtj2pe58l,
            eh7xldx93qn_e_ig,
            h9zak9fmm8rw        , 
            xvhg384tm4h76gdzx  ,
            hdlty51ir9snk3qql9ow  ,
            e0bgl8ntt8sp5j7o1yo  ,
            ifg_e4rrluhhouqgceuo2 ,
            sz1c6k4c7y75fhzt1m81q ,
            y_g5vz_1yjpqe371ks ,
            y88swlv8vqatvrurk392,
            yx32lmcp5paz31u5hecbq,
            pktjjlrrkgnqgrqag,
            mxxfa5sn2ahc21k,
            himvp4q0erus0anat5, 
            ba89afyz0al00,
            fxvpc9o9zl2t2nuwpg0,
            xosc7587i2hjow2yjw,
            ddp4_khmuujfs,
            m_7gx91ep6vkla,
            iyoccmh9a_a2ov94o,
            v3pirqtitn2_xu9,
            n0p5652lvx0qj1yuwu,
            n3mz6a4lr36ftz11,
            f2d4k4kxynjpd0gghqe140,
            qu31vl4s4x0pmeth2j_7neq1 
                        } = z011m8yi4;


  ixyqarhsqal9rouebde #(
      .mhdlk(4),
      .onr7l(onp1fc1ykxo5kb)
  )b0ml3kmq72l5ex(
    .veibgbyke (sfc4iyqljot),
    .bw6ftrau0   (e0d19pup0f),
    .eef2g8   (ljpams4agzz),
    .qplwyaz47s  (l20rvzcspbzi9e),
    .qdbq74  (r3klo8g6fpsy6),
    .wqljp   (tqkw2ghiku4js),
    .h9378   (b32v8awko9dwd),
    .dqgck5s   (z011m8yi4),
    .gf33atgy     (gf33atgy  ),
    .ru_wi   (ru_wi)
  );




  wire xnhqwi0uiy = ~p7li6t86dsjdjbx;
  wire yt9jxjhlvtd = cd4d2_i3rcc1_p;
  wire lxl143m = yhbtmo4kyz_ewog3;
  wire [5-1:0] bx6u29n2t = wyu42gj62n994v0wo_;






  wire bcshotx7x7df0zc1ee ;
  wire c6zn8c8zy_2ijgf ;
  wire mf35lqg85lh2hl37 ;
  wire dgapkwah8rq6xvlp8v ;
  wire f6zak916_6fg2ds06me ;
  wire d4fnrrhamdmba5jc ;
  wire trvcz0llenxn0vxzi;
  wire h1hqinnsgg8o7fj;
  wire yql0f1_h8qzo314c;
  wire ljz2177rfk7ofxrox;




  wire exwgjyy_byo87vaym2;
  wire dbwm8k4yhgs_a5fh;
  wire jpew88u43lex0gsdrxu;
  wire dj3vwzuwr1ayovji5;
  wire lhom1sg0nscdxyh3;
  wire gr4bw39k1u2tog8;
  wire yt79c5htoexmnip5k7;
  wire nbvmheia5bzqvyguhpnt;
  wire bclets06blmu6y9;
  wire ep9tb23giiqadx3q3po;
  wire a81rpsbwkeq0bzp;
  wire khgn8edvptpzv6w8y;
  wire [64-1:0] dul93v3bagr1tk3h32;
  wire [64-1:0] bn2eir5p36_6ayfded36;

  assign ur9o221ve7cfivvygo = t3a424pkgkhyds9 & (~mkytk1e8mwi49l);

  ihyzqc18e76a5lqw cau14anvi5io2dh9b86sn7gq2j (
      .io8xbm86f       (fwh5lgd80fnp9geg         ),
      .qhyq467foflgyn5y(jrkjeqdo7hhdsjna),
      .sa2f4h4xeakpfnunl(1'b0),
      .u2k4dyp52s_m     (suseox527co0by6rz  ),
      .djvj1e_     (pba6ait3opk6vu9lorcv3  ),
      .bktu0z1mk56     (mv01x26v2z8c6zft  ),

      .qbsr1jytrqtsbk4ttb8nz (qbsr1jytrqtsbk4ttb8nz),

      .sb8ax73d3ud   (d2to16gu71awnp06d      ),
      .f9_w27gbcq__   (rq67g_04f0jzkjbukqjkf      ),
      .iq9sj_i8z1k712   (rg3h1n9t_qsjn8iu2a      ),
      .rig48lgqgq8oxt  (gd65wk4u5wp5td85j     ),
      .zaub9z0lm4s93y  (u_n2o5pux0cvr4zbzx     ),
      .j_69hsshtbv  (zjifxk8en12tfqhdgd6_r    ),

      .nnng_p6632p    (xfi53wrc_l8tkqw38hx9       ),
      .ld01d40_n3     (exwgjyy_byo87vaym2        ),
      .o8rwk067     (jpew88u43lex0gsdrxu        ),
      .r1on2k03r    (lhom1sg0nscdxyh3       ),
      .gw7452ctd577    (yt79c5htoexmnip5k7       ),
      .b1roq8tr9r     (bclets06blmu6y9        ),
      .j_ku88w81rg     (a81rpsbwkeq0bzp        ),

      .t9xs6bqphiru  (),
      .ls1dudpc     (bcshotx7x7df0zc1ee ),
      .tzjssx03b     (mf35lqg85lh2hl37 ),
      .cni2453cuofb     (f6zak916_6fg2ds06me ),
      .kt04okvuth    (trvcz0llenxn0vxzi),
      .kq9gup8pu2    (yql0f1_h8qzo314c),
      .g_o2wra9n9s        (in62nwnhf8t6xb5tt),
      .nykwng_3anppxi  (xvppde5hc39p611bfgybe5nse ),
      .shpynlimbt55rj4  (hgct1tjvcv_169taj843hl ),
      .jycwup76klyed6d2  (ev298h4twlq88a66tah_ ),
      .i7pubsxfsb4uys  (),
      .jc4yg1pkylr2gonwcd (kn86nder0b7le4a1_71fi),
      .nd3cgvec1pogf2 (gqb1ts5dtrjcr4lemz25tvya5n),
      .f7crsrzernrwgmepy (s_w7o2mb9s0hc170_6d06768n),
      .pw085ct76po3c  (ntcj3nmpwv67z623k_ach),
      .g5usf8ixwjaxjs1m   (),
      .pxhhgm9746n    (),
      .fgm5kq4y725x6yylw (dczlby2rwj8daf3344jiifcy),
      .awld9ngcypgfxa (bn4f_e4qqgexxu51ah0e8ef2),
      .v5m66onlnmxeejfhn (qb3a5cpzsa87m6bukrkbmo2vfu),
      .kfz3mojvfh2fsfd  (kr3sxd5ylio9sn5szxxpznd),


      .ng_pudjzgnamv0es (),
      .bdhv0j4zhtx9nxmz (dul93v3bagr1tk3h32    )

  );


  ihyzqc18e76a5lqw x4o1mt0tubfdgce0hxeg3k (
      .io8xbm86f       (kxblx1rz1zw1140nes         ),
      .qhyq467foflgyn5y(cmvxg4cmkkrry),
      .sa2f4h4xeakpfnunl(1'b0),
      .u2k4dyp52s_m     (suseox527co0by6rz  ),
      .djvj1e_     (pba6ait3opk6vu9lorcv3  ),
      .bktu0z1mk56     (mv01x26v2z8c6zft  ),

      .qbsr1jytrqtsbk4ttb8nz (qbsr1jytrqtsbk4ttb8nz),

      .sb8ax73d3ud   (r3q_xx2nluna_ybk80      ),
      .f9_w27gbcq__   (x6pwowdnpxkoegubqh      ),
      .iq9sj_i8z1k712   (ycu7j7ypp2g_tz59w7      ),
      .rig48lgqgq8oxt  (a8hdcsvsn4jfp6ggx0     ),
      .zaub9z0lm4s93y  (n40qc_n1g3r0iys56ldo2v     ),
      .j_69hsshtbv  (h4o95esg4yb2e820pv     ),

      .nnng_p6632p    (f93ucku8ja3u7_7jfc       ),
      .ld01d40_n3     (dbwm8k4yhgs_a5fh        ),
      .o8rwk067     (dj3vwzuwr1ayovji5        ),
      .r1on2k03r    (gr4bw39k1u2tog8       ),
      .gw7452ctd577    (nbvmheia5bzqvyguhpnt       ),
      .b1roq8tr9r     (ep9tb23giiqadx3q3po        ),
      .j_ku88w81rg     (khgn8edvptpzv6w8y        ),

      .t9xs6bqphiru  (),
      .ls1dudpc     (c6zn8c8zy_2ijgf ),
      .tzjssx03b     (dgapkwah8rq6xvlp8v ),
      .cni2453cuofb     (d4fnrrhamdmba5jc ),
      .kt04okvuth    (h1hqinnsgg8o7fj),
      .kq9gup8pu2    (ljz2177rfk7ofxrox),

      .g_o2wra9n9s        (z5ernaentmhkissw),
      .nykwng_3anppxi  (fl8fierzzigw8tj75cbg ),
      .shpynlimbt55rj4  (g2dg49ff5vl0cadcmalf ),
      .jycwup76klyed6d2  (pnw4fl90e287i2d45hqtkgf7w ),
      .i7pubsxfsb4uys  (),
      .jc4yg1pkylr2gonwcd (g9ujasz2f7mtbry7s8motw),
      .nd3cgvec1pogf2 (h533q7tm9n7oflpyzj7d7iz),
      .f7crsrzernrwgmepy (v9oxvr4ndit7gq_f97xdbpw),
      .pw085ct76po3c  (rie7ralfn6d1m5cmw5ofhaq0x),
      .g5usf8ixwjaxjs1m   (),
      .pxhhgm9746n    (),
      .fgm5kq4y725x6yylw (d5lmrsu7qp9zpkuxrkcwg2h5r),
      .awld9ngcypgfxa (jvt8l7ep5r4tybm2531os520t),
      .v5m66onlnmxeejfhn (mfptziquqbpd0ydd8vtdnpcioo),
      .kfz3mojvfh2fsfd  (),


      .ng_pudjzgnamv0es (),
      .bdhv0j4zhtx9nxmz (bn2eir5p36_6ayfded36    )

  );


  pgil4p_zywsz2lytb w5ddmyjyn3zv8uhn(

    .s7eq8f6z1uyi2in (s7eq8f6z1uyi2in),

    .hab9b2zcdgrlbutx5  (hab9b2zcdgrlbutx5),
    .uub2rxsi1qvmca  (uub2rxsi1qvmca),
    .p_xqcszydp2j5d821j  (p_xqcszydp2j5d821j),
    .hwpkcsh2atrq              (hwpkcsh2atrq  ),
    .v3e6l1k7eo9k3             (v3e6l1k7eo9k3 ),
    .hxrmt706n071lic0f7            (hxrmt706n071lic0f7),
    .horqgj1y_r_5aplro             (d4d7ru_yllps7en_tto),
    .iqaziwvuq5463k3            (iqaziwvuq5463k3),
    .hs5w0q7r19myj9eezz            (hs5w0q7r19myj9eezz),
    .q1zci4ybfd7ftj8qxl2           (n_lam8gs1mljgiq8zi),
    .vp5_qftup10p3v7_jw8           (gkonom22e0fpa2_v3w0ab),
    .v7rzl8qveorn2jg6659m69     (v7rzl8qveorn2jg6659m69),
    .v_k8ohy_e2e9vlp6az04        (v_k8ohy_e2e9vlp6az04),
    .p54semfzu2zyfb            (p54semfzu2zyfb),
    .m2_t547jr8crh6jgy4c           (m2_t547jr8crh6jgy4c),
    .y_vw514j6xmphhfhc         (y_vw514j6xmphhfhc),
    .gtvau5cygdmb10dr_makqf        (gtvau5cygdmb10dr_makqf),
    .ct8_j4rs_zvw4xjl_ncf      (ct8_j4rs_zvw4xjl_ncf),
    .ovuaqnjxywro47yxbn20wg3m     (ovuaqnjxywro47yxbn20wg3m),      

    .vmfcanu2o                    (rtszu4lyr6770b),
    .v5uyqoe                    (wsbbvfhbclor6q),
    .agjzm78wm                    (rphdzcfsv024),
    .v0u85q8u16_pwgz7h17cl4       (v0u85q8u16_pwgz7h17cl4),
    .yov0d70301nwd4bbqbyv       (yov0d70301nwd4bbqbyv),

    .pz6cvxcjpgv                (pxc1y6acd93),
    .haezj87elp_               (haezj87elp_),

    .z1p1oekb0pd                (uzl99yf1fjxt8l),
    .js_7wqgsstbnxcjr29           (te83d5pk716t4mlgz7b),
    .eajem3pnezl               (eajem3pnezl),

    .lln3b7iev7jpvogh964ro_9bc_3y    (lln3b7iev7jpvogh964ro_9bc_3y),
    .q97rqfy8n7ixfm2a5wev4nd5sylpcq3j   (q97rqfy8n7ixfm2a5wev4nd5sylpcq3j),
    .hujgg6hjnhtbspbkekuz5_u          (hujgg6hjnhtbspbkekuz5_u),
    .v3pnt81kfrgbaanm1mhh51w           (v3pnt81kfrgbaanm1mhh51w),
    .i08eq60d_snxeq8si_ezod          (i08eq60d_snxeq8si_ezod),
    .y8wz7aud_fd6dfiakjtx2i0g          (y8wz7aud_fd6dfiakjtx2i0g),
    .dgnjyd9xs8efyxm0tdlsvfq4eop         (dgnjyd9xs8efyxm0tdlsvfq4eop),
    .a3xib90kwk4_hm1                (a3xib90kwk4_hm1),
    .nfzexr8q9g893gi                 (nfzexr8q9g893gi),
    .opkkwp3eg8g3448t                (opkkwp3eg8g3448t),

    .bnjz04i86zhxx6                  (jpew88u43lex0gsdrxu  ),
    .qpotfvbjdo6qtsy1                 (lhom1sg0nscdxyh3 ),
    .ua8gydukonfboz                 (yt79c5htoexmnip5k7 ),
    .vkfewi0rkx                  (bclets06blmu6y9 ),
    .iq5y0wse0y2                  (a81rpsbwkeq0bzp  ),
    .ueimo2s8tf29_f              (dul93v3bagr1tk3h32  ),
    .jzcjplpewzvpowh                 (xfi53wrc_l8tkqw38hx9),
    .jvcw7os6duv6_6                  (dj3vwzuwr1ayovji5  ),
    .k0q5465tih57fj                 (gr4bw39k1u2tog8 ),
    .sfgacjvxnybsqrx_                 (nbvmheia5bzqvyguhpnt ),
    .z9lf1gw3iz9e                  (ep9tb23giiqadx3q3po ),
    .m_pst8fyu48q6i4                  (khgn8edvptpzv6w8y  ),
    .xl0lr2g890tskf74yu8              (bn2eir5p36_6ayfded36  ),
    .jvt4ma57k62vz                 (f93ucku8ja3u7_7jfc),

    .tbs7se44h1m47t              (tbs7se44h1m47t),


    .rhrr146mr7lt9h              (rhrr146mr7lt9h    ),
    .io1uhjqtpgin_              (io1uhjqtpgin_    ),
    .gohm8ye7tw32so            (yxu62lq_npmss6p3vt),
    .d0q_15ed0hmwqygja          (v2r90qa11qssvr5tq98dbi961),      
    .jrkjeqdo7hhdsjna            (jrkjeqdo7hhdsjna  ),  
    .cmvxg4cmkkrry            (cmvxg4cmkkrry  ),  
    .r9arh0s0wxc_0                (r9arh0s0wxc_0      ),
    .vgno0maw8a                (vgno0maw8a      ),
    .gj95joew8j70jj4               (gj95joew8j70jj4     ),
    .cs_6ujj3b74              (cs_6ujj3b74    ),
    .g1iutrfs                  (g1iutrfs        ),
    .dwz7mnj7ox5              (dwz7mnj7ox5    ),
    .nmy2nw74r7gg              (nmy2nw74r7gg    ),
    .v4gayo0h8l6na             (v4gayo0h8l6na   ),

    .gf33atgy                      (gf33atgy  ) ,
    .ru_wi                    (ru_wi )                 
  );

  wire [64-1:0] iwo1igeb;

  wire [64-1:0] nah57z24;
  wire ut4y9bv_r7eob;
  wire rnkqkip5uke1_olq;
  wire r0lgv_bfa6a28k;
  wire vm2hkxepo_3udjn6;


  wire [64-1:0] ozyc_k8_rcbqufei66;
  wire plc7tlf2gws62oywdzj4ca2__kt;
  wire b2veu37paw81_f_5egxmngj;
  wire tusc6mfb4hc575qagmdo7e;
  wire lyq6iwa9d6a3y3ssr0nm0s9nc13;
  wire tyrnjwe8oh5yh__ee4inl0tlsfwh;
  wire [4-1:0] mbomfmdp_sgf2onp_wvkxk;
  wire [4-1:0] qbaslok75k5x7i_qq6yt;
  wire [4-1:0] mehggpt2hh21ueizwhm3t8;
  wire [4-1:0] ls21nfiggg0eh3kdmsb9g;

  wire [4-1:0] a16a70eac34inq1vax6dtrbqz6n;
  wire [4-1:0] igryv8wus5rnmwriqfx422;

  assign grzq9ca3wtx8fvla2 = pxc1y6acd93 + 64'd2;
  assign ermp9v8eg4wjm = pxc1y6acd93 + 64'd4;
  assign cedxz601zu3p26 = pxc1y6acd93 + 64'd6;
  assign kregni2q7skqhzcey = pxc1y6acd93 + 64'd8;

  assign vncx4r8ansja = xfi53wrc_l8tkqw38hx9;
  assign w2jm73vsinhrawnk = f93ucku8ja3u7_7jfc;
  assign haezj87elp_ = xfi53wrc_l8tkqw38hx9 ?  ermp9v8eg4wjm : grzq9ca3wtx8fvla2;
  assign vcjsen3a1rld3379dy = ermp9v8eg4wjm;

  assign eajem3pnezl = ({64{((~vncx4r8ansja) & (~w2jm73vsinhrawnk))}} & ermp9v8eg4wjm)
                    |  ({64{(vncx4r8ansja ^ w2jm73vsinhrawnk)}} & cedxz601zu3p26)
                    |  ({64{(vncx4r8ansja & w2jm73vsinhrawnk)}} & kregni2q7skqhzcey)
                    ;
  assign iwo1igeb = eajem3pnezl;


  m1691tbt1_d8b0d7avy69zn w8o2_0kc0tp5nz4pw7jg5pe(
      .n38s98n2ak7rvsds      (1'b1),
      .vncx4r8ansja      (vncx4r8ansja),
      .w2jm73vsinhrawnk      (w2jm73vsinhrawnk),
      .k2mmowd1vvq       (iwo1igeb),
      .yddzpj5oad_dtepf (qbaslok75k5x7i_qq6yt),
      .gf33atgy              (gf33atgy),
      .ru_wi            (ru_wi)
  );

  m1691tbt1_d8b0d7avy69zn wa3n20i5wwp80j3f36_t2eo(
      .n38s98n2ak7rvsds      (1'b0),
      .vncx4r8ansja      (vncx4r8ansja),
      .w2jm73vsinhrawnk      (w2jm73vsinhrawnk),
      .k2mmowd1vvq       (h01d94xsxbxe_req),
      .yddzpj5oad_dtepf (mehggpt2hh21ueizwhm3t8),
      .gf33atgy              (gf33atgy),
      .ru_wi            (ru_wi)
  );

  m1691tbt1_d8b0d7avy69zn em6erktk0bz0fuo0bdkod73rz(
      .n38s98n2ak7rvsds      (1'b0),
      .vncx4r8ansja      (vncx4r8ansja),
      .w2jm73vsinhrawnk      (w2jm73vsinhrawnk),
      .k2mmowd1vvq       (jkzw_f9anx55),
      .yddzpj5oad_dtepf (ls21nfiggg0eh3kdmsb9g),
      .gf33atgy              (gf33atgy),
      .ru_wi            (ru_wi)
  );











  m1691tbt1_d8b0d7avy69zn q4d95decnyfevkvhi1nh4ufbc0(
      .n38s98n2ak7rvsds      (1'b0),
      .vncx4r8ansja      (vncx4r8ansja),
      .w2jm73vsinhrawnk      (w2jm73vsinhrawnk),
      .k2mmowd1vvq       ({{64-32{1'b0}},m9u9kwx2_i51v[31:0]}),
      .yddzpj5oad_dtepf (a16a70eac34inq1vax6dtrbqz6n),
      .gf33atgy              (gf33atgy),
      .ru_wi            (ru_wi)
  );

  m1691tbt1_d8b0d7avy69zn sjx4ex0v5qrfwbs7j3hh(
      .n38s98n2ak7rvsds      (1'b0),
      .vncx4r8ansja      (vncx4r8ansja),
      .w2jm73vsinhrawnk      (w2jm73vsinhrawnk),
      .k2mmowd1vvq       (wd9dvepxj),
      .yddzpj5oad_dtepf (igryv8wus5rnmwriqfx422),
      .gf33atgy              (gf33atgy),
      .ru_wi            (ru_wi)
  );

  assign{
      ozyc_k8_rcbqufei66,
      plc7tlf2gws62oywdzj4ca2__kt,
      b2veu37paw81_f_5egxmngj,
      tusc6mfb4hc575qagmdo7e,
      lyq6iwa9d6a3y3ssr0nm0s9nc13,
      tyrnjwe8oh5yh__ee4inl0tlsfwh,
      mbomfmdp_sgf2onp_wvkxk
  } = 
             (~(iu24hrsmr_23sjn
              | x34niohsf97hpd0ryaqi2f 
              | ovuaqnjxywro47yxbn20wg3m
              | uy9oz74i74jxm7_shj)) ? {
                                   iwo1igeb,
                                   wsbbvfhbclor6q,
                                   rphdzcfsv024,
                                   rtszu4lyr6770b,
                                   1'b0,
                                   1'b0,
                                   qbaslok75k5x7i_qq6yt
                              } :
               iu24hrsmr_23sjn ? {
                                 {h01d94xsxbxe_req[64-1:1],1'b0} ,
                                  tvqijouldcgiz2dxdco7,
                                  zkxlkidschdubxpkpm,
                                  xmcrni1qngfvh9pil9j,  
                                  1'b0,  
                                  1'b0,
                                  mehggpt2hh21ueizwhm3t8
                              } :
               x34niohsf97hpd0ryaqi2f ? {
                                {dhnoc09bxu7[64-1:1],1'b0} ,
                                 wsbbvfhbclor6q,
                                 rphdzcfsv024,
                                 rtszu4lyr6770b,  
                                 t3a424pkgkhyds9,
                                 zx8m32pgevhs66owv,
                                 kcdxflfd2aoaky4s22wdxu
                              } :
                uy9oz74i74jxm7_shj ?  {wd9dvepxj,
                                   1'b1,
                                   1'b0,
                                   1'b0,
                                   1'b0,
                                   1'b0,
                                  igryv8wus5rnmwriqfx422
                                  } :
                                {
                                  m9u9kwx2_i51v[64-1:1],1'b0,
                                  wsbbvfhbclor6q,
                                  rphdzcfsv024,
                                  rtszu4lyr6770b,

                                  t3a424pkgkhyds9,

                                  1'b1,
                                  a16a70eac34inq1vax6dtrbqz6n
                                } ;

                   
                   
                   
                   
                   
                   
                   

          
            
          
            
  wire t32i4f_wean0fa1u = ovuaqnjxywro47yxbn20wg3m & sje9n_dhyhybd3336mypqp & hab9b2zcdgrlbutx5;
  wire h84jhwgq85e_8p8xajgs = enwn0u48p2_ls5az80;
  wire o58peml2v6pl11f_qm = t32i4f_wean0fa1u | h84jhwgq85e_8p8xajgs;
  wire ux352jntr209cy617p = t32i4f_wean0fa1u | (~h84jhwgq85e_8p8xajgs);
  ux607_gnrl_dfflr #(1) haqyswon8lj0s7qp1 (o58peml2v6pl11f_qm, ux352jntr209cy617p, enwn0u48p2_ls5az80, gf33atgy, ru_wi);

  wire npohtdyi385u8igamq = ovuaqnjxywro47yxbn20wg3m & t2_c88voetamgqvcje26 & hab9b2zcdgrlbutx5;
  wire mqyl3ytxg_7hvtvmx = miax48k27o484e8a;
  wire pql0xjpw3o9tucj = npohtdyi385u8igamq | mqyl3ytxg_7hvtvmx;
  wire iw9yiiknfmncl9m = npohtdyi385u8igamq | (~mqyl3ytxg_7hvtvmx);
  ux607_gnrl_dfflr #(1) tg_m8g_aualx90xu5r86t (pql0xjpw3o9tucj, iw9yiiknfmncl9m, miax48k27o484e8a, gf33atgy, ru_wi);

  assign {nah57z24,
          ut4y9bv_r7eob,
          rnkqkip5uke1_olq,
          r0lgv_bfa6a28k,
          vm2hkxepo_3udjn6,
          yplsjnahawnbssor2hz,
          veno8k7ang7x3cxp_hme
          }
         = 
               n56voih_ovca1tcmk ? { {jkzw_f9anx55[64-1:1],1'b0},
                                  r_edve7v9jcr26q6zk,
                                  vrqfzuog2k4pos133,
                                  bmw2yi333716crywk,
                                  k2sr7sw1plcmnki5ajtscw,

                                  1'b0,
                                  ls21nfiggg0eh3kdmsb9g
                                  }:
                                      {ozyc_k8_rcbqufei66,
                                       plc7tlf2gws62oywdzj4ca2__kt,
                                       b2veu37paw81_f_5egxmngj,
                                       tusc6mfb4hc575qagmdo7e,
                                       lyq6iwa9d6a3y3ssr0nm0s9nc13,
                                       tyrnjwe8oh5yh__ee4inl0tlsfwh, 
                                       mbomfmdp_sgf2onp_wvkxk
                                      };












  wire y9hro6vutoqx = (~p0olq02_hyvx0) & (~c4ughu0qm5sfai);








  wire mzym3mjyce6op7zn0m = y9hro6vutoqx | uy9oz74i74jxm7_shj | s_emxwh6glh2gqasb;
  assign n38s98n2ak7rvsds = (~s_emxwh6glh2gqasb) & (~uy9oz74i74jxm7_shj) 
                              
						 & (~ovuaqnjxywro47yxbn20wg3m) 
                     ;
  assign azm2vbkop_ll3 = s_emxwh6glh2gqasb;




  wire j8a_43cdx81pgt6;
  wire oanfk7pkpni9hzi;
  assign mvkvkx9jdo5tp = ((~oanfk7pkpni9hzi) | j8a_43cdx81pgt6)


                        & sj1gaizva5__by20e
                       ;
  assign o87j_xf7v0e87   = (~oanfk7pkpni9hzi) | p_xqcszydp2j5d821j;




  assign jnq99nw1wv9zocbz = mzym3mjyce6op7zn0m & 
                             (mvkvkx9jdo5tp
                             & (
                                 (
                                    (iu24hrsmr_23sjn & hjri7cufo9ckntq) |
                                    (x34niohsf97hpd0ryaqi2f & wuqmf3xlyidrg5jh6756go) |
                                    (iu24hrsmr_23sjn & w1casjl7bz73brz) |
                                    (x34niohsf97hpd0ryaqi2f & n2shp8eftjcvx91gh47ib)
                                 ) ?
                                 1'b0 
                                 : 1'b1)
                             );


  wire wf91ifcqtxkbqyerz9q6h18etr1 = fd4mgmurz46g ? r_edve7v9jcr26q6zk : tvqijouldcgiz2dxdco7;
  wire g4a279amg33ex6_57dy7uk;
  wire ors9wur0wmegu7qddxfpx2c4tf = fd4mgmurz46g ? vrqfzuog2k4pos133 : zkxlkidschdubxpkpm;
  wire jzlx94zw2acljk3im4hk15y2;
  wire nkwymbx0pd31qyr0aogxh3t = fd4mgmurz46g ? bmw2yi333716crywk : xmcrni1qngfvh9pil9j;
  wire lsb7ew69pgpemlur555lf01cw;
  ux607_gnrl_dfflr #(1) seqfk5mdjv9nyi5mmfryapqa9b (z5zyhwuzrigmw, wf91ifcqtxkbqyerz9q6h18etr1, g4a279amg33ex6_57dy7uk, gf33atgy, ru_wi);  
  ux607_gnrl_dfflr #(1) x_rxyg2c8x4vy4mbgyz_dlgrxyb (z5zyhwuzrigmw, ors9wur0wmegu7qddxfpx2c4tf, jzlx94zw2acljk3im4hk15y2, gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1) h9h3b3oo_u6usipf_5tgmaxhxd (z5zyhwuzrigmw, nkwymbx0pd31qyr0aogxh3t, lsb7ew69pgpemlur555lf01cw, gf33atgy, ru_wi);
  
  assign f48_2zc1qro_3dodmk8 = (x34niohsf97hpd0ryaqi2f & n2shp8eftjcvx91gh47ib);
  assign vaiscz5bqo4k6ql0519 = g4a279amg33ex6_57dy7uk;  
  assign w93is2iaq5aikcpaqxg3 = jzlx94zw2acljk3im4hk15y2;
  assign uuuoq6te8sq6lj_e02iqoc = lsb7ew69pgpemlur555lf01cw;


  assign qmd94avv02av64cbwaj42 = (x34niohsf97hpd0ryaqi2f & wuqmf3xlyidrg5jh6756go);

  wire bai8bpslnudl4850_4gb40xefa_;
  wire c4wbt8uizx0iyxrktx4_3fms4i7e0   = fd4mgmurz46g ? lwdhmuzyvcvv14mjbl0h2a41z   : yghffofulqa77bd7aw07badta1a;
  wire [27-1:0] aclq6lmgg_xmnub38cwpw9;
  wire [27-1:0] klnha10og8cfk6uwba7tw = fd4mgmurz46g ? l4ztejmt2__wxqm2rw : zddoxp22m1o11x30gbe;
  wire ohi6wdfgenq5dzrw8j5w4uxp57t52;
  wire ub7a4h1wtxrthc6wvuftt3dx_upd = fd4mgmurz46g ? xy48dugh009wtmazqug3kpy2a5h_ : rrl7evvmayt1_vvp74iq9h6_cjf;
  wire [16-1:0] ug2d3cahrnebnrkj75ae;
  wire [16-1:0] c52o9bjl0hfs48b7ajntopi = fd4mgmurz46g ? s3ujdp2a8n69bm6engxok : hwfethpzkuauejcgtbl6o;

  ux607_gnrl_dfflr #(1)                bq9loxwdxbmpp_gluxo_r3sru_zr (z5zyhwuzrigmw, c4wbt8uizx0iyxrktx4_3fms4i7e0, bai8bpslnudl4850_4gb40xefa_, gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(27) mctgtto4yqosrslhpz0jhqsuw     (z5zyhwuzrigmw, klnha10og8cfk6uwba7tw,     aclq6lmgg_xmnub38cwpw9,     gf33atgy, ru_wi);

  ux607_gnrl_dfflr #(1)                rx773qavdmsh2ilho39kygpfikzjb6 (z5zyhwuzrigmw, ub7a4h1wtxrthc6wvuftt3dx_upd, ohi6wdfgenq5dzrw8j5w4uxp57t52, gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(16) l7o8pr50_6he4i9nml9lh0dijta     (z5zyhwuzrigmw, c52o9bjl0hfs48b7ajntopi,     ug2d3cahrnebnrkj75ae,    gf33atgy, ru_wi);

  assign m4ndmqnlr5eisc8m2k6fd   = bai8bpslnudl4850_4gb40xefa_;
  assign jcczlhzxqzl5dx51l       = aclq6lmgg_xmnub38cwpw9;
  assign nkdn__tk5pvp4nczp7xysy5 = ohi6wdfgenq5dzrw8j5w4uxp57t52;
  assign fhzpp1p52pmfd3syoo     = ug2d3cahrnebnrkj75ae;











  wire q_sekh_a09jcd5gbzj4ft = (s_emxwh6glh2gqasb) ? 1'b1 :

                          (y3p3payhiarg5b & sj1gaizva5__by20e);



  assign ht929tfpovwde = q_sekh_a09jcd5gbzj4ft;


  wire hmsefsbc0hea = uub2rxsi1qvmca | bn5omzf486_lr86nad3q01;

  ux607_gnrl_dfflr #(64) tlxfjudygg3x (hmsefsbc0hea, nah57z24, dhnoc09bxu7, gf33atgy, ru_wi);

  ux607_gnrl_dfflr #(1) de_ct2ia6twycduwbp (hmsefsbc0hea, ut4y9bv_r7eob, wsbbvfhbclor6q, gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1) qayp_tck742s1v (hmsefsbc0hea, rnkqkip5uke1_olq, rphdzcfsv024, gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1) jbl9gx_7q46706q (hmsefsbc0hea, r0lgv_bfa6a28k, rtszu4lyr6770b, gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1) uvldncxx64q6rogs55b (hmsefsbc0hea, vm2hkxepo_3udjn6, t3a424pkgkhyds9, gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1) ytmqb_dyurxmr695zv6 (hmsefsbc0hea, yplsjnahawnbssor2hz, zx8m32pgevhs66owv, gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(4) dw1tycu67_757wt5wmx0hu6m (hmsefsbc0hea, veno8k7ang7x3cxp_hme, kcdxflfd2aoaky4s22wdxu, gf33atgy, ru_wi);


  assign nupfecm_6ycs = dhnoc09bxu7;



  assign k2mmowd1vvq    = ozyc_k8_rcbqufei66;
  assign zc2e7csnzgj98szggj = plc7tlf2gws62oywdzj4ca2__kt |

                         tusc6mfb4hc575qagmdo7e;
  assign ih_5pl6hw4ippiu = b2veu37paw81_f_5egxmngj;
  assign y4vtwevsvl03ho6h0 = tusc6mfb4hc575qagmdo7e;
  assign hto4un7x8fe6gc1 = lyq6iwa9d6a3y3ssr0nm0s9nc13 & (~tyrnjwe8oh5yh__ee4inl0tlsfwh);
  assign agsse3cpfshpa0xh48nu0 = mbomfmdp_sgf2onp_wvkxk;



  wire o3gomcf2a7of6 = uub2rxsi1qvmca;

  assign j8a_43cdx81pgt6 = hab9b2zcdgrlbutx5;
  wire m4as0_0mwn8i8ghd7 = o3gomcf2a7of6 | j8a_43cdx81pgt6;

  wire hdc75b1l2il1s3 = o3gomcf2a7of6 | (~j8a_43cdx81pgt6);

  ux607_gnrl_dfflr #(1) z2m50x5taz3pbhcdro (m4as0_0mwn8i8ghd7, hdc75b1l2il1s3, oanfk7pkpni9hzi, gf33atgy, ru_wi);













endmodule




















module mu0arb3ch40modhq7(





  input  jnq99nw1wv9zocbz, 
  output sj1gaizva5__by20e, 




  input  [64-1:0] k2mmowd1vvq, 
  input  y4vtwevsvl03ho6h0, 
  input  hto4un7x8fe6gc1, 
  input  zc2e7csnzgj98szggj, 
  input  ih_5pl6hw4ippiu, 
  input [4-1:0] agsse3cpfshpa0xh48nu0,
  input  n38s98n2ak7rvsds, 

  input  vncx4r8ansja, 
  input  w2jm73vsinhrawnk, 


  output p_xqcszydp2j5d821j, 
  input  ht929tfpovwde, 
  output mkytk1e8mwi49l,   
  output xr81_h9hnhjwec3la,   
  output tbs7se44h1m47t,   
  output krxdptqk3busoihx2f,   
  output gnmzf7svwij0ih7c7fh3,   
  output we422ti7i_fjt8z36n53,   
  output tylsyqg3frnshrlcfkd596,   
  output rk6m6hfluv6syr3pz6z,   
  output eygoo8ifqdnay_dhiskf_,   
  output xfxeg_cwdrq6mzr3teo, 
  output diw3rbg3tca7kp6uu3l2n, 
  output [32*2-1:0] m9u9kwx2_i51v,

  input  azm2vbkop_ll3,






  output c52ldkop361ts52m0, 
  input  x88wat37r_vjsn57a, 
  output [64-1:0]   z3k8ps_o7osj4uosf_6i5, 
  output w8k_3fawz__hfg4mk0mw7g, 
  output i88maxesdvq1fkint66, 
  output rzon56p292pybf35mi_, 
  output jn_zyepkhmn_mdbqe1, 
  output ewekc8h7f7w9i3v,


  input  ult8a6a0b4agydwsws, 
  input  gkbxrtlrxlk7_fk4,   
  input  bwdpzndejgg3liwep6q_,   
  input  glkxypl9rxder9fztnegf6,   
  input  qe9n3_xo49nzqdf6gl2rz2j, 
  input  [64-1:0] d27a6w261um4big8wy8, 



  input  gf33atgy,
  input  ru_wi
  );





  wire jgn947pmmcm9a77iuey    ;
  wire lkrl_gk1f715er9ueo   ;
  wire dwmx63ax2_grri9q93qee;
  wire k8wf2zd3daqs6q    ;
  wire mpfnaagjnjijyse09ut;
  wire nifwkqncj1hl346947pv;
  wire g15fpvpqce7y5e_av;





  wire slg57kzkbyqfi7p8    = agsse3cpfshpa0xh48nu0[0];
  wire vp_6uj6bszug_1g34      = agsse3cpfshpa0xh48nu0[1];
  wire v566qwjezf2ts2jxc    = agsse3cpfshpa0xh48nu0[2];
  wire gb01708ufzq16d8brgoq = agsse3cpfshpa0xh48nu0[3];
  wire fqofqqtniw0hyim2uev = gb01708ufzq16d8brgoq;
  wire ka3r2ypzdt7fk6ci4 = vp_6uj6bszug_1g34 | slg57kzkbyqfi7p8;

  wire u36kqiqxmd6pckn8zv4;
  wire w75ygrz0e7wt0jtj;
  wire s025plocuxvzgndohb94ord;
  wire magm6h97w4rnyo73oyt0xr;

  wire uub2rxsi1qvmca = jnq99nw1wv9zocbz & sj1gaizva5__by20e;
  wire hab9b2zcdgrlbutx5 = p_xqcszydp2j5d821j & ht929tfpovwde;

  wire k0v4r1pl1uucldofmt ;
  wire yea5qwj5l_vv88mad ;
  wire eb079qwm5qlu_m3 ;

  ux607_gnrl_dfflr #(1) mp6ttw9ifh_50hty3o1k3926       (uub2rxsi1qvmca, fqofqqtniw0hyim2uev, u36kqiqxmd6pckn8zv4      , gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1) ma6h3hzdy18pnhplc7kjewjd       (uub2rxsi1qvmca, ka3r2ypzdt7fk6ci4, w75ygrz0e7wt0jtj      , gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1) ql0g6cra2xhdk2nua_ecffibyg_ (uub2rxsi1qvmca, v566qwjezf2ts2jxc  , s025plocuxvzgndohb94ord, gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1) c7qicm4ng4aa8a5g64jhtfcra90mw6 (uub2rxsi1qvmca, slg57kzkbyqfi7p8  , magm6h97w4rnyo73oyt0xr, gf33atgy, ru_wi);

  ux607_gnrl_dfflr #(1) gchby5brutg_77k9etuz7       (uub2rxsi1qvmca, zc2e7csnzgj98szggj  , k0v4r1pl1uucldofmt      , gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1) dzfmvwtx8t1rb9r3rq7473y       (uub2rxsi1qvmca, ih_5pl6hw4ippiu  , yea5qwj5l_vv88mad      , gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1) y_94xsbedyp1jls19e1ob       (uub2rxsi1qvmca, y4vtwevsvl03ho6h0  , eb079qwm5qlu_m3      , gf33atgy, ru_wi);











  assign c52ldkop361ts52m0 = 
                   (g15fpvpqce7y5e_av & (~ka3r2ypzdt7fk6ci4))
                 | ( 
                     (
                         (
                              mpfnaagjnjijyse09ut 
                              & jgn947pmmcm9a77iuey & nifwkqncj1hl346947pv
                         )
                       |  dwmx63ax2_grri9q93qee 
                     )
                   ) 
                     ;






  wire d3ztptp5gozov = 
                              mpfnaagjnjijyse09ut &
                                (
                                     jgn947pmmcm9a77iuey 
                                  |  dwmx63ax2_grri9q93qee
                                );

  wire s_izrbbfbb_qxwyp7nhlydfau = v566qwjezf2ts2jxc | d3ztptp5gozov;

  wire [64-1:0] ul0qbiyjsvnbbuxywpo;
  wire [64-1:0] tnm6toeraapgm49f = s_izrbbfbb_qxwyp7nhlydfau ? (ul0qbiyjsvnbbuxywpo + 64'd8) : k2mmowd1vvq[64-1:0]; 

  assign z3k8ps_o7osj4uosf_6i5   = {tnm6toeraapgm49f[64-1:3],3'b0};
  assign rzon56p292pybf35mi_  = d3ztptp5gozov ? k0v4r1pl1uucldofmt : zc2e7csnzgj98szggj;
  assign jn_zyepkhmn_mdbqe1  = d3ztptp5gozov ? yea5qwj5l_vv88mad : ih_5pl6hw4ippiu;
  assign w8k_3fawz__hfg4mk0mw7g  = d3ztptp5gozov ? eb079qwm5qlu_m3 : y4vtwevsvl03ho6h0; 
  assign i88maxesdvq1fkint66  = d3ztptp5gozov ? 1'b0  
                                          : hto4un7x8fe6gc1;
  assign ewekc8h7f7w9i3v    = d3ztptp5gozov ? 1'b1  
                                          : n38s98n2ak7rvsds  ; 

  wire l27lppmdcfek4zfdhaysa;


  ux607_gnrl_dfflr #(64)ervkanw10kpl5ty(l27lppmdcfek4zfdhaysa, z3k8ps_o7osj4uosf_6i5, ul0qbiyjsvnbbuxywpo, gf33atgy,ru_wi);








  wire t5uzgtynfhtgf4olrgh1 = 1'b1;



  assign l27lppmdcfek4zfdhaysa = c52ldkop361ts52m0 & x88wat37r_vjsn57a;
  assign nifwkqncj1hl346947pv = ult8a6a0b4agydwsws & t5uzgtynfhtgf4olrgh1;







  localparam fnk0axwxfk4kr8z  = 2;

  localparam i3mg661fq9njsp5b = 2'd0;

  localparam v_qy6klyvlpd9v  = 2'd1;

  localparam w7jie_pve8zo265khr8  = 2'd2;

  localparam elevjtxw8s86z  = 2'd3;

  wire [fnk0axwxfk4kr8z-1:0] brgdc0amsvlnwf_2j;
  wire [fnk0axwxfk4kr8z-1:0] rc887zv55nqt;
  wire gsoquod_6th_uva;
  wire [fnk0axwxfk4kr8z-1:0] u99tnldu986760c5   ;
  wire [fnk0axwxfk4kr8z-1:0] g9natvym5lqakd    ;
  wire [fnk0axwxfk4kr8z-1:0] qyw9w17wm01o0ibqri8;
  wire [fnk0axwxfk4kr8z-1:0] evn7vmlv0q87c    ;
  wire wfoen161d4r42bkqp34lj     ;
  wire oz66a4n0vakndgbkbj6ds      ;
  wire odvuoxdd_64egspdavi73jis74  ;
  wire z5xqhvuiqp_g510lj8      ;


  assign lkrl_gk1f715er9ueo    = (rc887zv55nqt == i3mg661fq9njsp5b   );
  assign jgn947pmmcm9a77iuey     = (rc887zv55nqt == v_qy6klyvlpd9v    );
  assign dwmx63ax2_grri9q93qee = (rc887zv55nqt == w7jie_pve8zo265khr8);
  assign k8wf2zd3daqs6q     = (rc887zv55nqt == elevjtxw8s86z    );



  assign wfoen161d4r42bkqp34lj = lkrl_gk1f715er9ueo & uub2rxsi1qvmca;
  assign u99tnldu986760c5      = v_qy6klyvlpd9v;






  wire sxzqcctniika3q3dr = azm2vbkop_ll3;
  assign mpfnaagjnjijyse09ut = u36kqiqxmd6pckn8zv4 & (~sxzqcctniika3q3dr);
  wire drclftccumhjlefb60z7k;
  assign oz66a4n0vakndgbkbj6ds  = jgn947pmmcm9a77iuey & ( 


                                  mpfnaagjnjijyse09ut ? nifwkqncj1hl346947pv : 

                                                      hab9b2zcdgrlbutx5
                             );
  assign g9natvym5lqakd     = 
                (


                  (mpfnaagjnjijyse09ut & (~x88wat37r_vjsn57a)) ?  w7jie_pve8zo265khr8


                  : (mpfnaagjnjijyse09ut & x88wat37r_vjsn57a) ?  elevjtxw8s86z 




                  :  uub2rxsi1qvmca  ?  v_qy6klyvlpd9v 
                                    : i3mg661fq9njsp5b 
                ) ;



  assign odvuoxdd_64egspdavi73jis74 = dwmx63ax2_grri9q93qee &  x88wat37r_vjsn57a;
  assign qyw9w17wm01o0ibqri8      = elevjtxw8s86z;



  assign z5xqhvuiqp_g510lj8     =  k8wf2zd3daqs6q &  hab9b2zcdgrlbutx5;
  assign evn7vmlv0q87c          = 
                (

                  uub2rxsi1qvmca  ?  v_qy6klyvlpd9v : 

                      i3mg661fq9njsp5b
                );


  assign gsoquod_6th_uva = 
            wfoen161d4r42bkqp34lj | oz66a4n0vakndgbkbj6ds | odvuoxdd_64egspdavi73jis74 | z5xqhvuiqp_g510lj8;


  assign brgdc0amsvlnwf_2j = 
              ({fnk0axwxfk4kr8z{wfoen161d4r42bkqp34lj   }} & u99tnldu986760c5   )
            | ({fnk0axwxfk4kr8z{oz66a4n0vakndgbkbj6ds    }} & g9natvym5lqakd    )
            | ({fnk0axwxfk4kr8z{odvuoxdd_64egspdavi73jis74}} & qyw9w17wm01o0ibqri8)
            | ({fnk0axwxfk4kr8z{z5xqhvuiqp_g510lj8    }} & evn7vmlv0q87c    )
              ;

  ux607_gnrl_dfflr #(fnk0axwxfk4kr8z) qo3f12wu71_4hg0af7 (gsoquod_6th_uva, brgdc0amsvlnwf_2j, rc887zv55nqt, gf33atgy, ru_wi);








  wire b5673_7cv0l2qvl7qdx;









  assign sj1gaizva5__by20e     = b5673_7cv0l2qvl7qdx;
  assign g15fpvpqce7y5e_av = jnq99nw1wv9zocbz    ;

  assign b5673_7cv0l2qvl7qdx = x88wat37r_vjsn57a;





  wire f88xgiwsvo_ph;

  wire yziovh6rad45ktlh9i  ;
  wire hrv7jqit17o3bnxxqlq2;
  wire ijb9eb_o_apvphqjdrm3ej;
  wire xubyqgpogd9nm951t2x1qc;

  wire  [64-1:0] byf_5_o878wbhi;
  wire                      yu_vk_mwzns85eu26bb;
  assign yu_vk_mwzns85eu26bb = uub2rxsi1qvmca;
  ux607_gnrl_dfflr #(64)xot4d_xp_78w0_k5halrs(yu_vk_mwzns85eu26bb, k2mmowd1vvq, byf_5_o878wbhi, gf33atgy,ru_wi);

  wire [64-1:0] vyftcg_87ws8dhccfcxcr5ey;
  wire [64-1:0] pc49yt8z6klka99r6lnymm1f39h2x_ = f88xgiwsvo_ph ? vyftcg_87ws8dhccfcxcr5ey  : d27a6w261um4big8wy8;






  wire [63:0] mjsj2y4wst3gbfo948bcb3wqro = pc49yt8z6klka99r6lnymm1f39h2x_;
  wire af7zapjnbp4vrx0xe3dt1ts775h            = f88xgiwsvo_ph ? yziovh6rad45ktlh9i    : gkbxrtlrxlk7_fk4;
  wire snewez3w02aqsm8clo5vz9_4xz         = f88xgiwsvo_ph ? hrv7jqit17o3bnxxqlq2 : bwdpzndejgg3liwep6q_;
  wire iennlmu2g8s3s9jvfq4njz6t5v         = f88xgiwsvo_ph ? ijb9eb_o_apvphqjdrm3ej : glkxypl9rxder9fztnegf6;
  wire rwlhcfou0abji4pgetbn6aokf5_n       = f88xgiwsvo_ph ? xubyqgpogd9nm951t2x1qc : qe9n3_xo49nzqdf6gl2rz2j;

  wire u3bt0ih6tml06mvzphzxl7auozttv;



  wire lk71uv07lku2w__ua1 = vp_6uj6bszug_1g34 & uub2rxsi1qvmca;
  wire udqc7gx9pbk42mauqn_nwenx = slg57kzkbyqfi7p8 & uub2rxsi1qvmca;
  wire od43drkwbgj7631vplfe = (
                           ((~f88xgiwsvo_ph) & ult8a6a0b4agydwsws & (~drclftccumhjlefb60z7k) & (~u3bt0ih6tml06mvzphzxl7auozttv)) 




                         | (lk71uv07lku2w__ua1)
                         | (udqc7gx9pbk42mauqn_nwenx)
                         );

  wire czm566ybbr56rgyb3dbc = f88xgiwsvo_ph & u3bt0ih6tml06mvzphzxl7auozttv;
  wire sgotfmhe202l8xm3 = od43drkwbgj7631vplfe | czm566ybbr56rgyb3dbc;
  wire w83qw1sck_d373r4su9b = od43drkwbgj7631vplfe | (~czm566ybbr56rgyb3dbc);
  ux607_gnrl_dfflr #(1)  xr2_0zr1q9r5d5be5pzot(sgotfmhe202l8xm3, w83qw1sck_d373r4su9b, f88xgiwsvo_ph, gf33atgy, ru_wi);



  wire ig9w7qm367yi1ecue1d6 = od43drkwbgj7631vplfe & (~f88xgiwsvo_ph);
  ux607_gnrl_dfflr  #(1)  d_rswdq30k8zpopk    (ig9w7qm367yi1ecue1d6, af7zapjnbp4vrx0xe3dt1ts775h   , yziovh6rad45ktlh9i   , gf33atgy, ru_wi);
  ux607_gnrl_dfflr  #(1)  x3673xvlsa97hprlau (ig9w7qm367yi1ecue1d6, snewez3w02aqsm8clo5vz9_4xz, hrv7jqit17o3bnxxqlq2, gf33atgy, ru_wi);
  ux607_gnrl_dfflr  #(1)  zjse41x00b3ebwft7 (ig9w7qm367yi1ecue1d6, iennlmu2g8s3s9jvfq4njz6t5v, ijb9eb_o_apvphqjdrm3ej, gf33atgy, ru_wi);
  ux607_gnrl_dfflr  #(1)  zlqtpw4u0jowm821mcttm (ig9w7qm367yi1ecue1d6, rwlhcfou0abji4pgetbn6aokf5_n, xubyqgpogd9nm951t2x1qc, gf33atgy, ru_wi);
  ux607_gnrl_dfflr  #(64) prhesrqsbmy7umgnx2aj603  (ig9w7qm367yi1ecue1d6, d27a6w261um4big8wy8 , vyftcg_87ws8dhccfcxcr5ey , gf33atgy, ru_wi);


  wire jf7qdoy6ozeijw19x9dlfxrt1xhd = f88xgiwsvo_ph | ult8a6a0b4agydwsws;








  wire q4zlija4136s_s9d; 
  wire [47:0] aafyam17vrqz; 
  wire [47:0] h3p0wpn_ah; 
  wire laa1t5iskus82m9g; 
  wire omyw5_07_btxhfwq; 
  wire xr82kspf8yl7mns9yxa4; 
  wire r9y8upslfevdvznk53cw; 
  wire sq1cgn76v6bze84un8cin5; 
  wire npf9pi7xlc7xl4t4b; 
  wire qs2xflsg9gu850zbd7_28qz_; 
  wire i6plop1aymkh0pxvx0bf; 

  wire ivjbjr1mdk46llnbceap = uub2rxsi1qvmca & v566qwjezf2ts2jxc;
  wire hppr8ic01_x1ug5dfsrc = nifwkqncj1hl346947pv & drclftccumhjlefb60z7k;

  assign q4zlija4136s_s9d = ivjbjr1mdk46llnbceap | hppr8ic01_x1ug5dfsrc;



  assign aafyam17vrqz = pc49yt8z6klka99r6lnymm1f39h2x_[64-1:64-48];
  assign laa1t5iskus82m9g = af7zapjnbp4vrx0xe3dt1ts775h;
  assign xr82kspf8yl7mns9yxa4 = snewez3w02aqsm8clo5vz9_4xz;
  assign sq1cgn76v6bze84un8cin5 = iennlmu2g8s3s9jvfq4njz6t5v;
  assign qs2xflsg9gu850zbd7_28qz_ = rwlhcfou0abji4pgetbn6aokf5_n;

  ux607_gnrl_dfflr #(48) rpr642x346c2b6r4ln     (q4zlija4136s_s9d, aafyam17vrqz,     h3p0wpn_ah,     gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1) xss7uzg8azp04e_lz9fpk_ (q4zlija4136s_s9d, laa1t5iskus82m9g, omyw5_07_btxhfwq, gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1) hz_w2jxw_fgnuj8t_8r1fl (q4zlija4136s_s9d, xr82kspf8yl7mns9yxa4, r9y8upslfevdvznk53cw, gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1) d8bi5mvibjnpij5qm_rrdo (q4zlija4136s_s9d, sq1cgn76v6bze84un8cin5, npf9pi7xlc7xl4t4b, gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1) jnei71cnk4eklcqrxcvtpw6vb2u (q4zlija4136s_s9d, qs2xflsg9gu850zbd7_28qz_, i6plop1aymkh0pxvx0bf, gf33atgy, ru_wi);









  wire sh62jig2oeu1ga1pbr8f97lop3ye1c = jgn947pmmcm9a77iuey & w75ygrz0e7wt0jtj;





  assign drclftccumhjlefb60z7k = mpfnaagjnjijyse09ut & jgn947pmmcm9a77iuey;

  wire w0vcmzwl1n3hit2kqasddu4;
  wire igrebzi1pot9gibne_iy577x;

  assign p_xqcszydp2j5d821j = sh62jig2oeu1ga1pbr8f97lop3ye1c | igrebzi1pot9gibne_iy577x;
  assign w0vcmzwl1n3hit2kqasddu4 = ht929tfpovwde;
  assign igrebzi1pot9gibne_iy577x     = drclftccumhjlefb60z7k ? 1'b0 : jf7qdoy6ozeijw19x9dlfxrt1xhd;
  assign u3bt0ih6tml06mvzphzxl7auozttv = drclftccumhjlefb60z7k ? 1'b1 : w0vcmzwl1n3hit2kqasddu4;
















  wire bcv12lwzxo4ealg7fe9wog = (   jgn947pmmcm9a77iuey
                                  & s025plocuxvzgndohb94ord
                                )
                              | magm6h97w4rnyo73oyt0xr
                              | k8wf2zd3daqs6q;



  wire du89d6il56ogw5n1sdzzf = byf_5_o878wbhi[2:1] == 2'b00;
  wire wv9ucw6pn_cffizpe85bg = byf_5_o878wbhi[2:1] == 2'b01;
  wire w0xhd1q8_mibjwtvbnn = byf_5_o878wbhi[2:1] == 2'b10;
  wire nosxixgnhdcjj0ii2y = byf_5_o878wbhi[2:1] == 2'b11;
  wire [63:0] dni5qarmjaojzk3q8ytuhp9edxwt08 =  
                                                ({64{wv9ucw6pn_cffizpe85bg}} & {mjsj2y4wst3gbfo948bcb3wqro[15:0], h3p0wpn_ah[47:0]}) 
                                            |   ({64{w0xhd1q8_mibjwtvbnn}} & {mjsj2y4wst3gbfo948bcb3wqro[31:0], h3p0wpn_ah[47:16]}) 
                                            |   ({64{nosxixgnhdcjj0ii2y}} & {mjsj2y4wst3gbfo948bcb3wqro[47:0], h3p0wpn_ah[47:32]}) 
                                            ;

  assign m9u9kwx2_i51v  =  bcv12lwzxo4ealg7fe9wog ? dni5qarmjaojzk3q8ytuhp9edxwt08 : mjsj2y4wst3gbfo948bcb3wqro;


  assign tbs7se44h1m47t    =  bcv12lwzxo4ealg7fe9wog ? (|{af7zapjnbp4vrx0xe3dt1ts775h, omyw5_07_btxhfwq}) : af7zapjnbp4vrx0xe3dt1ts775h; 

  wire  o_ry9q1q7jm1wwv    =  bcv12lwzxo4ealg7fe9wog & (af7zapjnbp4vrx0xe3dt1ts775h & (~omyw5_07_btxhfwq));
  wire klrvngiy5eeicqbwnh_du1m = vncx4r8ansja & nosxixgnhdcjj0ii2y & o_ry9q1q7jm1wwv;
  wire e_w8wpj43wzby687fwgzx22 = ( (wv9ucw6pn_cffizpe85bg & vncx4r8ansja)
                            | (w0xhd1q8_mibjwtvbnn & (~vncx4r8ansja))) & w2jm73vsinhrawnk & o_ry9q1q7jm1wwv;
  assign krxdptqk3busoihx2f = ~klrvngiy5eeicqbwnh_du1m; 
  assign gnmzf7svwij0ih7c7fh3 = ~e_w8wpj43wzby687fwgzx22; 

  wire fgvaa79vt1ptlny6t5ljr_n_umyk1z = (nosxixgnhdcjj0ii2y & vncx4r8ansja) ? (snewez3w02aqsm8clo5vz9_4xz | r9y8upslfevdvznk53cw)
                                                              :  r9y8upslfevdvznk53cw;
  wire a8p0jz9dycmstf_fux7t5lnt06f = (
                               (
                                   du89d6il56ogw5n1sdzzf
                                | (wv9ucw6pn_cffizpe85bg & (~(vncx4r8ansja & w2jm73vsinhrawnk)))                                                                
                                | (w0xhd1q8_mibjwtvbnn & (~vncx4r8ansja) & (~w2jm73vsinhrawnk))
                                ) &     r9y8upslfevdvznk53cw)
                           | (
                               (
                                (wv9ucw6pn_cffizpe85bg & vncx4r8ansja & w2jm73vsinhrawnk) 
                              | (w0xhd1q8_mibjwtvbnn & (~vncx4r8ansja) & w2jm73vsinhrawnk)
                               ) & (snewez3w02aqsm8clo5vz9_4xz | r9y8upslfevdvznk53cw)
                             )
                           | (
                               (
                                (w0xhd1q8_mibjwtvbnn & vncx4r8ansja)
                              |  nosxixgnhdcjj0ii2y
                               ) & snewez3w02aqsm8clo5vz9_4xz 
                             )
                           ;

  wire fftdeu_8zbzxqpk6knsxnh2g_qz = (nosxixgnhdcjj0ii2y & vncx4r8ansja) ? (iennlmu2g8s3s9jvfq4njz6t5v | npf9pi7xlc7xl4t4b)
                                                              :  npf9pi7xlc7xl4t4b;
  wire m8t2ise7ogia9g4oodl405jx2b = (
                               (
                                   du89d6il56ogw5n1sdzzf
                                | (wv9ucw6pn_cffizpe85bg & (~(vncx4r8ansja & w2jm73vsinhrawnk)))                                                                
                                | (w0xhd1q8_mibjwtvbnn & (~vncx4r8ansja) & (~w2jm73vsinhrawnk))
                                ) &     npf9pi7xlc7xl4t4b)
                           | (
                               (
                                (wv9ucw6pn_cffizpe85bg & vncx4r8ansja & w2jm73vsinhrawnk) 
                              | (w0xhd1q8_mibjwtvbnn & (~vncx4r8ansja) & w2jm73vsinhrawnk)
                               ) & (iennlmu2g8s3s9jvfq4njz6t5v | npf9pi7xlc7xl4t4b)
                             )
                           | (
                               (
                                (w0xhd1q8_mibjwtvbnn & vncx4r8ansja)
                              |  nosxixgnhdcjj0ii2y
                               ) & iennlmu2g8s3s9jvfq4njz6t5v 
                             )
                           ;


  wire mv9qf6cuorsf29ydy5dt3io54te_z_nm = (nosxixgnhdcjj0ii2y & vncx4r8ansja) ? (rwlhcfou0abji4pgetbn6aokf5_n | i6plop1aymkh0pxvx0bf)
                                                              :  i6plop1aymkh0pxvx0bf;
  wire e34d0olqorsoa63c2x8o9zjlwj0gl = (
                               (
                                   du89d6il56ogw5n1sdzzf
                                | (wv9ucw6pn_cffizpe85bg & (~(vncx4r8ansja & w2jm73vsinhrawnk)))                                                                
                                | (w0xhd1q8_mibjwtvbnn & (~vncx4r8ansja) & (~w2jm73vsinhrawnk))
                                ) &     i6plop1aymkh0pxvx0bf)
                           | (
                               (
                                (wv9ucw6pn_cffizpe85bg & vncx4r8ansja & w2jm73vsinhrawnk) 
                              | (w0xhd1q8_mibjwtvbnn & (~vncx4r8ansja) & w2jm73vsinhrawnk)
                               ) & (rwlhcfou0abji4pgetbn6aokf5_n | i6plop1aymkh0pxvx0bf)
                             )
                           | (
                               (
                                (w0xhd1q8_mibjwtvbnn & vncx4r8ansja)
                              |  nosxixgnhdcjj0ii2y
                               ) & rwlhcfou0abji4pgetbn6aokf5_n 
                             )
                           ;

  assign we422ti7i_fjt8z36n53 =  bcv12lwzxo4ealg7fe9wog ? fgvaa79vt1ptlny6t5ljr_n_umyk1z : snewez3w02aqsm8clo5vz9_4xz;                            
  assign tylsyqg3frnshrlcfkd596 =  bcv12lwzxo4ealg7fe9wog ? a8p0jz9dycmstf_fux7t5lnt06f : snewez3w02aqsm8clo5vz9_4xz;                            
  assign rk6m6hfluv6syr3pz6z =  bcv12lwzxo4ealg7fe9wog ? fftdeu_8zbzxqpk6knsxnh2g_qz : iennlmu2g8s3s9jvfq4njz6t5v;                            
  assign eygoo8ifqdnay_dhiskf_ =  bcv12lwzxo4ealg7fe9wog ? m8t2ise7ogia9g4oodl405jx2b : iennlmu2g8s3s9jvfq4njz6t5v;                            
  assign xfxeg_cwdrq6mzr3teo =  bcv12lwzxo4ealg7fe9wog ? mv9qf6cuorsf29ydy5dt3io54te_z_nm : rwlhcfou0abji4pgetbn6aokf5_n;                            
  assign diw3rbg3tca7kp6uu3l2n =  bcv12lwzxo4ealg7fe9wog ? e34d0olqorsoa63c2x8o9zjlwj0gl : rwlhcfou0abji4pgetbn6aokf5_n;                            

  wire ijxng7c1h5vv59od5ph7yq4y4 = (nosxixgnhdcjj0ii2y & vncx4r8ansja) ? (af7zapjnbp4vrx0xe3dt1ts775h | omyw5_07_btxhfwq)
                                                              :  omyw5_07_btxhfwq;
  wire y9pn1aaitlj0xrjujkhbhx87 = (
                               (
                                   du89d6il56ogw5n1sdzzf
                                | (wv9ucw6pn_cffizpe85bg & (~(vncx4r8ansja & w2jm73vsinhrawnk)))                                                                
                                | (w0xhd1q8_mibjwtvbnn & (~vncx4r8ansja) & (~w2jm73vsinhrawnk))
                                ) &     omyw5_07_btxhfwq)
                           | (
                               (
                                (wv9ucw6pn_cffizpe85bg & vncx4r8ansja & w2jm73vsinhrawnk) 
                              | (w0xhd1q8_mibjwtvbnn & (~vncx4r8ansja) & w2jm73vsinhrawnk)
                               ) & (af7zapjnbp4vrx0xe3dt1ts775h | omyw5_07_btxhfwq)
                             )
                           | (
                               (
                                (w0xhd1q8_mibjwtvbnn & vncx4r8ansja)
                              |  nosxixgnhdcjj0ii2y
                               ) & af7zapjnbp4vrx0xe3dt1ts775h 
                             )
                           ;
  assign mkytk1e8mwi49l = bcv12lwzxo4ealg7fe9wog ? ijxng7c1h5vv59od5ph7yq4y4 : af7zapjnbp4vrx0xe3dt1ts775h;                            
  assign xr81_h9hnhjwec3la = bcv12lwzxo4ealg7fe9wog ? y9pn1aaitlj0xrjujkhbhx87 : af7zapjnbp4vrx0xe3dt1ts775h;                            









endmodule





















module ihyzqc18e76a5lqw(



  input  [32-1:0] io8xbm86f,

  input  qhyq467foflgyn5y,
  input  sa2f4h4xeakpfnunl,
  input  u2k4dyp52s_m,
  input  djvj1e_,
  input  bktu0z1mk56,




  input  qbsr1jytrqtsbk4ttb8nz,

  output g_o2wra9n9s,
  output nykwng_3anppxi,
  output shpynlimbt55rj4,
  output jycwup76klyed6d2,
  output i7pubsxfsb4uys,
  output [5-1:0] jc4yg1pkylr2gonwcd,
  output [5-1:0] nd3cgvec1pogf2,
  output [5-1:0] f7crsrzernrwgmepy,
  output [5-1:0] pw085ct76po3c,
  output [48-1:0] g5usf8ixwjaxjs1m,
  output [64-1:0] pxhhgm9746n,
  output fgm5kq4y725x6yylw,
  output awld9ngcypgfxa,
  output v5m66onlnmxeejfhn,
  output kfz3mojvfh2fsfd,


  output sb8ax73d3ud,
  output f9_w27gbcq__,

  output iq9sj_i8z1k712,
  output [5-1:0] rig48lgqgq8oxt,
  output [5-1:0] zaub9z0lm4s93y,
  output [5-1:0] j_69hsshtbv,

  output t9xs6bqphiru,
  output ls1dudpc   ,
  output tzjssx03b   ,
  output cni2453cuofb   ,
  output kt04okvuth  ,
  output kq9gup8pu2  ,

  output nnng_p6632p,
  output ld01d40_n3,
  output o8rwk067,
  output r1on2k03r,
  output gw7452ctd577,
  output b1roq8tr9r,
  output j_ku88w81rg,
  output [5-1:0] ng_pudjzgnamv0es,
  output [64-1:0] bdhv0j4zhtx9nxmz 

  );

  jgz9v2pi3n5adi7j41 b2163wfvtrtbqnnjbc0fx(

  .k0xug5g(io8xbm86f),
  .qhyq467foflgyn5y(qhyq467foflgyn5y),
  .sa2f4h4xeakpfnunl(sa2f4h4xeakpfnunl),

  .qbsr1jytrqtsbk4ttb8nz(qbsr1jytrqtsbk4ttb8nz),

  .b0ry73kp6sc2 (1'b0),
  .hr64e6c3gy  (1'b0),
  .cz1hh6af7xp2 (1'b0),

  .s1woka0byzgo    (1'b0),
  .al4xeg8mukgfg      (1'b0),
  .piwiqvrjoq     (1'b0),
  .wi_dfzp70x09hm1m  (1'b0),
  .jdyqycv3wdp2sgy(1'b0),


  .fpwql5ik7_sp0(),
  .dwci8hbxok739(),

  .mg0onistbzu9ys(),
  .g3btysb7vvv(),
  .yjgkn7vcv(),
  .sb8ax73d3ud(sb8ax73d3ud),
  .f9_w27gbcq__(f9_w27gbcq__),
  .iq9sj_i8z1k712(iq9sj_i8z1k712),

  .b6cv9yeaga7hf(),
  .rig48lgqgq8oxt(rig48lgqgq8oxt),
  .zaub9z0lm4s93y(zaub9z0lm4s93y),
  .j_69hsshtbv(j_69hsshtbv),
  .kd6v2vk601xpnm(),
  .t05leas4w4r(),

  .u2k4dyp52s_m(u2k4dyp52s_m),
  .djvj1e_(djvj1e_),
  .bktu0z1mk56(bktu0z1mk56),
  .fqizcmmfg (),
  .tbuacpjktio (),
  .ciftsjs2bvaxns (),
  .k_y4yq3crp_zqtg(),

  .qzdlalytscynhz1 (),

  .vfye1vj155_k  (),
  .vujduks2o30  (),
  .y4zqru1tedm  (),
  .q1coyps2cz7xe  (),
  .oli3_udj80h6urj  (),
  .rphjsg75001l2 (),
  .ch8qv98q9xu469etyz8oj(),
  .zj0wqwminaxn(),
  .jw1vgacy_r0vr(),


  .hgvdw0qnels8(),


  .rnx27onf2lbe     (1'b0),
  .g_o2wra9n9s        (g_o2wra9n9s),
  .nykwng_3anppxi  (nykwng_3anppxi ),
  .shpynlimbt55rj4  (shpynlimbt55rj4 ),
  .jycwup76klyed6d2  (jycwup76klyed6d2 ),
  .i7pubsxfsb4uys  (i7pubsxfsb4uys ),
  .jc4yg1pkylr2gonwcd (jc4yg1pkylr2gonwcd),
  .nd3cgvec1pogf2 (nd3cgvec1pogf2),
  .f7crsrzernrwgmepy (f7crsrzernrwgmepy),
  .pw085ct76po3c  (pw085ct76po3c),
  .g5usf8ixwjaxjs1m   (g5usf8ixwjaxjs1m ),
  .pxhhgm9746n    (pxhhgm9746n  ),
  .fgm5kq4y725x6yylw (fgm5kq4y725x6yylw),
  .awld9ngcypgfxa (awld9ngcypgfxa),
  .v5m66onlnmxeejfhn (v5m66onlnmxeejfhn),
  .kfz3mojvfh2fsfd  (kfz3mojvfh2fsfd),
  .m05tjqf24b1fabuu0e(),

   .d40y0va2l7xzj    (               ),
   .hhj5975j18r0n  (               ),

  .t9xs6bqphiru(t9xs6bqphiru),
  .ls1dudpc   (ls1dudpc   ),
  .tzjssx03b   (tzjssx03b   ),
  .cni2453cuofb   (cni2453cuofb   ),
  .kt04okvuth  (kt04okvuth  ),
  .kq9gup8pu2  (kq9gup8pu2  ),


  .eaxqugrf_ryu5rxxw41(),
  .tkm5u9dl8zav4(),
  .z8t7w6zr5woh649(),
  .mg4yq4mui7ruja(),
  .sibtd2rf5j(),


  .nnng_p6632p(nnng_p6632p),
  .ld01d40_n3 (ld01d40_n3 ),
  .o8rwk067 (o8rwk067 ),
  .r1on2k03r(r1on2k03r),
  .gw7452ctd577(gw7452ctd577),
  .b1roq8tr9r (b1roq8tr9r),
  .j_ku88w81rg (j_ku88w81rg ),
  .zk9uk90j08ogqpn(),
  .ng_pudjzgnamv0es(ng_pudjzgnamv0es),
  .bdhv0j4zhtx9nxmz    (bdhv0j4zhtx9nxmz    )  
  );


endmodule




















module ftui9s73ym2ff #(
  parameter nm_fj = 32,
  parameter s3xvyho = 32,
  parameter onr7l = 32
)(
  output ny26eoy00tenwa,

  input  c52ldkop361ts52m0,
  output x88wat37r_vjsn57a,
  input  [nm_fj-1:0] z3k8ps_o7osj4uosf_6i5,
  input  w8k_3fawz__hfg4mk0mw7g,
  input  i88maxesdvq1fkint66,
  input  rzon56p292pybf35mi_,
  input  jn_zyepkhmn_mdbqe1,
  input  ewekc8h7f7w9i3v,

  output ult8a6a0b4agydwsws,
  output gkbxrtlrxlk7_fk4,   
  output [s3xvyho-1:0] fw895kfvwds4i_6uy,
  output [onr7l-1:0] d27a6w261um4big8wy8, 

  output q9uknlmu4747layzj7,
  input  vlhrtmmnzbn11e0gw,
  output [nm_fj-1:0] ui2ziibknh_1uaiixo0m1,
  output kpptfyyykyfkwr_w7zz,
  output oz7xvqjtmxw3yf4j3,
  output mqdln_zof0pm8dvg2cb_e,
  output ll0zpg0jpkuqhp9f55h,

  input  hxhn_tu5eqc44_0avu,
  input  e9kdetktxle114zq31ok,   
  input  [s3xvyho-1:0] lqxbdzkfs0nroxbl0r1f,   
  input  [onr7l-1:0] pnsc2d5vs30dex7_jy61, 

  output bf61lpqg8z,

  input  gf33atgy,
  input  ru_wi
  );



  wire v9ov1b3vn5k4ctkb;
  wire ub9pjiu4juf6nuqoq2w6;
  wire [nm_fj-1:0] aw0a19a967dn7n0x25w;
  wire cwkq4r6_upg_2884r;
  wire air1drtzqvyz1ydvdej;
  wire ty6a2k41y0e9ir8_yzg;
  wire s4_gwe0uskrbhp37ksb;
  wire d4yudirhr1quwh;

  localparam f16zrowg1s1f5 = (nm_fj + 5);

  wire [f16zrowg1s1f5-1:0]djfdd4cy1d_i5vg;
  wire [f16zrowg1s1f5-1:0]lehbgtu_h616v3v3nzq;

  assign lehbgtu_h616v3v3nzq = {
                             z3k8ps_o7osj4uosf_6i5 
                            ,w8k_3fawz__hfg4mk0mw7g 
                            ,i88maxesdvq1fkint66 
                            ,rzon56p292pybf35mi_ 
                            ,jn_zyepkhmn_mdbqe1 
                            ,ewekc8h7f7w9i3v 
                          };

  assign {
                             aw0a19a967dn7n0x25w 
                            ,cwkq4r6_upg_2884r 
                            ,air1drtzqvyz1ydvdej 
                            ,ty6a2k41y0e9ir8_yzg 
                            ,s4_gwe0uskrbhp37ksb 
                            ,d4yudirhr1quwh 
                          } = djfdd4cy1d_i5vg;

  
  
  




  ux607_gnrl_bypbuf # (
    .DP(1),
    .DW(f16zrowg1s1f5) 
  ) eewsgqzf8478ca8abhd(
      .i_vld   (c52ldkop361ts52m0),
      .i_rdy   (x88wat37r_vjsn57a),

      .o_vld   (v9ov1b3vn5k4ctkb),
      .o_rdy   (ub9pjiu4juf6nuqoq2w6),

      .i_dat   (lehbgtu_h616v3v3nzq),
      .o_dat   (djfdd4cy1d_i5vg),
  
      .clk     (gf33atgy  ),
      .rst_n   (ru_wi)
  );


  wire fppz16b2vnxcgbxo5flw_ni5a; 
  wire otr0zqv99dzgqhnaqt3wmawo; 
  wire bo4tz80rb2i3jzf7tz05t39;
  wire v3ov4l_sfrqtd5gzo = q9uknlmu4747layzj7 & vlhrtmmnzbn11e0gw;
  wire t1y5bixqb70xoxpulhmy = hxhn_tu5eqc44_0avu;
  wire pl83axr4i6pmpf58jv1pqg_x = fppz16b2vnxcgbxo5flw_ni5a;

  wire nwjse95ua1izg3w0h4f;
     
  wire dr_nl9fj18dp_b8jcn = v9ov1b3vn5k4ctkb & ub9pjiu4juf6nuqoq2w6;
  
  wire atj5hrqo8hgpcem = ult8a6a0b4agydwsws;
  wire bfrjyl3w5yfnw5fneojkay = dr_nl9fj18dp_b8jcn;
     
  wire cq3l45rsxc6gmvfl5vcje = atj5hrqo8hgpcem;
  wire j9kahccisrvimcfsmyg0 = bfrjyl3w5yfnw5fneojkay | cq3l45rsxc6gmvfl5vcje;
     
  wire lzuix0hy34qwode9gpsgrna = bfrjyl3w5yfnw5fneojkay | (~cq3l45rsxc6gmvfl5vcje);

  ux607_gnrl_dfflr #(1) yep4r8guk9hnj0_spacsbfj35 (j9kahccisrvimcfsmyg0, lzuix0hy34qwode9gpsgrna, nwjse95ua1izg3w0h4f, gf33atgy, ru_wi);

  wire z5w_j675ghcegxz91   = (~nwjse95ua1izg3w0h4f);


  wire chbqdc7gjz5vh433w5m = z5w_j675ghcegxz91 | (cq3l45rsxc6gmvfl5vcje);



  wire kcv48ukn4yb7uxlfz_l76v6;
  wire ab3stth5phu3zhxwjv1re;

  wire rucga3znd8eyg82;
  wire qly6mxgi154d4;
  wire st7pytysu10a;
  wire w2w3fpyeldr0;

  
    
    
    
  wire j1rvopf2x3yuqsb = (~d4yudirhr1quwh) & chbqdc7gjz5vh433w5m;

  wire fpfmc99sca  = 1'b1;

  assign ub9pjiu4juf6nuqoq2w6 = 
       (fpfmc99sca ? qly6mxgi154d4 : 1'b1)
     & (j1rvopf2x3yuqsb ? ab3stth5phu3zhxwjv1re : 1'b1);

  assign rucga3znd8eyg82        = fpfmc99sca  & v9ov1b3vn5k4ctkb & (j1rvopf2x3yuqsb ? ab3stth5phu3zhxwjv1re : 1'b1);
  assign kcv48ukn4yb7uxlfz_l76v6 = j1rvopf2x3yuqsb & v9ov1b3vn5k4ctkb & (fpfmc99sca  ? qly6mxgi154d4        : 1'b1);


  ux607_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(1)
  ) vsmkuuhmv71me (
    .i_vld(rucga3znd8eyg82), 
    .i_rdy(qly6mxgi154d4), 
    .i_dat(1'b0),
    .o_vld(st7pytysu10a), 
    .o_rdy(w2w3fpyeldr0), 
    .o_dat(),
  
    .clk  (gf33atgy  ),
    .rst_n(ru_wi)  
   );

  wire x_ua3ig1haanymrcfrqq = kcv48ukn4yb7uxlfz_l76v6 & ab3stth5phu3zhxwjv1re;

  wire k4ycbfysqrx0usx5lyog437;
  wire lzsa6zlhsqoszi5p0r8q;

    
        
  assign ult8a6a0b4agydwsws = st7pytysu10a & k4ycbfysqrx0usx5lyog437;
  
    
  assign w2w3fpyeldr0 = k4ycbfysqrx0usx5lyog437;

    
  assign lzsa6zlhsqoszi5p0r8q = st7pytysu10a;

  wire bhlov58es2dpzr2ee = j1rvopf2x3yuqsb & v9ov1b3vn5k4ctkb;

  
  bh912j8o17nne6z_zsk9c # (
    .tcebpmbl7g (0),
    .mhdlk  (5),
    .onr7l  (onr7l+1+s3xvyho)
  ) nveohbhbnsoukk71dy7823fn (
        
    .veibgbyke(bhlov58es2dpzr2ee),
    .bw6ftrau0  (fppz16b2vnxcgbxo5flw_ni5a),
    .eef2g8  (otr0zqv99dzgqhnaqt3wmawo),
    .p3mxtqc2ivbcmm0(bo4tz80rb2i3jzf7tz05t39),
    .qbjvs30wtb  ({pnsc2d5vs30dex7_jy61, e9kdetktxle114zq31ok, lqxbdzkfs0nroxbl0r1f}),
    .wqljp  (k4ycbfysqrx0usx5lyog437),
    .h9378  (lzsa6zlhsqoszi5p0r8q),  
    .dqgck5s  ({d27a6w261um4big8wy8, gkbxrtlrxlk7_fk4, fw895kfvwds4i_6uy}),  
    .gf33atgy    (gf33atgy),
    .ru_wi  (ru_wi)
  );

  wire l2qiuit0jdaq2pbqot;
  wire h3tgasjwjf9pjoc3uvwxw = v3ov4l_sfrqtd5gzo & j1rvopf2x3yuqsb;
  wire bbi2mz3lt21kyervd = h3tgasjwjf9pjoc3uvwxw;
  wire z_9eqe_kqw352t = t1y5bixqb70xoxpulhmy & l2qiuit0jdaq2pbqot;
  wire l22dfv0bi6ta7i8 = bbi2mz3lt21kyervd | z_9eqe_kqw352t;
  wire lsn_s8i0xwjf_7o0k = bbi2mz3lt21kyervd | (~z_9eqe_kqw352t);
  wire k7w9hbbfq2amb;
  ux607_gnrl_dfflr #(1) u_43i10vfbwu1447 (l22dfv0bi6ta7i8, lsn_s8i0xwjf_7o0k, k7w9hbbfq2amb, gf33atgy, ru_wi);

  wire n8irj40n9ts5751 = k7w9hbbfq2amb & (~l2qiuit0jdaq2pbqot);
  wire afnouqeb8x1hrs_sjb1qx7q6 = v3ov4l_sfrqtd5gzo;
  wire l6ibn0emgp5ac27srn781jyqp8l;
  wire tu7pvnivwufqidxxqmpperpwks;
  wire uo358iz6xto41i2v7gdartvmtc = t1y5bixqb70xoxpulhmy;

  assign fppz16b2vnxcgbxo5flw_ni5a = n8irj40n9ts5751 ? 1'b0 : hxhn_tu5eqc44_0avu;

  ux607_gnrl_fifo # (
      .DP (4),
      .DW (1)
  ) k2cgh_scg4vicfxqvs1yyxallivmy6n(
    .i_vld  (afnouqeb8x1hrs_sjb1qx7q6),
    .i_rdy  (l6ibn0emgp5ac27srn781jyqp8l),
    .i_dat  (h3tgasjwjf9pjoc3uvwxw),
    .o_vld  (tu7pvnivwufqidxxqmpperpwks),
    .o_rdy  (uo358iz6xto41i2v7gdartvmtc),  
    .o_dat  (l2qiuit0jdaq2pbqot),  
    .clk    (gf33atgy),
    .rst_n  (ru_wi)
  );

  wire [nm_fj-1:0] i00quc3x43h;
     
     
     
  wire o5c5y3dn  = v3ov4l_sfrqtd5gzo & ( j1rvopf2x3yuqsb);
     
  wire j5a0kqjm6c3  = v3ov4l_sfrqtd5gzo & (~j1rvopf2x3yuqsb);
  wire qwiej1nsik  = o5c5y3dn | j5a0kqjm6c3;
  
  wire [nm_fj-1:0] fh_yhpdb9y4uv = ({i00quc3x43h[nm_fj-1:2],2'b0} + {{nm_fj-4{1'b0}},4'd8});
 
 
 
  wire [nm_fj-1:0] ur3nmlo0dzzyz = o5c5y3dn ? {aw0a19a967dn7n0x25w[nm_fj-1:2],2'b0} : fh_yhpdb9y4uv;
  ux607_gnrl_dfflr #(nm_fj) c3x_7a0gzdh083r (qwiej1nsik, ur3nmlo0dzzyz, i00quc3x43h, gf33atgy, ru_wi);

  wire f5yetvw_f7;
  wire e6scnj06m;

  wire l0npdj_cus6 = ty6a2k41y0e9ir8_yzg;
  wire bspkaws1evi = cwkq4r6_upg_2884r;

  wire w9w0t4t_5bw_h = o5c5y3dn;
  wire wgtzfsvtcij = o5c5y3dn;

  ux607_gnrl_dfflr #(1) vcj5axt7oqxq (wgtzfsvtcij, bspkaws1evi, e6scnj06m, gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1) dvhkwlqft931uz (w9w0t4t_5bw_h, l0npdj_cus6, f5yetvw_f7, gf33atgy, ru_wi);

  assign ui2ziibknh_1uaiixo0m1  = j1rvopf2x3yuqsb ? aw0a19a967dn7n0x25w  : fh_yhpdb9y4uv;
  assign kpptfyyykyfkwr_w7zz = j1rvopf2x3yuqsb ? cwkq4r6_upg_2884r : e6scnj06m;
  assign mqdln_zof0pm8dvg2cb_e = j1rvopf2x3yuqsb ? ty6a2k41y0e9ir8_yzg : f5yetvw_f7;
     
  assign oz7xvqjtmxw3yf4j3 = j1rvopf2x3yuqsb ? air1drtzqvyz1ydvdej : 1'b0;

  wire h2j202k2_h2;
  wire iqzc91c0a5f4 = s4_gwe0uskrbhp37ksb;
  wire tbd6yrxrp05 = o5c5y3dn;
  ux607_gnrl_dfflr #(1) iqn10kmwrodxpt (tbd6yrxrp05, iqzc91c0a5f4, h2j202k2_h2, gf33atgy, ru_wi);
  assign ll0zpg0jpkuqhp9f55h = j1rvopf2x3yuqsb ? s4_gwe0uskrbhp37ksb : h2j202k2_h2;

  wire zu5fzjwuao;
     
  wire vf6dvepfgo8uze = o5c5y3dn;
  wire nlvo362fup12 = vf6dvepfgo8uze;
  wire spi33jrk_u679k = vf6dvepfgo8uze;
  ux607_gnrl_dfflr #(1) wnkluf1qndbll48 (nlvo362fup12, spi33jrk_u679k, zu5fzjwuao, gf33atgy, ru_wi);

  
  
      
  
   
   
   
  
  
  
  wire jmfbolc77xbjjchjuk = (j1rvopf2x3yuqsb ? 1'b1 : bo4tz80rb2i3jzf7tz05t39) & l6ibn0emgp5ac27srn781jyqp8l;
  wire wpo33yfzo3tcd3ake9vdmwr = j1rvopf2x3yuqsb ? kcv48ukn4yb7uxlfz_l76v6 : zu5fzjwuao;
  wire w5zp09nvor1u7f9flxey8tzb2r = vlhrtmmnzbn11e0gw;
  assign q9uknlmu4747layzj7   = jmfbolc77xbjjchjuk & wpo33yfzo3tcd3ake9vdmwr;
  assign ab3stth5phu3zhxwjv1re = jmfbolc77xbjjchjuk & w5zp09nvor1u7f9flxey8tzb2r;

  assign bf61lpqg8z = 
                      tu7pvnivwufqidxxqmpperpwks 
                    | st7pytysu10a
                    | q9uknlmu4747layzj7 
                    | hxhn_tu5eqc44_0avu
                    | c52ldkop361ts52m0 
                    | v9ov1b3vn5k4ctkb 
                    | ult8a6a0b4agydwsws 
                    ;
      
  assign ny26eoy00tenwa = (~bf61lpqg8z);
      


endmodule

















module p651q_8n0fzsut5za #(
    parameter onr7l = 32,
    parameter mhdlk = 4
)(
   input  u22pp,
   input  irka0,
   input  [onr7l-1:0] qbjvs30wtb,
   output [onr7l-1:0] dqgck5s,
   output [onr7l*mhdlk-1:0] pc6rgvhuc_wry1q,
   output [mhdlk-1:0] ks96miyn2gm4,
   output [mhdlk-1:0] lexmfixlro03vle63iq,

   input  mhilu6fd3fe,
   input  [mhdlk-1:0] u60e_km0nn,
   input  [mhdlk*onr7l-1:0] vjgphsh5tfo,

   input  gf33atgy,
   input  ru_wi
);


  wire [onr7l-1:0] olf4xmxku9u9k8 [mhdlk-1:0];
  wire [mhdlk-1:0] cryhplg9_24tqw;
  wire [onr7l-1:0] d82dflwp06cax_ [mhdlk-1:0];



  wire [mhdlk-1:0] uipdtjs;
  wire [mhdlk-1:0] acm0zbhvam;
  wire [mhdlk-1:0] oi40qurrxr; 
  wire [mhdlk-1:0] n89fv;

  wire jlo7_b_z = (irka0 ^ u22pp) | mhilu6fd3fe;
  assign oi40qurrxr = mhilu6fd3fe ? u60e_km0nn :
                   irka0 ? (n89fv[0] ? {1'b1,{mhdlk-1{1'b0}}} : (n89fv >> 1)) :
                           (n89fv[mhdlk-1] ? {{mhdlk-1{1'b0}},1'b1} : (n89fv << 1))
                         ;  

  ux607_gnrl_dfflrs #(1)    svv3sz17bdpp(jlo7_b_z, oi40qurrxr[0]     , n89fv[0]     , gf33atgy, ru_wi);
  ux607_gnrl_dfflr  #(mhdlk-1) o0mc8mg4cq9iqbw(jlo7_b_z, oi40qurrxr[mhdlk-1:1], n89fv[mhdlk-1:1], gf33atgy, ru_wi);


  assign uipdtjs = n89fv; 
  assign acm0zbhvam = (n89fv == {{mhdlk-1{1'b0}},1'b1}) ? {1'b1, {mhdlk-1{1'b0}}}
                                                : (n89fv >> 1); 
  assign lexmfixlro03vle63iq = oi40qurrxr;                             
  assign ks96miyn2gm4 = n89fv;                                                

  genvar i;
  generate 

    for (i=0; i<mhdlk; i=i+1) begin:eyoclcjcy41
      assign cryhplg9_24tqw[i] = (u22pp & uipdtjs[i]) | mhilu6fd3fe ;      
      assign d82dflwp06cax_[i] =  mhilu6fd3fe ? vjgphsh5tfo[onr7l*(i+1)-1:onr7l*i] 
                                        : qbjvs30wtb;
      assign pc6rgvhuc_wry1q[onr7l*(i+1)-1:onr7l*i] = olf4xmxku9u9k8[i];
      ux607_gnrl_dfflr  #(onr7l) s3y1py6je3tms (cryhplg9_24tqw[i], d82dflwp06cax_[i], olf4xmxku9u9k8[i], gf33atgy, ru_wi);
    end
  endgenerate


  integer j;
  reg [onr7l-1:0] ui9y38d1t;
  always @*
  begin : e82692n5bc4eh
    ui9y38d1t = {onr7l{1'b0}};
    for(j=0; j<mhdlk; j=j+1) begin
      ui9y38d1t = ui9y38d1t | ({onr7l{acm0zbhvam[j]}} & olf4xmxku9u9k8[j]);
    end
  end

  assign dqgck5s = ui9y38d1t;

endmodule



















module m1691tbt1_d8b0d7avy69zn(
    input  n38s98n2ak7rvsds, 
    input  vncx4r8ansja, 
    input  w2jm73vsinhrawnk, 
    input [64-1:0] k2mmowd1vvq, 

    output [4-1:0] yddzpj5oad_dtepf,

    input gf33atgy,
    input ru_wi
);

































































  wire ty8m7nbkz9fhzegl = (k2mmowd1vvq[2:1] == 2'b0);
  wire y6yo9bz5y7x7v4 = ~ty8m7nbkz9fhzegl; 
  wire pywe6mcdv1jxh5bj88m3h = n38s98n2ak7rvsds & y6yo9bz5y7x7v4 & (~vncx4r8ansja) & (~w2jm73vsinhrawnk) & (k2mmowd1vvq[2:1] == 2'b11);

  assign yddzpj5oad_dtepf[0]    = pywe6mcdv1jxh5bj88m3h;
  assign yddzpj5oad_dtepf[1]      = n38s98n2ak7rvsds & ty8m7nbkz9fhzegl & (~(vncx4r8ansja & w2jm73vsinhrawnk));

  assign yddzpj5oad_dtepf[2]    = n38s98n2ak7rvsds & y6yo9bz5y7x7v4 & (~pywe6mcdv1jxh5bj88m3h);

  assign yddzpj5oad_dtepf[3] = (~n38s98n2ak7rvsds) & y6yo9bz5y7x7v4;



endmodule 



















module w3yn55ly7roq (
  output c4ughu0qm5sfai,


  input tw5xnp59d8x,
  input aw82i964do,
  input y8_gkxsfle,
  input pydatzxqqi,

  output h8xul8_er09on,

  input  [64-1:0] wd9dvepxj,  

















































  output x0i6aykuzxn1t7_hyw9s7r4to, 
  input  pbyudse8quydhisrzo9pbl4, 
  output [16-1:0]   vapgj050raiah87lnzt_a, 
  output cvksl3f95u8b10a3rmr6qvom,
  output togorwkvhfveb6zwndvww,
  output i036i6j05gm5ht39aak7k, 
  output xubhke6y45gk7d9bj7c1022icq,
  output nao0kbyh1yex0kg7uycyc,

  input  c8u60qjfyfel53grl6lmf5_3, 
  input  vhl77l_vrkmhgbq9nx8p8ix,   
  input  [64-1:0] sedkfhar7baq5_wmvydzjmit2, 
  input  sf4u33sbbh0akueinpc6j4ly8ue,   



  input  s7eq8f6z1uyi2in   ,
  input  w92a5o09fp9dg6   ,
  input  ous_emkpecrqhg5e7,
  input  qbsr1jytrqtsbk4ttb8nz,

  input  svlxg92fk8wh7_jgsa8x,

  output                           ldqpjrsj9dp8yg3uc,  
  output                           s70e4xdis3p67ndpn6fbx,  
  output [7-1:0] h9zlka3j3ih8ihpvwvky1, 
  
  output [54-1:0] tf_tmpul8i8qbm_djvtl5f,
  input  [54-1:0] qtsqtuxyont41a7h7i6,

  output                           w0ve66vjdz8lzwws3ic,  
  output                           df775k2ts6dn4528iq_ce5,  
  output [9-1:0] k3dychuj1pv4vw7cfj01ft8v, 
  
  output [64-1:0] jh4zf96qrsb31j072n,         
  input  [64-1:0] vfvtxk4jkkc3ql7_rqd,

  output                           hv6xxz3oswj4wy4j46,  
  output                           q6p7kcdd9o7j3e2c886,  
  output [7-1:0] ee_yaeclihal4dht69liwy6z, 
  
  output [54-1:0] thl4cxcuzntax8hnsn9bl4,         
  input  [54-1:0] mysqpp41yovfcis6f2dza47,

  
  output                           vp3x08mx4e27x4k26n,  
  output                           a7b829uahvy2i28yzgg,  
  output [9-1:0] kzxrmeg90fb06oya08h1, 
  
  output [64-1:0] kl5wycr14v5ukl7oqfhwe6,         
  input  [64-1:0] wt6c82_zmqgmt7if41t698,


  input  i_x3a8jgmo8qd81tcr,


  output wz_if_2q_23jhl2,
  input  n1wslu68m9v,

  output  x27lqkgq55knwoqsc6_bn0p, 
  input   ud5ygg9b8pmm93drtbfk4l8hv,
  output  [64-1:0] f_lrqmtz5mpqmbrhn6f05, 
  output  czjipv9hqkdx4jllt3ajsl,
  output  j92g3e8ublsg2d9sjj_i3,
  output  af3a5ot65per6f87crwmj, 
  output  bjucsszqg5d1sc5etnwvf1, 
  output  t37flu99i5ex1j3e_8   , 
  output  ss92bd8t5gyfjfl1_lp2,
  output  [2:0] z1beclu7k0_h4nn6njz05sbe1,
  output  [1:0] w1i6s2iwu2nnj7idywd,
  output  [1:0] wvjkzp74fi8ed7nnr7xlm3gt,

  input   phzkntckzzbndu4wevf1o6, 
  input   bpyef3a0dnkkyqdpymy, 
  input   [64-1:0] ba1ucnyekcm68i9wuqwmn,


  output bf61lpqg8z,
  input  dnl01g_,

  
  
  
  output  j8cjhcuf0m6xjvemdaz, 
  output  umc_2tn6um_9xaiy7_ksg0w,
  output  uiyh4da4134sjv7gnmc,
  output  q7ru87fmzxczveihcxcwh, 
  input   s_eowfyzlvx7gjv542upo,


  
  
  
  output d40pep591l63yhmefp7i,

  output t57d026x085pay,
  input  k5th293qdrtsytaehbsk,
  output g6gwjq519o1w1m3csgrrf3,
  output [27-1:0] lo_2ny7_v71by78q3,
  output hbdj3fcr8qkfkgzq58o1o2ozh,
  output [16-1:0] m_k_n75bb0f_im9fu_,




  input ozt73ngxbaqnefsu,

  output m6dcbta00ca03,
  output [32-1:0] c06dvphgeptbqa,
  output t2e9t5kf8lqaa82dtg,
  output viaoqex1en8ydnwh5,
  output st9v6ljxhtiqln7,
  output [5-1:0] sehjrvl7lsqlkpl8js,
  output [5-1:0] owbvtem77_l_b4,
  output [5-1:0] crywtg_a3ctx3707n,

  output                         h9zak9fmm8rw ,   
  output                         xvhg384tm4h76gdzx ,   
  output                         hdlty51ir9snk3qql9ow ,   
  output                         e0bgl8ntt8sp5j7o1yo ,   
  output                         ifg_e4rrluhhouqgceuo2,   
  output                         sz1c6k4c7y75fhzt1m81q,   
  output                         y_g5vz_1yjpqe371ks,  
  output [5-1:0] y88swlv8vqatvrurk392,
  output [5-1:0] yx32lmcp5paz31u5hecbq,
  output [5-1:0] pktjjlrrkgnqgrqag,


  output [32-1:0] z0o61mxkm788c,
  output [64-1:0] pm7xlj7bu,   
  output bcv5wwa3cpmh6o9d, 
  output pbiupof7z_siv68x2, 
  output eey8q1ex7jqqx0hm_,
  output hyzfgvg8iynh8zpa4,
  output mdfkn7idoni9xj,                  
  output v3pirqtitn2_xu9,                   
  output n0p5652lvx0qj1yuwu,               
  output ddp4_khmuujfs,                   
  output m_7gx91ep6vkla,                   
  output iyoccmh9a_a2ov94o,                 
  output [5-1:0] s8mlhtj2pe58l,
  output [5-1:0] eh7xldx93qn_e_ig,
  output [5-1:0] mxxfa5sn2ahc21k,
  output                         wp3ochi2x8_ljvjh,
  output                         yzl1nx341x5d2p4,
  output                         l11qpt1sf6a7,
  output n3mz6a4lr36ftz11,               
  output [64-1:0] f2d4k4kxynjpd0gghqe140, 
  output [4*8-1:0] uuy2zpbrzrwdf432a7_g,
  input  [4*8-1:0] d4d7ru_yllps7en_tto,
  output [7:0] ylmhlw32ex4fxli7,
  input  [7:0] n_lam8gs1mljgiq8zi,
  output [2:0] v_97hsna5xll5n1xslwe3,
  input  [2:0] v2r90qa11qssvr5tq98dbi961,
  output ba89afyz0al00,
  input  gkonom22e0fpa2_v3w0ab,
  output [2-1:0] fxvpc9o9zl2t2nuwpg0,
  input  [2-1:0] gtvau5cygdmb10dr_makqf,
  output qu31vl4s4x0pmeth2j_7neq1,
  output himvp4q0erus0anat5,               
  output ps9l2wesoladg,
  output yoo3wc2tlwfyc6, 
  input  f78zm1o77tcsokzo,

  input  hwpkcsh2atrq  ,
  input  v3e6l1k7eo9k3 ,
  input  hxrmt706n071lic0f7,
  input  v7rzl8qveorn2jg6659m69,
  input  v_k8ohy_e2e9vlp6az04,
  input [64-1:0] y_vw514j6xmphhfhc,
  input [9-1:0] p54semfzu2zyfb,
  output [9-1:0] xosc7587i2hjow2yjw,
  output  zsgl59ydqwjln,
  input   b9yq2alidby7zgom1,


  input   [64-1:0] h01d94xsxbxe_req,  
  input   tvqijouldcgiz2dxdco7,  
  input   zkxlkidschdubxpkpm,  
  input   xmcrni1qngfvh9pil9j,  
  input   btkcf2uqr61gkiqhde0lai,  
  input   w1casjl7bz73brz,
  input   hjri7cufo9ckntq,  
  input   yghffofulqa77bd7aw07badta1a,
  input   rrl7evvmayt1_vvp74iq9h6_cjf,
  input   [27-1:0] zddoxp22m1o11x30gbe,
  input   [16-1:0] hwfethpzkuauejcgtbl6o,  

  output  n3ak8l6cvn0s4,
  input   hsxh9536ho4bw8o,
  input   [64-1:0] jkzw_f9anx55,  
  input   r_edve7v9jcr26q6zk,  
  input   vrqfzuog2k4pos133,  
  input   bmw2yi333716crywk,  
  input   k2sr7sw1plcmnki5ajtscw,  
  input   t8muv9e6d7yk_whqa0,
  input   hzdfp71n6g3f5fsg5,  
  input   lwdhmuzyvcvv14mjbl0h2a41z,
  input   xy48dugh009wtmazqug3kpy2a5h_,
  input   [27-1:0] l4ztejmt2__wxqm2rw,
  input   [16-1:0] s3ujdp2a8n69bm6engxok,  






  input  p0olq02_hyvx0,
  output mneths0pu5slsnpiv,

  input q97rqfy8n7ixfm2a5wev4nd5sylpcq3j,
  input lln3b7iev7jpvogh964ro_9bc_3y,
  input hujgg6hjnhtbspbkekuz5_u,
  input v3pnt81kfrgbaanm1mhh51w,
  input [64-1:0] i08eq60d_snxeq8si_ezod,
  input dgnjyd9xs8efyxm0tdlsvfq4eop,
  input y8wz7aud_fd6dfiakjtx2i0g,
  input a3xib90kwk4_hm1,
  input nfzexr8q9g893gi,
  input [64-1:0] opkkwp3eg8g3448t,

  input  um28jgd2x4mbs,
  input  [64-1:0] l_imk5zs8ejjka,
  input  [64-1:0] lz3vnoxnz_z,
  input  yhbtmo4kyz_ewog3,
  input  cd4d2_i3rcc1_p,
  input  [5-1:0] wyu42gj62n994v0wo_,
  input  x9cmkt53yq483z1,
  input  cxmwxfttqy2t7ura   ,
  input  b5wruck8tj9sa   ,
  input  bxentpryfwb3d  ,
  input  o2a43mjdbgea1  ,
  output enwn0u48p2_ls5az80,
  output miax48k27o484e8a,
  input [8*32-1:0] pcr4upio7_tx37, 
  input [8*1-1:0] uzklqlncpqqm1rav,
  input [8*1-1:0] ortueunvnkx_l5m_j,
  input [8*1-1:0] hwuhtb7ucto_utk56,
  input [8*2-1:0] i1env2kmns7qvvuuc,
  input [8*1-1:0] g3s3vpafvy3i,


  
  
  
  input                                    e1jv60iid34gonwyukkue,           
  input  [74-1:0]       xz57o2ko5gkcbk8rq,          
  output                                   grv8y38uxakr22asia,         
  output                                   bvmb0d5jendar95w7nbnob8,           
  output [5:0]                             h47i__o10wyo2sbyt58zq1_h5,      

  
  
  
  input                                    vxwhhz9_cff6uy0x,
  
  output                                   moj77icm1kmex0900,                
  output  [27-1:0]     hib0x0rvcjwnn75a,                 
  output  [1:0]                            cgmsm8wvxc5kg90xwvwq0cga,                 
  
  input                                    w9mx37ezcezieq_9__94o,          
  input                                    hsnr3xtposirc7pmphtiko3xlz,     
  input                                    k1jkhgd9bvypwrti7ietjp0n7_nyzu,   
  input  [51-1:0]       qirelbyt49gkn46_f24yxtc,           
  input                                    jq4wiwydrozelhpru9snvs0,         
  input                                    j6muxslh7pud3298q9d8lc2,         

  input  gc4b3kdcan6do88ta_,
  input  o5q5hev,
  input  ru_wi
  );

  wire jnq99nw1wv9zocbz; 
  wire sj1gaizva5__by20e; 
  wire [64-1:0]   k2mmowd1vvq; 
  wire zc2e7csnzgj98szggj;
  wire ih_5pl6hw4ippiu;
  wire y4vtwevsvl03ho6h0;
  wire hto4un7x8fe6gc1;
  wire [4-1:0] agsse3cpfshpa0xh48nu0;
  wire n38s98n2ak7rvsds;
  wire vncx4r8ansja;
  wire w2jm73vsinhrawnk;
  wire p_xqcszydp2j5d821j; 
  wire ht929tfpovwde; 
  wire mkytk1e8mwi49l;   
  wire xr81_h9hnhjwec3la;   
  wire tbs7se44h1m47t;   
  wire krxdptqk3busoihx2f;   
  wire gnmzf7svwij0ih7c7fh3;   
  wire we422ti7i_fjt8z36n53;   
  wire tylsyqg3frnshrlcfkd596;   
  wire rk6m6hfluv6syr3pz6z;   
  wire eygoo8ifqdnay_dhiskf_;   
  wire xfxeg_cwdrq6mzr3teo;   
  wire diw3rbg3tca7kp6uu3l2n;   
  wire [32*2-1:0] m9u9kwx2_i51v; 


  wire ny26eoy00tenwa;

   wire f48_2zc1qro_3dodmk8 ;
   wire vaiscz5bqo4k6ql0519 ;
   wire w93is2iaq5aikcpaqxg3 ;
   wire uuuoq6te8sq6lj_e02iqoc ;
   wire azqy5qfm4kwm7vkwu6e;
   wire ig7796duzb8wqodp;

   wire qmd94avv02av64cbwaj42 ;
   wire hv9e7_hu5oyc6e87832pmb;
   wire m4ndmqnlr5eisc8m2k6fd;
   wire [27-1:0] jcczlhzxqzl5dx51l;
   wire nkdn__tk5pvp4nczp7xysy5;
   wire [16-1:0] fhzpp1p52pmfd3syoo;


  wire azm2vbkop_ll3;
  wire e8xevpvl7622ut;
  wire eb506yrftyyi;

  wire v4gayo0h8l6na;
  wire [64-1:0] nmy2nw74r7gg;
  wire ag7oznqt1davxt_ateix = aw82i964do;
  wire crissrnil1b81y9i4z5b = y8_gkxsfle;
  wire lff9k60vjdno23w3j = pydatzxqqi;
  wire kqepyrf26fkyy4nfbcb = 1'b0;
  wire hel4fu2nnjoq7fo5ajmx = 1'b0;
  wire mosnaiams7ws78b = 1'b0;
  wire v68_c8wty40tt9fiw7wr4126 = 1'b0;
  wire k0h81we1ir7v14ih_2h_ke4_ugx = 1'b0;
  wire [27-1:0] ok5b5bmabu8sw54j1dp = 27'b0;
  wire [16-1:0] awg6_wgvi09fsrjdjapqluj_m = 16'b0; 
  wire w2iw_tnc6hjryhl0x99;
  assign zsgl59ydqwjln = w2iw_tnc6hjryhl0x99;
  wire y3z3zpxfgxrbx38 = v4gayo0h8l6na | b9yq2alidby7zgom1;
  wire g5yf_4_mik =  b9yq2alidby7zgom1 | hsxh9536ho4bw8o;
  wire [64-1:0] g6ixtnv0p9i7t56z =  b9yq2alidby7zgom1 ? h01d94xsxbxe_req : nmy2nw74r7gg;
  wire pykis3m72999nbat1vr3i3s =  b9yq2alidby7zgom1 ? tvqijouldcgiz2dxdco7 : ag7oznqt1davxt_ateix;
  wire nx3fumqniblb3n80s0j99 =  b9yq2alidby7zgom1 ? zkxlkidschdubxpkpm : crissrnil1b81y9i4z5b;
  wire yp1uv8hz44sr7lcp0d9g8s =  b9yq2alidby7zgom1 ? xmcrni1qngfvh9pil9j : lff9k60vjdno23w3j;
  wire gsr_eo06m498skevdwc5 =  b9yq2alidby7zgom1 ? btkcf2uqr61gkiqhde0lai : kqepyrf26fkyy4nfbcb;
  wire nf0tdr1088vkc3n337km = b9yq2alidby7zgom1 ? w1casjl7bz73brz : hel4fu2nnjoq7fo5ajmx;
  wire bcy930rdd3kchj6zz25          = b9yq2alidby7zgom1 ? hjri7cufo9ckntq                   : mosnaiams7ws78b;
  wire swj1ts__7_b_1ty7m6npb47x7   = b9yq2alidby7zgom1 ? yghffofulqa77bd7aw07badta1a   : v68_c8wty40tt9fiw7wr4126;
  wire bi9aryftwbjsj2lmk6_15fkfoa9mdau1 = b9yq2alidby7zgom1 ? rrl7evvmayt1_vvp74iq9h6_cjf : k0h81we1ir7v14ih_2h_ke4_ugx;
  wire [27-1:0] otat8qurqhuymsh77h3nqv   = b9yq2alidby7zgom1 ? zddoxp22m1o11x30gbe   : ok5b5bmabu8sw54j1dp;
  wire [16-1:0]    snmuzlxp_djsvf0z4gtma23 = b9yq2alidby7zgom1 ? hwfethpzkuauejcgtbl6o : awg6_wgvi09fsrjdjapqluj_m; 
  f5fy2w73p7p_y5b   uh9o5ee_7d8aky56swv(
    .nupfecm_6ycs   (),
    .wd9dvepxj      (wd9dvepxj),  
    .jnq99nw1wv9zocbz (jnq99nw1wv9zocbz),
    .sj1gaizva5__by20e (sj1gaizva5__by20e),
    .k2mmowd1vvq    (k2mmowd1vvq   ),
    .zc2e7csnzgj98szggj (zc2e7csnzgj98szggj),
    .ih_5pl6hw4ippiu (ih_5pl6hw4ippiu),
    .y4vtwevsvl03ho6h0 (y4vtwevsvl03ho6h0),
    .hto4un7x8fe6gc1 (hto4un7x8fe6gc1),
    .agsse3cpfshpa0xh48nu0 (agsse3cpfshpa0xh48nu0),
    .n38s98n2ak7rvsds     (n38s98n2ak7rvsds     ),
    .vncx4r8ansja     (vncx4r8ansja),
    .w2jm73vsinhrawnk     (w2jm73vsinhrawnk),

    .p_xqcszydp2j5d821j (p_xqcszydp2j5d821j),
    .ht929tfpovwde (ht929tfpovwde),
    .mkytk1e8mwi49l(mkytk1e8mwi49l  ),
    .xr81_h9hnhjwec3la(xr81_h9hnhjwec3la  ),
    .tbs7se44h1m47t   (tbs7se44h1m47t  ),
    .krxdptqk3busoihx2f(krxdptqk3busoihx2f),
    .gnmzf7svwij0ih7c7fh3(gnmzf7svwij0ih7c7fh3),
    .we422ti7i_fjt8z36n53(we422ti7i_fjt8z36n53  ),
    .tylsyqg3frnshrlcfkd596(tylsyqg3frnshrlcfkd596  ),
    .rk6m6hfluv6syr3pz6z(rk6m6hfluv6syr3pz6z  ),
    .eygoo8ifqdnay_dhiskf_(eygoo8ifqdnay_dhiskf_  ),
    .xfxeg_cwdrq6mzr3teo(xfxeg_cwdrq6mzr3teo),
    .diw3rbg3tca7kp6uu3l2n(diw3rbg3tca7kp6uu3l2n),
    .m9u9kwx2_i51v (m9u9kwx2_i51v),

    .azm2vbkop_ll3  (azm2vbkop_ll3),
    .e8xevpvl7622ut    (e8xevpvl7622ut),
    .eb506yrftyyi    (eb506yrftyyi),

    .enwn0u48p2_ls5az80   (enwn0u48p2_ls5az80),
    .miax48k27o484e8a   (miax48k27o484e8a),

    .m6dcbta00ca03    (m6dcbta00ca03    ),
    .rnx27onf2lbe    (ozt73ngxbaqnefsu    ),
    .c06dvphgeptbqa    (c06dvphgeptbqa    ),
    .t2e9t5kf8lqaa82dtg(t2e9t5kf8lqaa82dtg),
    .viaoqex1en8ydnwh5(viaoqex1en8ydnwh5),
    .st9v6ljxhtiqln7(st9v6ljxhtiqln7),
    .sehjrvl7lsqlkpl8js(sehjrvl7lsqlkpl8js),
    .owbvtem77_l_b4(owbvtem77_l_b4),
    .crywtg_a3ctx3707n(crywtg_a3ctx3707n),
    .h9zak9fmm8rw       (h9zak9fmm8rw       ),   
    .xvhg384tm4h76gdzx (xvhg384tm4h76gdzx ),   
    .hdlty51ir9snk3qql9ow (hdlty51ir9snk3qql9ow ),   
    .e0bgl8ntt8sp5j7o1yo (e0bgl8ntt8sp5j7o1yo ),   
    .ifg_e4rrluhhouqgceuo2(ifg_e4rrluhhouqgceuo2),   
    .sz1c6k4c7y75fhzt1m81q(sz1c6k4c7y75fhzt1m81q),   
    .y_g5vz_1yjpqe371ks(y_g5vz_1yjpqe371ks), 
    .y88swlv8vqatvrurk392(y88swlv8vqatvrurk392),
    .yx32lmcp5paz31u5hecbq(yx32lmcp5paz31u5hecbq),
    .pktjjlrrkgnqgrqag(pktjjlrrkgnqgrqag),
    .z0o61mxkm788c      (z0o61mxkm788c     ),
    .pm7xlj7bu  (pm7xlj7bu     ),
    .bcv5wwa3cpmh6o9d(bcv5wwa3cpmh6o9d),
    .pbiupof7z_siv68x2(pbiupof7z_siv68x2),
    .eey8q1ex7jqqx0hm_(eey8q1ex7jqqx0hm_),
    .hyzfgvg8iynh8zpa4  (hyzfgvg8iynh8zpa4 ),
    .mdfkn7idoni9xj (mdfkn7idoni9xj),
    .v3pirqtitn2_xu9  (v3pirqtitn2_xu9 ),
    .n0p5652lvx0qj1yuwu  (n0p5652lvx0qj1yuwu ),
    .ddp4_khmuujfs  (ddp4_khmuujfs ),
    .m_7gx91ep6vkla  (m_7gx91ep6vkla ),
    .iyoccmh9a_a2ov94o(iyoccmh9a_a2ov94o),
    .s8mlhtj2pe58l  (s8mlhtj2pe58l),
    .eh7xldx93qn_e_ig  (eh7xldx93qn_e_ig),
    .mxxfa5sn2ahc21k  (mxxfa5sn2ahc21k),
    .wp3ochi2x8_ljvjh   (wp3ochi2x8_ljvjh ),
    .yzl1nx341x5d2p4   (yzl1nx341x5d2p4 ),
    .l11qpt1sf6a7   (l11qpt1sf6a7 ),
    .n3mz6a4lr36ftz11     (n3mz6a4lr36ftz11),
    .f2d4k4kxynjpd0gghqe140    (f2d4k4kxynjpd0gghqe140),
    .uuy2zpbrzrwdf432a7_g   (uuy2zpbrzrwdf432a7_g),
    .d4d7ru_yllps7en_tto   (d4d7ru_yllps7en_tto),
    .ylmhlw32ex4fxli7       (ylmhlw32ex4fxli7       ),
    .n_lam8gs1mljgiq8zi       (n_lam8gs1mljgiq8zi       ),
    .v_97hsna5xll5n1xslwe3  (v_97hsna5xll5n1xslwe3),
    .v2r90qa11qssvr5tq98dbi961(v2r90qa11qssvr5tq98dbi961),
    .ba89afyz0al00        (ba89afyz0al00        ),
    .gkonom22e0fpa2_v3w0ab     (gkonom22e0fpa2_v3w0ab     ),
    .fxvpc9o9zl2t2nuwpg0    (fxvpc9o9zl2t2nuwpg0    ),
    .gtvau5cygdmb10dr_makqf    (gtvau5cygdmb10dr_makqf    ),
    .qu31vl4s4x0pmeth2j_7neq1(qu31vl4s4x0pmeth2j_7neq1),
    .himvp4q0erus0anat5     (himvp4q0erus0anat5),
    .ps9l2wesoladg           (ps9l2wesoladg),
    .yoo3wc2tlwfyc6          (yoo3wc2tlwfyc6  ),
    .f78zm1o77tcsokzo          (f78zm1o77tcsokzo  ),
    .hwpkcsh2atrq  (hwpkcsh2atrq  ),
    .v3e6l1k7eo9k3 (v3e6l1k7eo9k3 ),
    .hxrmt706n071lic0f7(hxrmt706n071lic0f7),
    .v7rzl8qveorn2jg6659m69 (v7rzl8qveorn2jg6659m69),
    .v_k8ohy_e2e9vlp6az04   (v_k8ohy_e2e9vlp6az04),
    .y_vw514j6xmphhfhc (y_vw514j6xmphhfhc),
    .p54semfzu2zyfb    (p54semfzu2zyfb   ), 
    .xosc7587i2hjow2yjw    (xosc7587i2hjow2yjw   ), 
    .v4gayo0h8l6na     (v4gayo0h8l6na    ),
    .nmy2nw74r7gg      (nmy2nw74r7gg     ),
    .zsgl59ydqwjln     (w2iw_tnc6hjryhl0x99    ), 
    .b9yq2alidby7zgom1     (y3z3zpxfgxrbx38    ),


    .g5yf_4_mik         (g5yf_4_mik),
    .h01d94xsxbxe_req      (g6ixtnv0p9i7t56z),  
    .w1casjl7bz73brz  (nf0tdr1088vkc3n337km),
    .hjri7cufo9ckntq          (bcy930rdd3kchj6zz25         ),
    .yghffofulqa77bd7aw07badta1a   (swj1ts__7_b_1ty7m6npb47x7  ),
    .rrl7evvmayt1_vvp74iq9h6_cjf (bi9aryftwbjsj2lmk6_15fkfoa9mdau1),
    .zddoxp22m1o11x30gbe       (otat8qurqhuymsh77h3nqv      ),
    .hwfethpzkuauejcgtbl6o     (snmuzlxp_djsvf0z4gtma23    ),
    .xmcrni1qngfvh9pil9j(yp1uv8hz44sr7lcp0d9g8s),
    .btkcf2uqr61gkiqhde0lai(gsr_eo06m498skevdwc5),
    .tvqijouldcgiz2dxdco7(pykis3m72999nbat1vr3i3s),
    .zkxlkidschdubxpkpm(nx3fumqniblb3n80s0j99),
    .n3ak8l6cvn0s4       (n3ak8l6cvn0s4     ),
    .hsxh9536ho4bw8o       (hsxh9536ho4bw8o     ),
    .jkzw_f9anx55        (jkzw_f9anx55      ),
    .r_edve7v9jcr26q6zk  (r_edve7v9jcr26q6zk),
    .vrqfzuog2k4pos133  (vrqfzuog2k4pos133),
    .bmw2yi333716crywk  (bmw2yi333716crywk),
    .k2sr7sw1plcmnki5ajtscw  (k2sr7sw1plcmnki5ajtscw),
    .t8muv9e6d7yk_whqa0    (t8muv9e6d7yk_whqa0),
    .hzdfp71n6g3f5fsg5          (hzdfp71n6g3f5fsg5),
    .lwdhmuzyvcvv14mjbl0h2a41z   (lwdhmuzyvcvv14mjbl0h2a41z  ),
    .xy48dugh009wtmazqug3kpy2a5h_ (xy48dugh009wtmazqug3kpy2a5h_),
    .l4ztejmt2__wxqm2rw       (l4ztejmt2__wxqm2rw      ),
    .s3ujdp2a8n69bm6engxok     (s3ujdp2a8n69bm6engxok    ),

    .ny26eoy00tenwa  (ny26eoy00tenwa),

    .p0olq02_hyvx0  (p0olq02_hyvx0 ),
    .mneths0pu5slsnpiv  (mneths0pu5slsnpiv ),

    .lln3b7iev7jpvogh964ro_9bc_3y (lln3b7iev7jpvogh964ro_9bc_3y),
    .q97rqfy8n7ixfm2a5wev4nd5sylpcq3j (q97rqfy8n7ixfm2a5wev4nd5sylpcq3j),
    .hujgg6hjnhtbspbkekuz5_u(hujgg6hjnhtbspbkekuz5_u),
    .v3pnt81kfrgbaanm1mhh51w (v3pnt81kfrgbaanm1mhh51w),
    .i08eq60d_snxeq8si_ezod(i08eq60d_snxeq8si_ezod),
    .y8wz7aud_fd6dfiakjtx2i0g (y8wz7aud_fd6dfiakjtx2i0g),
    .dgnjyd9xs8efyxm0tdlsvfq4eop (dgnjyd9xs8efyxm0tdlsvfq4eop),
    .a3xib90kwk4_hm1(a3xib90kwk4_hm1),
    .nfzexr8q9g893gi (nfzexr8q9g893gi),
    .opkkwp3eg8g3448t(opkkwp3eg8g3448t),

    .um28jgd2x4mbs    (um28jgd2x4mbs   ),
    .l_imk5zs8ejjka     (l_imk5zs8ejjka    ),
    .lz3vnoxnz_z    (lz3vnoxnz_z   ),
    .yhbtmo4kyz_ewog3  (yhbtmo4kyz_ewog3 ),
    .cd4d2_i3rcc1_p (cd4d2_i3rcc1_p),
    .wyu42gj62n994v0wo_ (wyu42gj62n994v0wo_),
    .x9cmkt53yq483z1(x9cmkt53yq483z1),
    .cxmwxfttqy2t7ura   (cxmwxfttqy2t7ura   ),
    .b5wruck8tj9sa   (b5wruck8tj9sa   ),
    .bxentpryfwb3d  (bxentpryfwb3d  ),
    .o2a43mjdbgea1  (o2a43mjdbgea1  ),

    .c4ughu0qm5sfai  (c4ughu0qm5sfai),
    .f48_2zc1qro_3dodmk8 (f48_2zc1qro_3dodmk8),
    .vaiscz5bqo4k6ql0519(vaiscz5bqo4k6ql0519),
    .w93is2iaq5aikcpaqxg3(w93is2iaq5aikcpaqxg3),
    .uuuoq6te8sq6lj_e02iqoc(uuuoq6te8sq6lj_e02iqoc),
    .azqy5qfm4kwm7vkwu6e(azqy5qfm4kwm7vkwu6e),
    .ig7796duzb8wqodp   (ig7796duzb8wqodp),
    .qmd94avv02av64cbwaj42      (qmd94avv02av64cbwaj42      ),
    .hv9e7_hu5oyc6e87832pmb     (hv9e7_hu5oyc6e87832pmb     ),
    .m4ndmqnlr5eisc8m2k6fd   (m4ndmqnlr5eisc8m2k6fd   ),
    .jcczlhzxqzl5dx51l       (jcczlhzxqzl5dx51l       ),
    .nkdn__tk5pvp4nczp7xysy5 (nkdn__tk5pvp4nczp7xysy5 ),
    .fhzpp1p52pmfd3syoo     (fhzpp1p52pmfd3syoo     ),
    .ous_emkpecrqhg5e7(ous_emkpecrqhg5e7),
    .s7eq8f6z1uyi2in   (s7eq8f6z1uyi2in),
    .qbsr1jytrqtsbk4ttb8nz   (qbsr1jytrqtsbk4ttb8nz),

    .gf33atgy           (o5q5hev      ),
    .ru_wi         (ru_wi        ) 
  );


  wire l3fd1x5l3xpi3bbwblpsrwwruvvw; 
  wire awh5wdqsak51daa1xam8ipi9;
  wire [64-1:0] r_ktqd4uca5y4b3gnhz03iwd; 
  wire mi8oba8vxuze_93cxrid23bv ;
  wire kya1iiz3vedj6v1ucdydery90b ;
  wire y0ozra0qgen9l9te2u_pqq0bx4a ;
  wire mfxhd3_j98125z7zj4spfnef1m6rw ;


  wire wv8wwd_1gm9_e7vubue9gb29; 
  wire yijhfr84p7xs3yctj1skm24t02_; 
  wire jz08e92smloz0op1zfo3g9ungcnbc;   
  wire crrw2ei1pk6riohtoykjv9qeuen;   
  wire ttqo192f6935w8y576tjxiwa30fd;   
  wire [64-1:0] e45yjvds31b0kqjvsynzmgpf; 



  wire c52ldkop361ts52m0;
  wire x88wat37r_vjsn57a;
  wire [64-1:0]   z3k8ps_o7osj4uosf_6i5;
  wire w8k_3fawz__hfg4mk0mw7g;
  wire i88maxesdvq1fkint66;
  wire rzon56p292pybf35mi_;
  wire jn_zyepkhmn_mdbqe1;
  wire ewekc8h7f7w9i3v;

  wire ult8a6a0b4agydwsws;
  wire gkbxrtlrxlk7_fk4;
  wire bwdpzndejgg3liwep6q_;
  wire glkxypl9rxder9fztnegf6;
  wire qe9n3_xo49nzqdf6gl2rz2j;
  wire [64-1:0] d27a6w261um4big8wy8;


  mu0arb3ch40modhq7 yz6lns_lj8xc109if9_2 (
    .jnq99nw1wv9zocbz (jnq99nw1wv9zocbz),
    .sj1gaizva5__by20e (sj1gaizva5__by20e),
    .k2mmowd1vvq    (k2mmowd1vvq   ),
    .zc2e7csnzgj98szggj (zc2e7csnzgj98szggj),
    .ih_5pl6hw4ippiu (ih_5pl6hw4ippiu),
    .y4vtwevsvl03ho6h0 (y4vtwevsvl03ho6h0),
    .hto4un7x8fe6gc1 (hto4un7x8fe6gc1),
    .agsse3cpfshpa0xh48nu0(agsse3cpfshpa0xh48nu0),
    .n38s98n2ak7rvsds     (n38s98n2ak7rvsds     ),
    .vncx4r8ansja     (vncx4r8ansja),
    .w2jm73vsinhrawnk     (w2jm73vsinhrawnk),

    .p_xqcszydp2j5d821j (p_xqcszydp2j5d821j),
    .ht929tfpovwde (ht929tfpovwde),
    .mkytk1e8mwi49l (mkytk1e8mwi49l  ),
    .xr81_h9hnhjwec3la (xr81_h9hnhjwec3la  ),
    .tbs7se44h1m47t    (tbs7se44h1m47t  ),
    .krxdptqk3busoihx2f(krxdptqk3busoihx2f),
    .gnmzf7svwij0ih7c7fh3(gnmzf7svwij0ih7c7fh3),
    .we422ti7i_fjt8z36n53(we422ti7i_fjt8z36n53  ),
    .tylsyqg3frnshrlcfkd596(tylsyqg3frnshrlcfkd596  ),
    .rk6m6hfluv6syr3pz6z(rk6m6hfluv6syr3pz6z  ),
    .eygoo8ifqdnay_dhiskf_(eygoo8ifqdnay_dhiskf_  ),
    .xfxeg_cwdrq6mzr3teo(xfxeg_cwdrq6mzr3teo),
    .diw3rbg3tca7kp6uu3l2n(diw3rbg3tca7kp6uu3l2n),
    .m9u9kwx2_i51v (m9u9kwx2_i51v),

    .azm2vbkop_ll3 (azm2vbkop_ll3),


    .c52ldkop361ts52m0 (c52ldkop361ts52m0 ),
    .x88wat37r_vjsn57a (x88wat37r_vjsn57a ),
    .z3k8ps_o7osj4uosf_6i5  (z3k8ps_o7osj4uosf_6i5  ),
    .w8k_3fawz__hfg4mk0mw7g (w8k_3fawz__hfg4mk0mw7g ),
    .i88maxesdvq1fkint66 (i88maxesdvq1fkint66 ),
    .rzon56p292pybf35mi_ (rzon56p292pybf35mi_ ),
    .jn_zyepkhmn_mdbqe1 (jn_zyepkhmn_mdbqe1 ),
    .ewekc8h7f7w9i3v   (ewekc8h7f7w9i3v   ), 

    .ult8a6a0b4agydwsws (ult8a6a0b4agydwsws ),
    .gkbxrtlrxlk7_fk4   (gkbxrtlrxlk7_fk4   ),
    .bwdpzndejgg3liwep6q_(bwdpzndejgg3liwep6q_),
    .glkxypl9rxder9fztnegf6(glkxypl9rxder9fztnegf6),
    .qe9n3_xo49nzqdf6gl2rz2j(qe9n3_xo49nzqdf6gl2rz2j),
    .d27a6w261um4big8wy8 (d27a6w261um4big8wy8 ),


    .gf33atgy           (o5q5hev   ),
    .ru_wi         (ru_wi     ) 
  );












  x9ryvjofa0kbj48adfm   f80p1z9rdysrssz3do6(
    .w92a5o09fp9dg6   (w92a5o09fp9dg6   ),
    .ous_emkpecrqhg5e7(ous_emkpecrqhg5e7),
    .vxwhhz9_cff6uy0x    (vxwhhz9_cff6uy0x     ),

    .c52ldkop361ts52m0 (c52ldkop361ts52m0 ),
    .x88wat37r_vjsn57a (x88wat37r_vjsn57a ),
    .z3k8ps_o7osj4uosf_6i5  (z3k8ps_o7osj4uosf_6i5  ),
    .w8k_3fawz__hfg4mk0mw7g (w8k_3fawz__hfg4mk0mw7g ),
    .i88maxesdvq1fkint66 (i88maxesdvq1fkint66 ), 
    .rzon56p292pybf35mi_ (rzon56p292pybf35mi_ ),
    .jn_zyepkhmn_mdbqe1 (jn_zyepkhmn_mdbqe1 ),
    .ewekc8h7f7w9i3v   (ewekc8h7f7w9i3v   ), 

    .ult8a6a0b4agydwsws (ult8a6a0b4agydwsws ),
    .gkbxrtlrxlk7_fk4   (gkbxrtlrxlk7_fk4   ),
    .bwdpzndejgg3liwep6q_(bwdpzndejgg3liwep6q_),
    .glkxypl9rxder9fztnegf6(glkxypl9rxder9fztnegf6),
    .qe9n3_xo49nzqdf6gl2rz2j(qe9n3_xo49nzqdf6gl2rz2j),
    .d27a6w261um4big8wy8 (d27a6w261um4big8wy8 ),





























    .x0i6aykuzxn1t7_hyw9s7r4to(x0i6aykuzxn1t7_hyw9s7r4to),
    .pbyudse8quydhisrzo9pbl4(pbyudse8quydhisrzo9pbl4),
    .vapgj050raiah87lnzt_a (vapgj050raiah87lnzt_a ),
    .cvksl3f95u8b10a3rmr6qvom(cvksl3f95u8b10a3rmr6qvom ),
    .togorwkvhfveb6zwndvww(togorwkvhfveb6zwndvww ),
    .i036i6j05gm5ht39aak7k(i036i6j05gm5ht39aak7k ),
    .xubhke6y45gk7d9bj7c1022icq (xubhke6y45gk7d9bj7c1022icq),
	.nao0kbyh1yex0kg7uycyc(nao0kbyh1yex0kg7uycyc),
	.tw5xnp59d8x(tw5xnp59d8x),
                                                  
    .c8u60qjfyfel53grl6lmf5_3(c8u60qjfyfel53grl6lmf5_3),
    .vhl77l_vrkmhgbq9nx8p8ix  (vhl77l_vrkmhgbq9nx8p8ix  ),
    .sedkfhar7baq5_wmvydzjmit2(sedkfhar7baq5_wmvydzjmit2),
    .sf4u33sbbh0akueinpc6j4ly8ue  (sf4u33sbbh0akueinpc6j4ly8ue ), 
                                                  



    .l3fd1x5l3xpi3bbwblpsrwwruvvw (l3fd1x5l3xpi3bbwblpsrwwruvvw),
    .awh5wdqsak51daa1xam8ipi9 (awh5wdqsak51daa1xam8ipi9),
    .r_ktqd4uca5y4b3gnhz03iwd  (r_ktqd4uca5y4b3gnhz03iwd ),
    .mi8oba8vxuze_93cxrid23bv  (mi8oba8vxuze_93cxrid23bv ),
    .kya1iiz3vedj6v1ucdydery90b  (kya1iiz3vedj6v1ucdydery90b ),
    .y0ozra0qgen9l9te2u_pqq0bx4a  (y0ozra0qgen9l9te2u_pqq0bx4a ),
    .mfxhd3_j98125z7zj4spfnef1m6rw  (mfxhd3_j98125z7zj4spfnef1m6rw ),


    .wv8wwd_1gm9_e7vubue9gb29 (wv8wwd_1gm9_e7vubue9gb29),
    .yijhfr84p7xs3yctj1skm24t02_   (yijhfr84p7xs3yctj1skm24t02_  ),
    .jz08e92smloz0op1zfo3g9ungcnbc   (jz08e92smloz0op1zfo3g9ungcnbc  ),
    .crrw2ei1pk6riohtoykjv9qeuen   (crrw2ei1pk6riohtoykjv9qeuen  ),
    .ttqo192f6935w8y576tjxiwa30fd (ttqo192f6935w8y576tjxiwa30fd),
    .e45yjvds31b0kqjvsynzmgpf (e45yjvds31b0kqjvsynzmgpf),


    .ny26eoy00tenwa  (ny26eoy00tenwa),

    .bf61lpqg8z    (bf61lpqg8z),
    .o5q5hev       (o5q5hev   ),
    .dnl01g_       (dnl01g_   ),
    .ru_wi         (ru_wi     ) 
  );



























































































  gdyqy_u6w0mpgo co871e52ji_6rwj(
     .pp7hxkc1fr9z2qqw    (ous_emkpecrqhg5e7),
     .i_x3a8jgmo8qd81tcr (i_x3a8jgmo8qd81tcr ),
     .nvyp85muxi8p9u1y8brs(svlxg92fk8wh7_jgsa8x),

     .f48_2zc1qro_3dodmk8  (f48_2zc1qro_3dodmk8  ),
     .vaiscz5bqo4k6ql0519(vaiscz5bqo4k6ql0519),
     .w93is2iaq5aikcpaqxg3(w93is2iaq5aikcpaqxg3),
     .uuuoq6te8sq6lj_e02iqoc(uuuoq6te8sq6lj_e02iqoc),
     .azqy5qfm4kwm7vkwu6e (azqy5qfm4kwm7vkwu6e ),
     .ig7796duzb8wqodp    (ig7796duzb8wqodp    ),

     .qmd94avv02av64cbwaj42      (qmd94avv02av64cbwaj42      ),
     .hv9e7_hu5oyc6e87832pmb     (hv9e7_hu5oyc6e87832pmb     ),
     .m4ndmqnlr5eisc8m2k6fd   (m4ndmqnlr5eisc8m2k6fd   ),
     .jcczlhzxqzl5dx51l       (jcczlhzxqzl5dx51l       ),
     .nkdn__tk5pvp4nczp7xysy5 (nkdn__tk5pvp4nczp7xysy5 ),
     .fhzpp1p52pmfd3syoo     (fhzpp1p52pmfd3syoo     ),

     .j8cjhcuf0m6xjvemdaz  (j8cjhcuf0m6xjvemdaz  ),
     .umc_2tn6um_9xaiy7_ksg0w(umc_2tn6um_9xaiy7_ksg0w),
     .uiyh4da4134sjv7gnmc(uiyh4da4134sjv7gnmc),
     .q7ru87fmzxczveihcxcwh(q7ru87fmzxczveihcxcwh),
     .s_eowfyzlvx7gjv542upo (s_eowfyzlvx7gjv542upo ),

     .d40pep591l63yhmefp7i      (d40pep591l63yhmefp7i      ),

     .t57d026x085pay       (t57d026x085pay       ),
     .k5th293qdrtsytaehbsk      (k5th293qdrtsytaehbsk      ),
     .g6gwjq519o1w1m3csgrrf3  (g6gwjq519o1w1m3csgrrf3  ),
     .lo_2ny7_v71by78q3        (lo_2ny7_v71by78q3        ),
     .hbdj3fcr8qkfkgzq58o1o2ozh(hbdj3fcr8qkfkgzq58o1o2ozh),
     .m_k_n75bb0f_im9fu_      (m_k_n75bb0f_im9fu_      ),

     .jgm2b78on4di5vswgsdt               (e1jv60iid34gonwyukkue                  ),           
     .tuui0ewt7j2chov1tdfd              (xz57o2ko5gkcbk8rq                 ),          
     .u_g5yts7tlcxo7ykedbqiv4ji0             (grv8y38uxakr22asia                ),         
     .qdiqiuzopx36bi3s6fbh7mc16h2cj0         (bvmb0d5jendar95w7nbnob8            ),           
     .urdbh4qug0s4u_dxqek3ejkxxgejj          (h47i__o10wyo2sbyt58zq1_h5             ),      

     .dep51yq                           (vxwhhz9_cff6uy0x                     ),
     .wk9s3wmc2q0yaa13                   (moj77icm1kmex0900                    ),                
     .s7re1eyp36bjvie                    (hib0x0rvcjwnn75a                     ),                 
     .a1pnq3ko2aaldi7h3xwme             (cgmsm8wvxc5kg90xwvwq0cga              ),                 
     .oq4nxgat71_rnebbasjmv9             (w9mx37ezcezieq_9__94o              ),          
     .rj1ewmv16hujp9xlnpm6a3hhu9y8ml        (hsnr3xtposirc7pmphtiko3xlz         ),     
     .ryfblq1f8us1a8u3gy2gijl12x085ja      (k1jkhgd9bvypwrti7ietjp0n7_nyzu       ),   
     .j6q7tn13h_mjup45od1mu              (qirelbyt49gkn46_f24yxtc               ),           
     .x81uu_gb6esoi095hudjgylqn            (jq4wiwydrozelhpru9snvs0             ),         
     .ql2if76ihe_ppb4rp3buw7            (j6muxslh7pud3298q9d8lc2             ),         

     .ldqpjrsj9dp8yg3uc    (ldqpjrsj9dp8yg3uc  ),
     .s70e4xdis3p67ndpn6fbx    (s70e4xdis3p67ndpn6fbx  ),
     .h9zlka3j3ih8ihpvwvky1  (h9zlka3j3ih8ihpvwvky1),
     
     .tf_tmpul8i8qbm_djvtl5f   (tf_tmpul8i8qbm_djvtl5f ),        
     .qtsqtuxyont41a7h7i6  (qtsqtuxyont41a7h7i6),
                                             
     .w0ve66vjdz8lzwws3ic    (w0ve66vjdz8lzwws3ic  ),
     .df775k2ts6dn4528iq_ce5    (df775k2ts6dn4528iq_ce5  ),
     .k3dychuj1pv4vw7cfj01ft8v  (k3dychuj1pv4vw7cfj01ft8v),
     
     .jh4zf96qrsb31j072n   (jh4zf96qrsb31j072n ),        
     .vfvtxk4jkkc3ql7_rqd  (vfvtxk4jkkc3ql7_rqd),
                                            
     .hv6xxz3oswj4wy4j46    (hv6xxz3oswj4wy4j46  ),
     .q6p7kcdd9o7j3e2c886    (q6p7kcdd9o7j3e2c886  ),
     .ee_yaeclihal4dht69liwy6z  (ee_yaeclihal4dht69liwy6z),
     
     .thl4cxcuzntax8hnsn9bl4   (thl4cxcuzntax8hnsn9bl4 ),        
     .mysqpp41yovfcis6f2dza47  (mysqpp41yovfcis6f2dza47),
                                             
     .vp3x08mx4e27x4k26n    (vp3x08mx4e27x4k26n  ),
     .a7b829uahvy2i28yzgg    (a7b829uahvy2i28yzgg  ),
     .kzxrmeg90fb06oya08h1  (kzxrmeg90fb06oya08h1),
     
     .kl5wycr14v5ukl7oqfhwe6   (kl5wycr14v5ukl7oqfhwe6 ),        
     .wt6c82_zmqgmt7if41t698  (wt6c82_zmqgmt7if41t698),

                                            


    .c4ughu0qm5sfai(c4ughu0qm5sfai),

    .gc4b3kdcan6do88ta_  (gc4b3kdcan6do88ta_),






     .wz_if_2q_23jhl2    (wz_if_2q_23jhl2    ),


      .pcr4upio7_tx37     (pcr4upio7_tx37   ), 
      .uzklqlncpqqm1rav  (uzklqlncpqqm1rav),
      .ortueunvnkx_l5m_j  (ortueunvnkx_l5m_j),
      .hwuhtb7ucto_utk56  (hwuhtb7ucto_utk56),
      .i1env2kmns7qvvuuc  (i1env2kmns7qvvuuc),
      .g3s3vpafvy3i  (g3s3vpafvy3i),


     .th06du2c8e2_b7k  (l3fd1x5l3xpi3bbwblpsrwwruvvw),
     .irjoi8wvo25u209f_5  (awh5wdqsak51daa1xam8ipi9),
     .zvk11dhgg2s67mkq   (r_ktqd4uca5y4b3gnhz03iwd ),
     .fbzs0o4ysyuzeg_qdj  (mi8oba8vxuze_93cxrid23bv),
     .me1n4pvwxa7n3u8l05  (kya1iiz3vedj6v1ucdydery90b),
     .qaidts35dk5jcji0n  (mfxhd3_j98125z7zj4spfnef1m6rw),
     .r8nzx6_1no31zeloft  (y0ozra0qgen9l9te2u_pqq0bx4a),


     .phzkntckzzbndu4wevf1o6  (wv8wwd_1gm9_e7vubue9gb29),
     .bpyef3a0dnkkyqdpymy    (yijhfr84p7xs3yctj1skm24t02_  ),
     .wv442dsr_nxty0qoldk7qmqg (jz08e92smloz0op1zfo3g9ungcnbc),   
     .b2loifdzo9b2smec06r0t (crrw2ei1pk6riohtoykjv9qeuen),   
     .tx07brh7_ullbwlubonaqwg2(ttqo192f6935w8y576tjxiwa30fd),   
     .ba1ucnyekcm68i9wuqwmn  (e45yjvds31b0kqjvsynzmgpf),


     .rinamilgle00i5xmx_vt (x27lqkgq55knwoqsc6_bn0p), 
     .j8wlfupbw25hdmohz5q0 (ud5ygg9b8pmm93drtbfk4l8hv),
     .z64bwdr23steb7s9y9j  (f_lrqmtz5mpqmbrhn6f05 ),
     .bg1spy6_v2kbo75pz1d6  (ss92bd8t5gyfjfl1_lp2 ),
     .b7aet1zp_fcfxn8h7rw0u1 (z1beclu7k0_h4nn6njz05sbe1),
     .t3szwnvfo2nj3wk6r5kvt  (w1i6s2iwu2nnj7idywd),
     .cneu8a119tg3vmie6zr2h_ (czjipv9hqkdx4jllt3ajsl),
     .jw2dzv9gi7gygudyqql6fz (j92g3e8ublsg2d9sjj_i3),
     .o_7kpry6inkqpqi1bf1nd (af3a5ot65per6f87crwmj),
     .ybcilssdlw64sqj1jf2uuk (bjucsszqg5d1sc5etnwvf1),
     .znotwr53pu47f5m1agm    (t37flu99i5ex1j3e_8   ),
     .bngbyv57e7juc0vkk2y8i  (wvjkzp74fi8ed7nnr7xlm3gt   ),

     .ze2bfnigu62i9937pcxnjc (phzkntckzzbndu4wevf1o6), 
     .dm5b92mx0redfbuhs1u3d   (bpyef3a0dnkkyqdpymy),
     .c3vtv1izxu7rm5646jsmmke (ba1ucnyekcm68i9wuqwmn),


    .gf33atgy           (n1wslu68m9v    ),
    .ru_wi         (ru_wi        ) 
  );




  assign h8xul8_er09on = (~tw5xnp59d8x);



endmodule






















module hpwm3nya3 #(
   parameter xio4kx7ep1ojwa_r      = 79,
   parameter cmnocc9r2aiw8za       = 8,
   parameter xholqktr732apzsv8d0  = 3
) (
    input                                    mv5to8v6,                       
    
    input                                    k3n1uuckanw669a,               
    input  [27-1:0]      qfy7pr76nvqld1f,               
    input  [1:0]                             nowfs1y75z9hmhv6r0ppp6vjly,        
    
    output                                   f_8ecse5wf0jrndlozy2070bja,        
    
    output  [20-1:0]        c_lxwlogrc590ejlmhjdrmfmj,          
    
    
    output                                   ugixcggahb26m1glzpuqvpq,         
    output                                   vbpz6tidsg3o93kih6nmamlyg9wmr1zz,   
    output                                   j2dtuvq0m4iir947lery9tpxqwhjj2g3, 
    output                                   wo834bx1b9sidvkaqiq_b7jk,        
    output                                   faamp7iz46_jj1ci8a,             
    
    
    
    
    output                                   v66ux9ovjkzt3jn,                
    output  [27-1:0]     cd3lo77nievm4v3,                 
    output  [1:0]                            rgnht1zljy67subvhyua_,          
    
    input                                    nmlix317bu48vgct7x02m7vgn,          
    input                                    s6zb15tq6xjiqgce5nwjcg7be4,     
    input                                    ry0rypry86op3l_hqbwk8pe32ena3e,   
    input  [xio4kx7ep1ojwa_r-1:0]              h4zmq2srkdf5iaeagd8d7i87,           
    input                                    dzo70vq3_1_kyxyiurxy1d20ed,         
    input                                    b0c0o6unssb9h3tgqck870,         

    output                                   c2_546oy8pb0vifo,                 

    
    input                                    gf33atgy,
    input                                    ru_wi,
    input                                    gc4b3kdcan6do88ta_
);

    localparam pse_9oeblmiqo   = 0;
    
    
    localparam skhfe86rjzr       = 1;
    
    
    localparam c6bt4uxhjt76ybdb  = 2;
    localparam ir1y97hv4a9oct4l  = 3;
    
    localparam pvu039o1s9t1m9x_  = xio4kx7ep1ojwa_r-1;
    localparam obu455a2wnp4vu0  = pvu039o1s9t1m9x_+1-27;
    localparam snj9jgmwt45902 = obu455a2wnp4vu0-1;
    localparam la40sjjy7dga49 = snj9jgmwt45902+1-20;

    localparam rqzr_eaa     = 2'b00;
    localparam eri_rah_b     = 2'b01;
    localparam ib1cruu      = 2'b10;

    localparam b1lh2fnh92    = 2;

    localparam cpuuvz0x4_r5s = cmnocc9r2aiw8za-1;    




    genvar i;
    wire [cmnocc9r2aiw8za-1:0]                  i25ll1dii3u_d2n76;




    wire pj9rc44fi;
    wire vkm_fyjfzj9 = mv5to8v6 | b0c0o6unssb9h3tgqck870;
  ux607_clkgate u_oq26k57nedglq(
    .clk_in        (gf33atgy                   ),
    .clkgate_bypass(gc4b3kdcan6do88ta_        ),
    .clock_en      (vkm_fyjfzj9                ),
    .clk_out       (pj9rc44fi               )
  );




    wire [cmnocc9r2aiw8za-1:0]                 hw9pzy7xw26mqd67;
    
    
    wire [cmnocc9r2aiw8za-1:0]                 pjisxg4auax56ugw;
    
    
    wire [1:0]                               wpxfw0jit8znrgcnnkq3he [cmnocc9r2aiw8za-1:0];
    wire [27-1:0]        ipk9h7z3cggz0wdxsb6yj_3p [cmnocc9r2aiw8za-1:0];
    wire [20-1:0]           bzfogmie89cgtvfq27e3aswmuil9 [cmnocc9r2aiw8za-1:0];
    wire [cmnocc9r2aiw8za-1:0]                 wskyn9jef_ao7fnlha;
    wire [cmnocc9r2aiw8za-1:0]                 yo5yfpeiuk3zechv7ry;
    wire [cmnocc9r2aiw8za-1:0]                 a_jrytlfkm3zom4pys8;
    
    wire [20-1:0]           ufhrnwb_tir83f [cmnocc9r2aiw8za-1:0];
    wire [27-1:0]        da5jkvbuwnfukf5p [cmnocc9r2aiw8za-1:0];

    wire [cmnocc9r2aiw8za-1:0]                 dqb744wwgwrkj8pmzlqz;
    
    

    
    
    reg                                      cpznd0fzt2newpz7w_;
    
    
    
    reg [20-1:0]            rtdki0i0xl5hvqfbkj371;


    wire [cmnocc9r2aiw8za-1:0]                 sgncc5i359h6_b7y9;
    wire [xio4kx7ep1ojwa_r-1:0]                unj96xqpx4osi2 [cmnocc9r2aiw8za-1:0];
    wire [xio4kx7ep1ojwa_r-1:0]                vsbxpc1qp3j8l [cmnocc9r2aiw8za-1:0];
    wire udqn4evfqnp;
    wire eqb83t6;
    wire ku0a1r2r_h4;


generate 
    for(i=0; i<cmnocc9r2aiw8za; i=i+1) begin: n5jg7z9942w5zidr6
        assign hw9pzy7xw26mqd67[i] = vsbxpc1qp3j8l[i][pse_9oeblmiqo];
        
        
        assign pjisxg4auax56ugw[i] = vsbxpc1qp3j8l[i][skhfe86rjzr];
        
        
        assign wpxfw0jit8znrgcnnkq3he[i] = vsbxpc1qp3j8l[i][ir1y97hv4a9oct4l:c6bt4uxhjt76ybdb];
        assign wskyn9jef_ao7fnlha[i] = wpxfw0jit8znrgcnnkq3he[i] == 2'b00;
        assign yo5yfpeiuk3zechv7ry[i] = wpxfw0jit8znrgcnnkq3he[i] == 2'b01;
        assign a_jrytlfkm3zom4pys8[i] = wpxfw0jit8znrgcnnkq3he[i] == 2'b10;
        assign ipk9h7z3cggz0wdxsb6yj_3p[i] = wskyn9jef_ao7fnlha[i] ? {27{1'b1}} : 
                                         yo5yfpeiuk3zechv7ry[i] ? {{27-9{1'b1}}, 9'b0} : 
                                         {{27-18{1'b1}}, 18'b0};
        assign bzfogmie89cgtvfq27e3aswmuil9[i] = wskyn9jef_ao7fnlha[i] ? {20{1'b1}} : 
                                            yo5yfpeiuk3zechv7ry[i] ? {{20-9{1'b1}}, 9'b0} : 
                                            {{20-18{1'b1}}, 18'b0};
        
        assign ufhrnwb_tir83f[i] = vsbxpc1qp3j8l[i][snj9jgmwt45902:la40sjjy7dga49];
        assign da5jkvbuwnfukf5p[i] = vsbxpc1qp3j8l[i][pvu039o1s9t1m9x_:obu455a2wnp4vu0];
        assign dqb744wwgwrkj8pmzlqz[i] = ((qfy7pr76nvqld1f & ipk9h7z3cggz0wdxsb6yj_3p[i]) == (da5jkvbuwnfukf5p[i] & ipk9h7z3cggz0wdxsb6yj_3p[i])) & hw9pzy7xw26mqd67[i];
        
    end
endgenerate

    assign ku0a1r2r_h4 = (|dqb744wwgwrkj8pmzlqz) | mv5to8v6;
    assign eqb83t6 = ku0a1r2r_h4 & k3n1uuckanw669a;
    assign udqn4evfqnp = ~ku0a1r2r_h4 & k3n1uuckanw669a;

    wire [20-1:0]           tup8n0fn9pth5itu3f_au;

    assign tup8n0fn9pth5itu3f_au = {{20-18{1'b0}}, qfy7pr76nvqld1f[17:0]};

    integer j;
    always @(*) begin: vsxvdv5in4v_1f267wqv_2v
        
        
        
        cpznd0fzt2newpz7w_ = 1'b0;
        
        
        
        rtdki0i0xl5hvqfbkj371 = 20'b0;

        for (j=0; j<cmnocc9r2aiw8za; j=j+1) begin: wio55hb7s7eikmtdkw6
            
            
            
            cpznd0fzt2newpz7w_ = cpznd0fzt2newpz7w_ | (pjisxg4auax56ugw[j] & dqb744wwgwrkj8pmzlqz[j]);
            
            
            
            rtdki0i0xl5hvqfbkj371 = rtdki0i0xl5hvqfbkj371 | (((ufhrnwb_tir83f[j] & bzfogmie89cgtvfq27e3aswmuil9[j]) | (tup8n0fn9pth5itu3f_au & ~bzfogmie89cgtvfq27e3aswmuil9[j])) & {20{dqb744wwgwrkj8pmzlqz[j]}}); 
        end
    end


    wire                                     twm0b4dd7ahh8f = dzo70vq3_1_kyxyiurxy1d20ed & ~wo834bx1b9sidvkaqiq_b7jk;
    wire                                     pubj1y308jtf6 =  1'b0 
                                                             | (nmlix317bu48vgct7x02m7vgn  & s6zb15tq6xjiqgce5nwjcg7be4)
                                                             | (nmlix317bu48vgct7x02m7vgn  & ry0rypry86op3l_hqbwk8pe32ena3e); 
    wire                                     h624jgnv03hp4iysjt03z = eqb83t6 | twm0b4dd7ahh8f;

    
    wire [cmnocc9r2aiw8za-1:0]                 cs4v4br38e3kc1mou;
    wire [cmnocc9r2aiw8za-1:0]                 jsb3cun4k6fukeall7w71;
    wire                                     prkeaifroj4g2dpakqjw;
    wire [cmnocc9r2aiw8za-1:0]                 kvpghm6ix33yptbkacv4v8xgof;

    assign prkeaifroj4g2dpakqjw = h624jgnv03hp4iysjt03z;
    assign jsb3cun4k6fukeall7w71 = eqb83t6 ? dqb744wwgwrkj8pmzlqz : kvpghm6ix33yptbkacv4v8xgof;
    ux607_gnrl_dfflr #(cmnocc9r2aiw8za) i_cj4uews4woe6jhe8zk4h (prkeaifroj4g2dpakqjw, jsb3cun4k6fukeall7w71, cs4v4br38e3kc1mou, gf33atgy, ru_wi);

    
    wire                                     pukahq7l38_zm0c_t;
    wire                                     mke2bj8i42idruey0et0;
    wire                                     a9_ke8p4rgkl0e_;

    assign a9_ke8p4rgkl0e_ = h624jgnv03hp4iysjt03z;
    assign mke2bj8i42idruey0et0 = eqb83t6 ? 1'b1 : h4zmq2srkdf5iaeagd8d7i87[pse_9oeblmiqo] & twm0b4dd7ahh8f;
    ux607_gnrl_dfflr #(1) xk5zybrc9dvh6c9vna_0j (a9_ke8p4rgkl0e_, mke2bj8i42idruey0et0, pukahq7l38_zm0c_t, gf33atgy, ru_wi);

    
    
    
    

    
    
    

    
    
    
    

    
    
    

    
    wire                                     zjwl1qdz34pwx9l;
    wire                                     zh3m_2uvc6wm91jm9;
    wire                                     wessf0r1ohspioxg;

    assign wessf0r1ohspioxg = h624jgnv03hp4iysjt03z;
    assign zh3m_2uvc6wm91jm9 = eqb83t6 ? cpznd0fzt2newpz7w_ : h4zmq2srkdf5iaeagd8d7i87[skhfe86rjzr];
    ux607_gnrl_dfflr #(1) q4alfwn_r3zsamq34_tnu (wessf0r1ohspioxg, zh3m_2uvc6wm91jm9, zjwl1qdz34pwx9l, gf33atgy, ru_wi);

    
    
    
    

    
    
    

    
    
    
    

    
    
    

    
    
    
    

    
    
    

    
    wire [20-1:0]           p5gbqclsvfry9on1w1v0;
    wire [20-1:0]           lhmal8igxxt9iviaydtu;
    wire                                     j57nla9hf28_ar8ek7apg;
    wire [20-1:0]           i4bgot3pzg0n4juoif;
    wire [1:0]                               io6sh2oqx3bsah15unjfp2l_97b;
    wire                                     ujykf7uo0adtw5zvngkq8t1i;
    wire                                     bxmci6y3rhm4tcn1t6cxjv;
    wire [20-1:0]           pn91hcl3rg1c11q9t5ccdlcbkq6dp;
    wire [20-1:0]           u5k65gvbjzxn790cd7fsnipre9zf;

    
    assign i4bgot3pzg0n4juoif        = {{20-18{1'b0}}, cd3lo77nievm4v3[17:0]};
    assign io6sh2oqx3bsah15unjfp2l_97b = h4zmq2srkdf5iaeagd8d7i87[ir1y97hv4a9oct4l:c6bt4uxhjt76ybdb];
    assign ujykf7uo0adtw5zvngkq8t1i = (io6sh2oqx3bsah15unjfp2l_97b == 2'b00);
    assign bxmci6y3rhm4tcn1t6cxjv = (io6sh2oqx3bsah15unjfp2l_97b == 2'b01);
    assign pn91hcl3rg1c11q9t5ccdlcbkq6dp = ujykf7uo0adtw5zvngkq8t1i ? {20{1'b1}} :
                                      bxmci6y3rhm4tcn1t6cxjv ? {{20-9{1'b1}}, 9'b0} :
                                      {{20-18{1'b1}}, 18'b0};
    assign u5k65gvbjzxn790cd7fsnipre9zf = (pn91hcl3rg1c11q9t5ccdlcbkq6dp & h4zmq2srkdf5iaeagd8d7i87[snj9jgmwt45902:la40sjjy7dga49]) | (~pn91hcl3rg1c11q9t5ccdlcbkq6dp & i4bgot3pzg0n4juoif);

    assign j57nla9hf28_ar8ek7apg = h624jgnv03hp4iysjt03z;
    assign lhmal8igxxt9iviaydtu = eqb83t6 ? rtdki0i0xl5hvqfbkj371 : u5k65gvbjzxn790cd7fsnipre9zf;
    ux607_gnrl_dfflr #(20) x8azcwrk7rdz0suqs8j9_ (j57nla9hf28_ar8ek7apg, lhmal8igxxt9iviaydtu, p5gbqclsvfry9on1w1v0, gf33atgy, ru_wi);

    
    wire [27-1:0]        bue4c0f7wem;
    wire [27-1:0]        c8g3mt3pg2jlm;
    wire                                     ltew2bxq6eu9aq;

    assign ltew2bxq6eu9aq = udqn4evfqnp;   
    assign c8g3mt3pg2jlm = qfy7pr76nvqld1f;
    ux607_gnrl_dfflr #(27) e05s_wh1wka33p0z1 (ltew2bxq6eu9aq, c8g3mt3pg2jlm, bue4c0f7wem, gf33atgy, ru_wi);

    
    wire [1:0]                               zw6ebpxucv29fhmsar7lgm;
    wire [1:0]                               geg04wqhw3xlb8kdlk4fsut1lp;
    wire                                     r8uj6dter_go27zb47a_th3048v0s;

    assign r8uj6dter_go27zb47a_th3048v0s = udqn4evfqnp;   
    assign geg04wqhw3xlb8kdlk4fsut1lp = nowfs1y75z9hmhv6r0ppp6vjly;
    ux607_gnrl_dfflr #(2) qe94e6sl1210uw3gnz6eiycgn8 (r8uj6dter_go27zb47a_th3048v0s, geg04wqhw3xlb8kdlk4fsut1lp, zw6ebpxucv29fhmsar7lgm, gf33atgy, ru_wi);




generate 
    for(i=0; i<cmnocc9r2aiw8za; i=i+1) begin: mpi9jkoirzo4ev3ab
        assign sgncc5i359h6_b7y9[i] = mv5to8v6 | (twm0b4dd7ahh8f & kvpghm6ix33yptbkacv4v8xgof[i]);
        assign unj96xqpx4osi2[i] = mv5to8v6 ? {xio4kx7ep1ojwa_r{1'b0}} : h4zmq2srkdf5iaeagd8d7i87;

        ux607_gnrl_dfflr #(1) mg4hio46oqao1_ij4 (sgncc5i359h6_b7y9[i], unj96xqpx4osi2[i][0], vsbxpc1qp3j8l[i][0], pj9rc44fi, ru_wi);
        ux607_gnrl_dfflr #(xio4kx7ep1ojwa_r-1) koqjnfv662ks1 (sgncc5i359h6_b7y9[i], unj96xqpx4osi2[i][xio4kx7ep1ojwa_r-1:1], vsbxpc1qp3j8l[i][xio4kx7ep1ojwa_r-1:1], pj9rc44fi, ru_wi);
    end
endgenerate




wire [cpuuvz0x4_r5s-1:0] blk93p1i16xx;
wire xtuu_xtcsg4icbv_ = &hw9pzy7xw26mqd67; 
wire [cpuuvz0x4_r5s-1:0] vs7xk5fv2idvsx3b;
wire [cmnocc9r2aiw8za-1:0] j6u1lgj0jf7udo;
wire [cmnocc9r2aiw8za-1:0] bnrmlmaiin9wudfye9v7j7; 

generate
if(cmnocc9r2aiw8za ==16) begin:vt5kaq6
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
    assign bnrmlmaiin9wudfye9v7j7 =  dqb744wwgwrkj8pmzlqz;

    assign i25ll1dii3u_d2n76[0]  = ~blk93p1i16xx[7]  &  ~blk93p1i16xx[3] & ~blk93p1i16xx[1] &  ~blk93p1i16xx[0] & xtuu_xtcsg4icbv_;
    assign i25ll1dii3u_d2n76[1]  =  blk93p1i16xx[7]  &  ~blk93p1i16xx[3] & ~blk93p1i16xx[1] &  ~blk93p1i16xx[0] & xtuu_xtcsg4icbv_;
    assign i25ll1dii3u_d2n76[2]  = ~blk93p1i16xx[8]  &   blk93p1i16xx[3] & ~blk93p1i16xx[1] &  ~blk93p1i16xx[0] & xtuu_xtcsg4icbv_;
    assign i25ll1dii3u_d2n76[3]  =  blk93p1i16xx[8]  &   blk93p1i16xx[3] & ~blk93p1i16xx[1] &  ~blk93p1i16xx[0] & xtuu_xtcsg4icbv_;
    assign i25ll1dii3u_d2n76[4]  = ~blk93p1i16xx[9]  &  ~blk93p1i16xx[4] &  blk93p1i16xx[1] &  ~blk93p1i16xx[0] & xtuu_xtcsg4icbv_;
    assign i25ll1dii3u_d2n76[5]  =  blk93p1i16xx[9]  &  ~blk93p1i16xx[4] &  blk93p1i16xx[1] &  ~blk93p1i16xx[0] & xtuu_xtcsg4icbv_;
    assign i25ll1dii3u_d2n76[6]  = ~blk93p1i16xx[10] &   blk93p1i16xx[4] &  blk93p1i16xx[1] &  ~blk93p1i16xx[0] & xtuu_xtcsg4icbv_;
    assign i25ll1dii3u_d2n76[7]  =  blk93p1i16xx[10] &   blk93p1i16xx[4] &  blk93p1i16xx[1] &  ~blk93p1i16xx[0] & xtuu_xtcsg4icbv_;
    assign i25ll1dii3u_d2n76[8]  = ~blk93p1i16xx[11] &  ~blk93p1i16xx[5] & ~blk93p1i16xx[2] &   blk93p1i16xx[0] & xtuu_xtcsg4icbv_;
    assign i25ll1dii3u_d2n76[9]  =  blk93p1i16xx[11] &  ~blk93p1i16xx[5] & ~blk93p1i16xx[2] &   blk93p1i16xx[0] & xtuu_xtcsg4icbv_;
    assign i25ll1dii3u_d2n76[10] = ~blk93p1i16xx[12] &   blk93p1i16xx[5] & ~blk93p1i16xx[2] &   blk93p1i16xx[0] & xtuu_xtcsg4icbv_;
    assign i25ll1dii3u_d2n76[11] =  blk93p1i16xx[12] &   blk93p1i16xx[5] & ~blk93p1i16xx[2] &   blk93p1i16xx[0] & xtuu_xtcsg4icbv_;
    assign i25ll1dii3u_d2n76[12] = ~blk93p1i16xx[13] &  ~blk93p1i16xx[6] &  blk93p1i16xx[2] &   blk93p1i16xx[0] & xtuu_xtcsg4icbv_;
    assign i25ll1dii3u_d2n76[13] =  blk93p1i16xx[13] &  ~blk93p1i16xx[6] &  blk93p1i16xx[2] &   blk93p1i16xx[0] & xtuu_xtcsg4icbv_;
    assign i25ll1dii3u_d2n76[14] = ~blk93p1i16xx[14] &   blk93p1i16xx[6] &  blk93p1i16xx[2] &   blk93p1i16xx[0] & xtuu_xtcsg4icbv_;
    assign i25ll1dii3u_d2n76[15] =  blk93p1i16xx[14] &   blk93p1i16xx[6] &  blk93p1i16xx[2] &   blk93p1i16xx[0] & xtuu_xtcsg4icbv_;

    assign vs7xk5fv2idvsx3b = ({15{j6u1lgj0jf7udo[0]}} & {blk93p1i16xx[14:8],1'b1,blk93p1i16xx[6:4],1'b1,blk93p1i16xx[2], 2'b11}) |
                             ({15{j6u1lgj0jf7udo[1]}} & {blk93p1i16xx[14:8],1'b0,blk93p1i16xx[6:4],1'b1,blk93p1i16xx[2], 2'b11}) |
                             ({15{j6u1lgj0jf7udo[2]}} & {blk93p1i16xx[14:9],1'b1,blk93p1i16xx[7:4],1'b0,blk93p1i16xx[2], 2'b11}) |
                             ({15{j6u1lgj0jf7udo[3]}} & {blk93p1i16xx[14:9],1'b0,blk93p1i16xx[7:4],1'b0,blk93p1i16xx[2], 2'b11}) |
                             ({15{j6u1lgj0jf7udo[4]}} & {blk93p1i16xx[14:10],1'b1,blk93p1i16xx[8:5],1'b1,blk93p1i16xx[3:2], 2'b01}) |
                             ({15{j6u1lgj0jf7udo[5]}} & {blk93p1i16xx[14:10],1'b0,blk93p1i16xx[8:5],1'b1,blk93p1i16xx[3:2], 2'b01}) |
                             ({15{j6u1lgj0jf7udo[6]}} & {blk93p1i16xx[14:11],1'b1,blk93p1i16xx[9:5],1'b0,blk93p1i16xx[3:2], 2'b01}) |
                             ({15{j6u1lgj0jf7udo[7]}} & {blk93p1i16xx[14:11],1'b0,blk93p1i16xx[9:5],1'b0,blk93p1i16xx[3:2], 2'b01}) |
                             ({15{j6u1lgj0jf7udo[8]}} & {blk93p1i16xx[14:12],1'b1,blk93p1i16xx[10:6],1'b1,blk93p1i16xx[4:3],  1'b1,blk93p1i16xx[1],1'b0}) |
                             ({15{j6u1lgj0jf7udo[9]}} & {blk93p1i16xx[14:12],1'b0,blk93p1i16xx[10:6],1'b1,blk93p1i16xx[4:3],  1'b1,blk93p1i16xx[1],1'b0}) |
                             ({15{j6u1lgj0jf7udo[10]}} & {blk93p1i16xx[14:13],1'b1,blk93p1i16xx[11:6],1'b0,blk93p1i16xx[4:3], 1'b1,blk93p1i16xx[1],1'b0}) |
                             ({15{j6u1lgj0jf7udo[11]}} & {blk93p1i16xx[14:13],1'b0,blk93p1i16xx[11:6],1'b0,blk93p1i16xx[4:3], 1'b1,blk93p1i16xx[1],1'b0}) |
                             ({15{j6u1lgj0jf7udo[12]}} & {blk93p1i16xx[14],1'b1,blk93p1i16xx[12:7],1'b1,blk93p1i16xx[5:3],  1'b0,blk93p1i16xx[1],1'b0}) |
                             ({15{j6u1lgj0jf7udo[13]}} & {blk93p1i16xx[14],1'b0,blk93p1i16xx[12:7],1'b1,blk93p1i16xx[5:3],  1'b0,blk93p1i16xx[1],1'b0}) |
                             ({15{j6u1lgj0jf7udo[14]}} & {1'b1,blk93p1i16xx[13:7],1'b0,blk93p1i16xx[5:3], 1'b0,blk93p1i16xx[1],1'b0}) |
                             ({15{j6u1lgj0jf7udo[15]}} & {1'b0,blk93p1i16xx[13:7],1'b0,blk93p1i16xx[5:3], 1'b0,blk93p1i16xx[1],1'b0});
end
else if(cmnocc9r2aiw8za ==8) begin:g62rpi2e
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
    assign bnrmlmaiin9wudfye9v7j7 =  dqb744wwgwrkj8pmzlqz;

    assign i25ll1dii3u_d2n76[0]  = ~blk93p1i16xx[3] & ~blk93p1i16xx[1] &  ~blk93p1i16xx[0] & xtuu_xtcsg4icbv_;
    assign i25ll1dii3u_d2n76[1]  =  blk93p1i16xx[3] & ~blk93p1i16xx[1] &  ~blk93p1i16xx[0] & xtuu_xtcsg4icbv_;
    assign i25ll1dii3u_d2n76[2]  = ~blk93p1i16xx[4] &  blk93p1i16xx[1] &  ~blk93p1i16xx[0] & xtuu_xtcsg4icbv_;
    assign i25ll1dii3u_d2n76[3]  =  blk93p1i16xx[4] &  blk93p1i16xx[1] &  ~blk93p1i16xx[0] & xtuu_xtcsg4icbv_;
    assign i25ll1dii3u_d2n76[4]  = ~blk93p1i16xx[5] & ~blk93p1i16xx[2] &   blk93p1i16xx[0] & xtuu_xtcsg4icbv_;
    assign i25ll1dii3u_d2n76[5]  =  blk93p1i16xx[5] & ~blk93p1i16xx[2] &   blk93p1i16xx[0] & xtuu_xtcsg4icbv_;
    assign i25ll1dii3u_d2n76[6]  = ~blk93p1i16xx[6] &  blk93p1i16xx[2] &   blk93p1i16xx[0] & xtuu_xtcsg4icbv_;
    assign i25ll1dii3u_d2n76[7]  =  blk93p1i16xx[6] &  blk93p1i16xx[2] &   blk93p1i16xx[0] & xtuu_xtcsg4icbv_;

                          

    assign vs7xk5fv2idvsx3b = ({7{j6u1lgj0jf7udo[0]}} & {blk93p1i16xx[6:4],1'b1,blk93p1i16xx[2],2'b11})
                           | ({7{j6u1lgj0jf7udo[1]}} & {blk93p1i16xx[6:4],1'b0,blk93p1i16xx[2],2'b11})
                           | ({7{j6u1lgj0jf7udo[2]}} & {blk93p1i16xx[6:5],1'b1,blk93p1i16xx[3:2],2'b01})
                           | ({7{j6u1lgj0jf7udo[3]}} & {blk93p1i16xx[6:5],1'b0,blk93p1i16xx[3:2],2'b01})
                           | ({7{j6u1lgj0jf7udo[4]}} & {blk93p1i16xx[6],1'b1,blk93p1i16xx[4:3],1'b1,blk93p1i16xx[1],1'b0})
                           | ({7{j6u1lgj0jf7udo[5]}} & {blk93p1i16xx[6],1'b0,blk93p1i16xx[4:3],1'b1,blk93p1i16xx[1],1'b0})
                           | ({7{j6u1lgj0jf7udo[6]}} & {1'b1,blk93p1i16xx[5:3],1'b0,blk93p1i16xx[1],1'b0})
                           | ({7{j6u1lgj0jf7udo[7]}} & {1'b0,blk93p1i16xx[5:3],1'b0,blk93p1i16xx[1],1'b0})
                           ;
end
else begin:g4j8p5
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
    assign bnrmlmaiin9wudfye9v7j7 =  dqb744wwgwrkj8pmzlqz;

    assign i25ll1dii3u_d2n76[0]  =  ~blk93p1i16xx[1] &  ~blk93p1i16xx[0] & xtuu_xtcsg4icbv_;
    assign i25ll1dii3u_d2n76[1]  =   blk93p1i16xx[1] &  ~blk93p1i16xx[0] & xtuu_xtcsg4icbv_;
    assign i25ll1dii3u_d2n76[2]  =  ~blk93p1i16xx[2] &   blk93p1i16xx[0] & xtuu_xtcsg4icbv_;
    assign i25ll1dii3u_d2n76[3]  =   blk93p1i16xx[2] &   blk93p1i16xx[0] & xtuu_xtcsg4icbv_;

                          

    assign vs7xk5fv2idvsx3b = ({3{j6u1lgj0jf7udo[0]}} & {blk93p1i16xx[2],2'b11})
                           | ({3{j6u1lgj0jf7udo[1]}} & {blk93p1i16xx[2],2'b01})
                           | ({3{j6u1lgj0jf7udo[2]}} & {1'b1,blk93p1i16xx[1],1'b0})
                           | ({3{j6u1lgj0jf7udo[3]}} & {1'b0,blk93p1i16xx[1],1'b0})
                           ;
end
endgenerate

assign j6u1lgj0jf7udo = mv5to8v6 ? {cmnocc9r2aiw8za{1'b0}} : eqb83t6 ? bnrmlmaiin9wudfye9v7j7 : i25ll1dii3u_d2n76;

wire ou029l35_79b7g0uc00638i = (xtuu_xtcsg4icbv_ & (eqb83t6 | twm0b4dd7ahh8f)) | mv5to8v6;
ux607_gnrl_dfflr #(cpuuvz0x4_r5s) paca0uqimbbvs4d0n933f(ou029l35_79b7g0uc00638i,vs7xk5fv2idvsx3b,blk93p1i16xx,gf33atgy,ru_wi); 

wire [cmnocc9r2aiw8za-1:0] dc3tx2ejpweplpq8ck1f27 =  {hw9pzy7xw26mqd67[cmnocc9r2aiw8za-2:0],1'b1} ^ hw9pzy7xw26mqd67;
wire [cmnocc9r2aiw8za-1:0] re7qj5c2go8inyaoucg;

generate
for(i=0;i<cmnocc9r2aiw8za;i=i+1) begin:sxq_amt5geudw_mtdr8g2d41y2
    if(i==0) begin:t9w81cc3ejd_
        assign re7qj5c2go8inyaoucg[i] = dc3tx2ejpweplpq8ck1f27[0];
    end
    else begin:cghdgmfjwlvv
        assign re7qj5c2go8inyaoucg[i] = |dc3tx2ejpweplpq8ck1f27[i:0];
    end
end
endgenerate

wire [cmnocc9r2aiw8za-1:0] ridudot9q3ozuzce_05rf = {re7qj5c2go8inyaoucg[cmnocc9r2aiw8za-2:0],1'b0} ^ re7qj5c2go8inyaoucg;

assign kvpghm6ix33yptbkacv4v8xgof =  (xtuu_xtcsg4icbv_ ? i25ll1dii3u_d2n76 : ridudot9q3ozuzce_05rf);












    wire [b1lh2fnh92-1:0]         sat482scl8zle;
    wire [b1lh2fnh92-1:0]         fdr3d671e7dw6;
    wire                         h8ghyl6u7gffe;
    wire [b1lh2fnh92-1:0]         u99tnldu986760c5;
    wire [b1lh2fnh92-1:0]         y5ramxcxkrqsz12gk;
    wire [b1lh2fnh92-1:0]         frmnwpwxl1k1l;
    wire                         wfoen161d4r42bkqp34lj;
    wire                         hln5byq3t_zxwy8c51dq;
    wire                         klef245vk22hxpmozv2gww9;
    
    wire                         uoozmjtee2uc_8o;
    wire                         ejae6qevtda080dzd5d;
    

    assign c2_546oy8pb0vifo = (sat482scl8zle == rqzr_eaa);
    assign uoozmjtee2uc_8o = (sat482scl8zle == eri_rah_b);
    assign ejae6qevtda080dzd5d  = (sat482scl8zle == ib1cruu);

    
    assign wfoen161d4r42bkqp34lj = c2_546oy8pb0vifo & k3n1uuckanw669a;
    assign u99tnldu986760c5 = udqn4evfqnp ? eri_rah_b : ib1cruu;

    
    assign hln5byq3t_zxwy8c51dq = uoozmjtee2uc_8o & nmlix317bu48vgct7x02m7vgn;
    assign y5ramxcxkrqsz12gk = ib1cruu;

    
    assign klef245vk22hxpmozv2gww9 = ejae6qevtda080dzd5d;
    assign frmnwpwxl1k1l = k3n1uuckanw669a ? (udqn4evfqnp ? eri_rah_b : ib1cruu) : rqzr_eaa;

    

    assign h8ghyl6u7gffe = wfoen161d4r42bkqp34lj | hln5byq3t_zxwy8c51dq | klef245vk22hxpmozv2gww9;
    assign fdr3d671e7dw6 =    ({b1lh2fnh92{wfoen161d4r42bkqp34lj}} & u99tnldu986760c5)
                            | ({b1lh2fnh92{hln5byq3t_zxwy8c51dq}} & y5ramxcxkrqsz12gk)
                            | ({b1lh2fnh92{klef245vk22hxpmozv2gww9 }} & frmnwpwxl1k1l )
                            ; 

    ux607_gnrl_dfflr #(b1lh2fnh92) afp_kqyn5ft8m (h8ghyl6u7gffe, fdr3d671e7dw6, sat482scl8zle, gf33atgy, ru_wi);




    assign v66ux9ovjkzt3jn = uoozmjtee2uc_8o;
    assign cd3lo77nievm4v3  = bue4c0f7wem;
    assign rgnht1zljy67subvhyua_  = zw6ebpxucv29fhmsar7lgm;





    wire               lvn1okew4e1jm302yzyht;                      
    wire               yzpvj2cp44tuel91z9tankq;                      
    wire               jl9t_wr0467jngt74lx01c1i;                      
    wire               cz553_d0qlsc1tvrmb0pkrz5uv;                     
    wire               sxfvetk5l8uqosb5bso;                     

    
    assign lvn1okew4e1jm302yzyht = ejae6qevtda080dzd5d;
    assign yzpvj2cp44tuel91z9tankq =  (s6zb15tq6xjiqgce5nwjcg7be4 & nmlix317bu48vgct7x02m7vgn)
                                  
                                  ;
    assign jl9t_wr0467jngt74lx01c1i = lvn1okew4e1jm302yzyht | yzpvj2cp44tuel91z9tankq;
    assign cz553_d0qlsc1tvrmb0pkrz5uv = (~lvn1okew4e1jm302yzyht) | yzpvj2cp44tuel91z9tankq;
    ux607_gnrl_dfflr #(1) vosya7d_jl9ii7cu (jl9t_wr0467jngt74lx01c1i, cz553_d0qlsc1tvrmb0pkrz5uv, sxfvetk5l8uqosb5bso, gf33atgy, ru_wi);


    wire               aw85z9wxo3a1iwczeohvkpc;                      
    wire               s979qn1uap58cnr3kge2j6pl0;                      
    wire               g838isxs19zm_951h0biuas7dc;                      
    wire               fu89finup50npmbs18hvxyxvv;                     
    wire               omud9qoq5c70_nn_efulbdo3;                     

    
    assign aw85z9wxo3a1iwczeohvkpc = ejae6qevtda080dzd5d;
    assign s979qn1uap58cnr3kge2j6pl0 = ry0rypry86op3l_hqbwk8pe32ena3e & nmlix317bu48vgct7x02m7vgn;
    assign g838isxs19zm_951h0biuas7dc = aw85z9wxo3a1iwczeohvkpc | s979qn1uap58cnr3kge2j6pl0;
    assign fu89finup50npmbs18hvxyxvv = (~aw85z9wxo3a1iwczeohvkpc) | s979qn1uap58cnr3kge2j6pl0;
    ux607_gnrl_dfflr #(1) wg3u77daogjarffm_ise9b (g838isxs19zm_951h0biuas7dc, fu89finup50npmbs18hvxyxvv, omud9qoq5c70_nn_efulbdo3, gf33atgy, ru_wi);




    wire               bdfdk1o4b6647hu3qx82;
    wire               l1tts73djyx9lk4r;
    wire               gu63gtn9gi__3y_9oyq9;
    wire               f4fljw8rmon9pad98riz;
    wire               p0xp_q1lw16gkpbca;
    
    assign bdfdk1o4b6647hu3qx82 = k3n1uuckanw669a & udqn4evfqnp;
    
    assign l1tts73djyx9lk4r = (k3n1uuckanw669a & eqb83t6) | nmlix317bu48vgct7x02m7vgn;
    assign gu63gtn9gi__3y_9oyq9 = bdfdk1o4b6647hu3qx82 | l1tts73djyx9lk4r;
    assign f4fljw8rmon9pad98riz = ~bdfdk1o4b6647hu3qx82 | l1tts73djyx9lk4r;
    ux607_gnrl_dfflr #(1) q3enzpsnyzym2_yoktd (gu63gtn9gi__3y_9oyq9, f4fljw8rmon9pad98riz, p0xp_q1lw16gkpbca, gf33atgy, ru_wi);

    assign f_8ecse5wf0jrndlozy2070bja = p0xp_q1lw16gkpbca;
    assign c_lxwlogrc590ejlmhjdrmfmj   = p5gbqclsvfry9on1w1v0;
    
    
    assign ugixcggahb26m1glzpuqvpq  = zjwl1qdz34pwx9l;






    assign vbpz6tidsg3o93kih6nmamlyg9wmr1zz = sxfvetk5l8uqosb5bso;                             
    assign j2dtuvq0m4iir947lery9tpxqwhjj2g3 = omud9qoq5c70_nn_efulbdo3;

    assign faamp7iz46_jj1ci8a = uoozmjtee2uc_8o;
    wire              j5djvpfvkybh06fizld9;
    wire              a_s7yn5lzc5x3rkfn0;
    wire              rvo8smiyof7vbbmkg;
    wire              ibvvquk0srq6e9x7y;
    wire              p3ds83l6ptt7zw;

    
    assign j5djvpfvkybh06fizld9 = k3n1uuckanw669a;
    
    assign a_s7yn5lzc5x3rkfn0 = ((k3n1uuckanw669a & eqb83t6) | uoozmjtee2uc_8o) & mv5to8v6;
    assign rvo8smiyof7vbbmkg = j5djvpfvkybh06fizld9 | a_s7yn5lzc5x3rkfn0;
    assign ibvvquk0srq6e9x7y = a_s7yn5lzc5x3rkfn0 | (~j5djvpfvkybh06fizld9);
    ux607_gnrl_dfflr #(1) x90eei5lbts5in0rj0c5z0p (rvo8smiyof7vbbmkg, ibvvquk0srq6e9x7y, p3ds83l6ptt7zw, gf33atgy, ru_wi);

    
    assign wo834bx1b9sidvkaqiq_b7jk = p3ds83l6ptt7zw;

endmodule





















module ux607_gnrl_axi2icb # (
  parameter AW = 32,
  parameter DW = 32,
  parameter ID_W = 4,
  parameter USR_W = 4,
  parameter FIFO_OUTS_NUM = 4,
  parameter ALLOW_BURST = 0,
  parameter MW = 4
)(

  output axi_slave_active,


  output                           axi_arready,
  input                            axi_arvalid,
  input [ID_W-1:0]        axi_arid,
  input [AW-1:0]      axi_araddr,
  input [7:0]                      axi_arlen,
  input [2:0]                      axi_arsize,
  input [1:0]                      axi_arburst,
  input                            axi_arlock,
  input [3:0]                      axi_arcache,
  input [2:0]                      axi_arprot,
  input [3:0]                      axi_arqos,
  input [3:0]                      axi_arregion,
  input [USR_W-1:0]          axi_aruser,

  output                           axi_awready,
  input                            axi_awvalid,
  input [ID_W-1:0]        axi_awid,
  input [AW-1:0]      axi_awaddr,
  input [7:0]                      axi_awlen,
  input [2:0]                      axi_awsize,
  input [1:0]                      axi_awburst,
  input                            axi_awlock,
  input [3:0]                      axi_awcache,
  input [2:0]                      axi_awprot,
  input [3:0]                      axi_awqos,
  input [3:0]                      axi_awregion,
  input [USR_W-1:0]          axi_awuser, 

  output                           axi_wready,
  input                            axi_wvalid,
  input [ID_W-1:0]        axi_wid,
  input [DW-1:0]           axi_wdata,
  input [MW-1:0]        axi_wstrb,
  input                            axi_wlast,

  input                            axi_rready,
  output                           axi_rvalid,
  output [ID_W-1:0]       axi_rid,
  output [DW-1:0]          axi_rdata,
  output [1:0]                     axi_rresp,
  output                           axi_rlast,

  input                            axi_bready,
  output                           axi_bvalid,
  output [ID_W-1:0]       axi_bid,
  output [1:0]                     axi_bresp,

  input                            axi_bus_clk_en,

  output                         icb_cmd_valid ,
  input                          icb_cmd_ready ,
  output [AW-1:0]                icb_cmd_addr  , 
  output                         icb_cmd_read  , 
  output [3-1:0]                 icb_cmd_burst ,
  output [2-1:0]                 icb_cmd_beat  ,
  output [        DW-1:0]        icb_cmd_wdata ,
  output [        MW-1:0]        icb_cmd_wmask ,
  output                         icb_cmd_lock  ,
  output                         icb_cmd_excl  ,
  output [1:0]                   icb_cmd_size  ,
  output                         icb_cmd_sel   ,
  output [USR_W-1:0]             icb_cmd_user   ,

  input                          icb_rsp_valid ,
  output                         icb_rsp_ready ,
  input                          icb_rsp_err   ,
  input                          icb_rsp_excl_ok,
  input  [        DW-1:0]        icb_rsp_rdata ,

  input  clk,
  input  rst_n
  );




  wire          g4k11xiitgz962r  ;
  wire          nxfnmkeh2_oxuinwhs  ;
  wire [AW-1:0] kez7oy1hkm0x_mba   ;
  wire          qozylwb2v0y4igv8   ;
  wire [DW-1:0] d6w6ulxl95ras8b4jl  ;
  wire [MW-1:0] hdfxyj_9lnc9x9ls099  ;
  wire [2:0]    p6apzeecwtoem_e2x87  ;
  wire [1:0]    xmas5gu2txl3r66b1f   ;
  wire          mrpmr1jpfod77q   ;             
  wire [1:0]    om7id6y4jtcq4   ;
  wire [USR_W-1:0]   jq3nag_rg7k24ivb   ;             

  wire          ee0gaim_5o2cowj8cc  ;
  wire          iy0c52aia8jldt99i  ;
  wire [DW-1:0] wtmpbfqxajai_cc  ; 
  wire          dt4m1v705h0fe    ;
  wire          t_xyazag81f8t2zmg8b4;

  wire          hivak1ik74xuevh7l0f_4513   ;             

  ux607_gnrl_axi2icb_read # (
  .AW(AW),
  .DW(DW),
  .MW(MW),
  .BUFFER_DP(2),
  .FIFO_OUTS_NUM(FIFO_OUTS_NUM),
  .ALLOW_BURST (ALLOW_BURST), 
  .ID_W (ID_W),
  .USR_W (USR_W)
  ) laz5u5wq_1914kwviiicc (

    .axi_arready  (axi_arready ),
    .axi_arvalid  (axi_arvalid ),
    .axi_arid     (axi_arid    ),
    .axi_araddr   (axi_araddr  ),
    .axi_arlen    (axi_arlen   ),
    .axi_arsize   (axi_arsize  ),
    .axi_arburst  (axi_arburst ),
    .axi_arlock   (axi_arlock  ),
    .axi_arcache  (axi_arcache ),
    .axi_arprot   (axi_arprot  ),
    .axi_arqos    (axi_arqos   ),
    .axi_arregion (axi_arregion),
    .axi_aruser   (axi_aruser  ),


    .axi_rready   (axi_rready   ),
    .axi_rvalid   (axi_rvalid   ),
    .axi_rid      (axi_rid      ),
    .axi_rdata    (axi_rdata    ),
    .axi_rresp    (axi_rresp    ),
    .axi_rlast    (axi_rlast    ),


    .icb_rcmd_valid (g4k11xiitgz962r ),
    .icb_rcmd_ready (nxfnmkeh2_oxuinwhs ),
    .icb_rcmd_addr  (kez7oy1hkm0x_mba  ),
    .icb_rcmd_read  (qozylwb2v0y4igv8  ),
    .icb_rcmd_wdata (d6w6ulxl95ras8b4jl ),
    .icb_rcmd_wmask (hdfxyj_9lnc9x9ls099 ),
    .icb_rcmd_burst (p6apzeecwtoem_e2x87 ),
    .icb_rcmd_beat  (xmas5gu2txl3r66b1f  ),
    .icb_rcmd_excl  (mrpmr1jpfod77q  ),             
    .icb_rcmd_size  (om7id6y4jtcq4  ),
    .icb_rcmd_usr   (jq3nag_rg7k24ivb  ),

    .icb_rrsp_ready  (ee0gaim_5o2cowj8cc  ), 
    .icb_rrsp_valid  (iy0c52aia8jldt99i  ), 
    .icb_rrsp_rdata  (wtmpbfqxajai_cc  ), 
    .icb_rrsp_err    (dt4m1v705h0fe    ), 
    .icb_rrsp_excl_ok(t_xyazag81f8t2zmg8b4), 

    .axi_bus_clk_en  (axi_bus_clk_en),

    .axi2icb_read_active  (hivak1ik74xuevh7l0f_4513),

    .clk  (clk  ),
    .rst_n(rst_n)  
  );



  wire           v5brbv_o0cwz8ltkbnv ;
  wire           h6vhmpdy12279cq0xb6 ;
  wire [AW-1:0]  zh16cx29t0l33  ;
  wire           kg6c6siv37bjp1  ;
  wire [DW-1:0]  ka4nz5iwhho4_t ;
  wire [MW-1:0]  fzedypimn06pveo8 ;
  wire [2:0]     gsh3nost5unqiaqgo ;
  wire [1:0]     ld9htofs52b7nj  ;
  wire           f22pg5kqjpfmk83h2e  ;             
  wire [1:0]     iwvo07en81_3rvne  ;
  wire [USR_W-1:0]hi_0bv4ttpvt3lv  ;             

  wire           i5ydr9vb80xsvdjv2lm ;
  wire           pimisco33wy7hvy ;
  wire [DW-1:0]  tz3bvqjneeev42ye ; 
  wire           nnqpeie69utf9y5h   ;
  wire           o0d8x1ga2vq5_p_g__k;

  wire           ix0lsijxqslj1lxk0dtiy2fsq;

  ux607_gnrl_axi2icb_write # (
  .AW(AW),
  .DW(DW),
  .MW(MW),
  .BUFFER_DP(2),
  .FIFO_OUTS_NUM(FIFO_OUTS_NUM),
  .ALLOW_BURST (ALLOW_BURST),
  .ID_W (ID_W),
  .USR_W (USR_W)
  ) m216l1l7y9vjvbtp1t44 (

    .axi_awready   (axi_awready   ),
    .axi_awvalid   (axi_awvalid   ),
    .axi_awid      (axi_awid      ),
    .axi_awaddr    (axi_awaddr    ),
    .axi_awlen     (axi_awlen     ),
    .axi_awsize    (axi_awsize    ),
    .axi_awburst   (axi_awburst   ),
    .axi_awlock    (axi_awlock    ),
    .axi_awcache   (axi_awcache   ),
    .axi_awprot    (axi_awprot    ),
    .axi_awqos     (axi_awqos     ),
    .axi_awregion  (axi_awregion  ),
    .axi_awuser    (axi_awuser    ), 

    .axi_wready    (axi_wready    ),
    .axi_wvalid    (axi_wvalid    ),
    .axi_wid       (axi_wid       ),
    .axi_wdata     (axi_wdata     ),
    .axi_wstrb     (axi_wstrb     ),
    .axi_wlast     (axi_wlast     ),

    .axi_bready    (axi_bready    ),
    .axi_bvalid    (axi_bvalid    ),
    .axi_bid       (axi_bid       ),
    .axi_bresp     (axi_bresp     ),

    .icb_wcmd_valid (v5brbv_o0cwz8ltkbnv ),
    .icb_wcmd_ready (h6vhmpdy12279cq0xb6 ),
    .icb_wcmd_addr  (zh16cx29t0l33  ),
    .icb_wcmd_read  (kg6c6siv37bjp1  ), 
    .icb_wcmd_wdata (ka4nz5iwhho4_t ),
    .icb_wcmd_wmask (fzedypimn06pveo8 ),
    .icb_wcmd_burst (gsh3nost5unqiaqgo ),
    .icb_wcmd_beat  (ld9htofs52b7nj  ),
    .icb_wcmd_lock  (               ),
    .icb_wcmd_excl  (f22pg5kqjpfmk83h2e  ),
    .icb_wcmd_size  (iwvo07en81_3rvne  ),
    .icb_wcmd_usr   (hi_0bv4ttpvt3lv ),

    .icb_wrsp_valid  (pimisco33wy7hvy  ),
    .icb_wrsp_ready  (i5ydr9vb80xsvdjv2lm  ),
    .icb_wrsp_err    (nnqpeie69utf9y5h    ),
    .icb_wrsp_excl_ok(o0d8x1ga2vq5_p_g__k),

    .axi_bus_clk_en  (axi_bus_clk_en),

    .axi2icb_write_active  (ix0lsijxqslj1lxk0dtiy2fsq),

    .clk   (clk  ),
    .rst_n (rst_n)
  );





  localparam ubq4gj1kd8vql_2k2 = 2;
  localparam v7uxeap96r379eztgx_ = 1;

  wire [ubq4gj1kd8vql_2k2*1-1:0] k1_j5ubhqqpfrl3p0bi186va9;
  wire [ubq4gj1kd8vql_2k2*1-1:0] w0hjg2xow0ymilw7bcxpm2l;
  wire [ubq4gj1kd8vql_2k2*AW-1:0] xzpsiztjmn62eb967x1xkc6;
  wire [ubq4gj1kd8vql_2k2*1-1:0] a_dm6kd_qbw2cv84wtboltif01;
  wire [ubq4gj1kd8vql_2k2*1-1:0] wspjbjcpf459zy17qhyz8jmqy7;
  wire [ubq4gj1kd8vql_2k2*2-1:0] y7jg1o7n3jl52fxr0isdv8;
  wire [ubq4gj1kd8vql_2k2*DW-1:0] ae00o9ay050qc5d5zxf18282b92;
  wire [ubq4gj1kd8vql_2k2*MW-1:0] puxr8jzij0m30qcwmdz2sufl51;
  wire [ubq4gj1kd8vql_2k2*3-1:0] sxjmcdip1m7ighns0k5aue59fj;
  wire [ubq4gj1kd8vql_2k2*2-1:0] noyjdh392j1x0s9g1b_lk;
  wire [ubq4gj1kd8vql_2k2  -1:0] s6vj39lt1yt7f1ytk3pr3 = {ubq4gj1kd8vql_2k2{1'b0}};
  wire [ubq4gj1kd8vql_2k2*USR_W-1:0] w8o2oxw46tp1zf4rujrx4zyxw ;

  wire [ubq4gj1kd8vql_2k2*1-1:0] qkiytqsa_fo9x5ls7yb_x1k2;
  wire [ubq4gj1kd8vql_2k2*1-1:0] idw2i93am7m9wy_5hzipgymj5k3;
  wire [ubq4gj1kd8vql_2k2*1-1:0] wzmdtyq65i82w_tt0juwqle;
  wire [ubq4gj1kd8vql_2k2*1-1:0] kz10yoaxkacgm38dwv37tl2ixfv;
  wire [ubq4gj1kd8vql_2k2*DW-1:0] fyvkbec2dn4rlcslyiyttfrx;
  wire [ubq4gj1kd8vql_2k2*USR_W-1:0] od5a1yudx9bmyqpwleexh4h9;















  assign k1_j5ubhqqpfrl3p0bi186va9 =
                           {
                             g4k11xiitgz962r,
                             v5brbv_o0cwz8ltkbnv
                           } ;

  wire[ubq4gj1kd8vql_2k2-1:0] ccxw7l8izxzjj14ozqkgvvyd6 =









                           {ubq4gj1kd8vql_2k2{1'b0}};

  assign xzpsiztjmn62eb967x1xkc6 =
                           {
                             kez7oy1hkm0x_mba,
                             zh16cx29t0l33
                           } ;

  assign a_dm6kd_qbw2cv84wtboltif01 =
                           {
                             qozylwb2v0y4igv8,
                             kg6c6siv37bjp1
                           } ;

  assign ae00o9ay050qc5d5zxf18282b92 =
                           {
                             d6w6ulxl95ras8b4jl,
                             ka4nz5iwhho4_t
                           } ;

  assign puxr8jzij0m30qcwmdz2sufl51 =
                           {
                             hdfxyj_9lnc9x9ls099,
                             fzedypimn06pveo8
                           } ;

  assign sxjmcdip1m7ighns0k5aue59fj =
                           {
                             p6apzeecwtoem_e2x87,
                             gsh3nost5unqiaqgo
                           } ;

  assign noyjdh392j1x0s9g1b_lk =
                           {
                             xmas5gu2txl3r66b1f,
                             ld9htofs52b7nj
                           } ;

  assign wspjbjcpf459zy17qhyz8jmqy7 =
                           {
                             mrpmr1jpfod77q,
                             f22pg5kqjpfmk83h2e
                           } ;

  assign y7jg1o7n3jl52fxr0isdv8 =
                           {
                             om7id6y4jtcq4,
                             iwvo07en81_3rvne
                           } ;

  assign w8o2oxw46tp1zf4rujrx4zyxw =
                           {
                             jq3nag_rg7k24ivb,
                             hi_0bv4ttpvt3lv
                           } ;

  assign                   {
                             nxfnmkeh2_oxuinwhs,
                             h6vhmpdy12279cq0xb6
                           } = w0hjg2xow0ymilw7bcxpm2l;


  assign                   {
                             iy0c52aia8jldt99i,
                             pimisco33wy7hvy
                           } = qkiytqsa_fo9x5ls7yb_x1k2;

  assign                   {
                             dt4m1v705h0fe,
                             nnqpeie69utf9y5h
                           } = wzmdtyq65i82w_tt0juwqle;

  assign                   {
                             t_xyazag81f8t2zmg8b4,
                             o0d8x1ga2vq5_p_g__k
                           } = kz10yoaxkacgm38dwv37tl2ixfv;

  assign                   {
                             wtmpbfqxajai_cc,
                             tz3bvqjneeev42ye
                           } = fyvkbec2dn4rlcslyiyttfrx;

  assign idw2i93am7m9wy_5hzipgymj5k3 = {
                             ee0gaim_5o2cowj8cc,
                             i5ydr9vb80xsvdjv2lm
                           };

  wire l0_5x2ohgu6m77k54mg;

  ux607_gnrl_icb_arbt # (

  .ALLOW_BURST (ALLOW_BURST),

  .ARBT_SCHEME (1),
  .FIFO_CUT_READY  (0),
  .ALLOW_0CYCL_RSP (0),

  .FIFO_OUTS_NUM   (FIFO_OUTS_NUM),
  .ARBT_NUM   (ubq4gj1kd8vql_2k2),
  .ARBT_PTR_W (v7uxeap96r379eztgx_),
  .USR_W      (USR_W),
  .AW         (AW),
  .DW         (DW) 
  ) jxbdlhwd92pzn3e(
  .arbt_active            (l0_5x2ohgu6m77k54mg),                      
  .o_icb_cmd_valid        (icb_cmd_valid ),                     
  .o_icb_cmd_ready        (icb_cmd_ready ),                     
  .o_icb_cmd_read         (icb_cmd_read  ),                     
  .o_icb_cmd_addr         (icb_cmd_addr  ),                     
  .o_icb_cmd_wdata        (icb_cmd_wdata ),                     
  .o_icb_cmd_wmask        (icb_cmd_wmask ),                     
  .o_icb_cmd_burst        (icb_cmd_burst ),                     
  .o_icb_cmd_beat         (icb_cmd_beat  ),                     
  .o_icb_cmd_excl         (icb_cmd_excl  ),                     
  .o_icb_cmd_lock         (icb_cmd_lock  ),                     
  .o_icb_cmd_size         (icb_cmd_size  ),                     
  .o_icb_cmd_usr          (icb_cmd_user  ),

  .o_icb_rsp_valid        (icb_rsp_valid  ),                     
  .o_icb_rsp_ready        (icb_rsp_ready  ),                     
  .o_icb_rsp_err          (icb_rsp_err    ),                     
  .o_icb_rsp_excl_ok      (icb_rsp_excl_ok),                     
  .o_icb_rsp_rdata        (icb_rsp_rdata  ),                    
  .o_icb_rsp_usr          ({USR_W{1'b0}}  ), 

  .i_bus_icb_cmd_sel_vec  (ccxw7l8izxzjj14ozqkgvvyd6) ,

  .i_bus_icb_cmd_ready    (w0hjg2xow0ymilw7bcxpm2l ),
  .i_bus_icb_cmd_valid    (k1_j5ubhqqpfrl3p0bi186va9 ),
  .i_bus_icb_cmd_read     (a_dm6kd_qbw2cv84wtboltif01  ),
  .i_bus_icb_cmd_addr     (xzpsiztjmn62eb967x1xkc6  ),
  .i_bus_icb_cmd_wdata    (ae00o9ay050qc5d5zxf18282b92 ),
  .i_bus_icb_cmd_wmask    (puxr8jzij0m30qcwmdz2sufl51 ),
  .i_bus_icb_cmd_burst    (sxjmcdip1m7ighns0k5aue59fj ),
  .i_bus_icb_cmd_beat     (noyjdh392j1x0s9g1b_lk  ),
  .i_bus_icb_cmd_excl     (wspjbjcpf459zy17qhyz8jmqy7  ),
  .i_bus_icb_cmd_lock     (s6vj39lt1yt7f1ytk3pr3 ), 
  .i_bus_icb_cmd_size     (y7jg1o7n3jl52fxr0isdv8 ), 
  .i_bus_icb_cmd_usr      (w8o2oxw46tp1zf4rujrx4zyxw  ), 

  .i_bus_icb_rsp_valid    (qkiytqsa_fo9x5ls7yb_x1k2 ) ,
  .i_bus_icb_rsp_ready    (idw2i93am7m9wy_5hzipgymj5k3 ) ,
  .i_bus_icb_rsp_err      (wzmdtyq65i82w_tt0juwqle)    ,
  .i_bus_icb_rsp_excl_ok  (kz10yoaxkacgm38dwv37tl2ixfv),
  .i_bus_icb_rsp_rdata    (fyvkbec2dn4rlcslyiyttfrx ) ,
  .i_bus_icb_rsp_usr      (od5a1yudx9bmyqpwleexh4h9) ,

  .clk                    (clk  )                     ,
  .rst_n                  (rst_n)
  );


  assign icb_cmd_sel  = icb_cmd_valid ; 






  wire stljptivoymm8t1vi8 = axi_arvalid | axi_awvalid | axi_wvalid | axi_rvalid | axi_bvalid ;

  assign axi_slave_active = (stljptivoymm8t1vi8 | hivak1ik74xuevh7l0f_4513 | ix0lsijxqslj1lxk0dtiy2fsq | l0_5x2ohgu6m77k54mg);



endmodule







module  ux607_gnrl_axi2icb_write # (
  parameter BUFFER_DP = 2,
  parameter AW = 32,
  parameter DW = 32,
  parameter MW = 4,
  parameter ALLOW_BURST = 0,
  parameter FIFO_OUTS_NUM = 4,
  parameter ID_W = 4,
  parameter USR_W = 1
) (

  output                           axi_awready,
  input                            axi_awvalid,
  input [ID_W-1:0]        axi_awid,
  input [AW-1:0]      axi_awaddr,
  input [7:0]                      axi_awlen,
  input [2:0]                      axi_awsize,
  input [1:0]                      axi_awburst,
  input                            axi_awlock,
  input [3:0]                      axi_awcache,
  input [2:0]                      axi_awprot,
  input [3:0]                      axi_awqos,
  input [3:0]                      axi_awregion,
  input [USR_W-1:0]          axi_awuser, 

  output                           axi_wready,
  input                            axi_wvalid,
  input [ID_W-1:0]        axi_wid,
  input [DW-1:0]           axi_wdata,
  input [MW-1:0]        axi_wstrb,
  input                            axi_wlast,

  input                            axi_bready,
  output                           axi_bvalid,
  output [ID_W-1:0]       axi_bid,
  output [1:0]                     axi_bresp,

  output                           icb_wcmd_valid,
  input                            icb_wcmd_ready,
  output [AW-1:0]                  icb_wcmd_addr,
  output                           icb_wcmd_read, 
  output [DW-1:0]                  icb_wcmd_wdata,
  output [MW-1:0]                  icb_wcmd_wmask,
  output [2:0]                     icb_wcmd_burst,
  output [1:0]                     icb_wcmd_beat,
  output                           icb_wcmd_lock,
  output                           icb_wcmd_excl,
  output [1:0]                     icb_wcmd_size,
  output [USR_W-1:0]               icb_wcmd_usr,

  input                            icb_wrsp_valid,
  output                           icb_wrsp_ready,
  input                            icb_wrsp_err,
  input                            icb_wrsp_excl_ok,

  input                            axi_bus_clk_en,

  output                           axi2icb_write_active,

  input  clk,
  input  rst_n
  );



  assign icb_wcmd_lock = 1'b0;


    localparam m2obdmbm7lrjdsvysr = ID_W+AW+8+3+2+1+4+3+4+4+USR_W;
    wire [m2obdmbm7lrjdsvysr-1:0] dcvm0a_dxcft7n72yw = {
                                             axi_awid    ,  
                                             axi_awaddr  ,
                                             axi_awlen   ,
                                             axi_awsize  ,
                                             axi_awburst ,
                                             axi_awlock  ,
                                             axi_awcache ,
                                             axi_awprot  ,
                                             axi_awqos   ,
                                             axi_awregion,
                                             axi_awuser   
                                            };
    wire [ID_W-1:0]    blcn1yvo8nt6t6xf    ; 
    wire [AW-1:0]  z1671m7vv3evkpne  ; 
    wire [7:0]                  vo3k0n9qzg9ph6m46   ; 
    wire [2:0]                  ar_rw9t62wsvom697rvi2  ; 
    wire [1:0]                  ixnmstf7hr62573gcwlidw ; 
    wire                        hby4soro9kdqiigwkgo  ; 
    wire [3:0]                  wd3g7w63oc93a6iv3ji ; 
    wire [2:0]                  oxns2iuot0xry0uk  ; 
    wire [3:0]                  be7f9j0jjk4nmku   ; 
    wire [3:0]                  to6cvmot263x2om2n8l8;
    wire [USR_W-1:0]      fml_np4pbuynvqwadm23  ; 

    wire [m2obdmbm7lrjdsvysr-1:0] z4hb9xf1ol2vbztjx ;

    assign  { 
              blcn1yvo8nt6t6xf    , 
              z1671m7vv3evkpne  , 
              vo3k0n9qzg9ph6m46   , 
              ar_rw9t62wsvom697rvi2  , 
              ixnmstf7hr62573gcwlidw , 
              hby4soro9kdqiigwkgo  , 
              wd3g7w63oc93a6iv3ji , 
              oxns2iuot0xry0uk  , 
              be7f9j0jjk4nmku   , 
              to6cvmot263x2om2n8l8,
              fml_np4pbuynvqwadm23    
            } = z4hb9xf1ol2vbztjx ;

    wire gut_a3vqb7tl6ve4jp1x0 ;    
    wire bkksqlu67uceqisenl ; 
    wire rsk12alll4cr ; 

    vq28fpkbg0dxljs8bf0k # (
      .hejad2_b4dywimoxw5 (1),
      .evi4vkasjp742kf4 (0),
      .mhdlk  (BUFFER_DP),
      .onr7l  (m2obdmbm7lrjdsvysr)
    ) mv67njo098wtgffd(
    .geml8twgru(axi_bus_clk_en), 
    .bw6ftrau0(axi_awvalid  ), 
    .eef2g8(axi_awready  ), 
    .qbjvs30wtb(dcvm0a_dxcft7n72yw),

    .td5hjljc_(1'b1),
    .wqljp(gut_a3vqb7tl6ve4jp1x0), 
    .h9378(bkksqlu67uceqisenl), 
    .dqgck5s(z4hb9xf1ol2vbztjx    ),

    .i0lklnhw28rc7dj(rsk12alll4cr),
    .gf33atgy  (clk  ),
    .ru_wi(rst_n)  
   );

    localparam z9_r__ensx481kjfcq_ = ID_W+DW+MW+1;
    wire [z9_r__ensx481kjfcq_-1:0] ry3h44oh0crn1dmx = {
                                             axi_wid        ,  
                                             axi_wdata      , 
                                             axi_wstrb      , 
                                             axi_wlast        
                                            };
    wire [ID_W-1:0]    eli2g_3s8txx4    ; 
    wire [DW-1:0]       on8q6jgldwnfhnxl  ; 
    wire [MW-1:0]    v2_7ykv6_69q6p5  ; 
    wire                        xxdd8qrecxg1h0_nwe  ; 

    wire [z9_r__ensx481kjfcq_-1:0] xc62eedzo559b ;

    assign  { 
              eli2g_3s8txx4    , 
              on8q6jgldwnfhnxl  , 
              v2_7ykv6_69q6p5  , 
              xxdd8qrecxg1h0_nwe    
            } = xc62eedzo559b ;

    wire iydg6q2hl9i8dyd18x_01 ;    
    wire miyqp0up17we11liuz_sz ; 
    wire bjd0di16hl3k6r37 ; 

    vq28fpkbg0dxljs8bf0k # (
      .hejad2_b4dywimoxw5 (1),
      .evi4vkasjp742kf4 (0),
      .mhdlk  (BUFFER_DP),
      .onr7l  (z9_r__ensx481kjfcq_)
    ) jfz87di8otj6(
    .geml8twgru(axi_bus_clk_en),
    .bw6ftrau0(axi_wvalid  ), 
    .eef2g8(axi_wready  ), 
    .qbjvs30wtb(ry3h44oh0crn1dmx),

    .td5hjljc_(1'b1),
    .wqljp(iydg6q2hl9i8dyd18x_01), 
    .h9378(miyqp0up17we11liuz_sz), 
    .dqgck5s(xc62eedzo559b    ),

    .i0lklnhw28rc7dj(bjd0di16hl3k6r37),
    .gf33atgy  (clk  ),
    .ru_wi(rst_n)  
   );

  wire izooaeazskwyqjnotwclm74;
  wire u7w75sbjtfwd1wf2aw84p;
  wire hgdqv2pzcv388wrnwbg;

  assign bkksqlu67uceqisenl     = hgdqv2pzcv388wrnwbg & izooaeazskwyqjnotwclm74;
  assign u7w75sbjtfwd1wf2aw84p = hgdqv2pzcv388wrnwbg & gut_a3vqb7tl6ve4jp1x0    ;

  ux607_gnrl_axi2icb_aw # (
    .AW (AW),
    .DW (DW),
    .MW (MW),
    .ALLOW_BURST(ALLOW_BURST),
    .ID_W (ID_W),
    .USR_W (USR_W)
  ) d7n4vmtvx890f9lbs0s(
    .axi_awready  (izooaeazskwyqjnotwclm74 ),
    .axi_awvalid  (u7w75sbjtfwd1wf2aw84p ),
    .axi_awid     (blcn1yvo8nt6t6xf    ),
    .axi_awaddr   (z1671m7vv3evkpne  ),
    .axi_awlen    (vo3k0n9qzg9ph6m46   ),
    .axi_awsize   (ar_rw9t62wsvom697rvi2  ),
    .axi_awburst  (ixnmstf7hr62573gcwlidw ),
    .axi_awlock   (hby4soro9kdqiigwkgo  ),
    .axi_awcache  (wd3g7w63oc93a6iv3ji ),
    .axi_awprot   (oxns2iuot0xry0uk  ),
    .axi_awqos    (be7f9j0jjk4nmku   ),
    .axi_awregion (to6cvmot263x2om2n8l8),
    .axi_awuser   (fml_np4pbuynvqwadm23),

    .axi_wready   (miyqp0up17we11liuz_sz),
    .axi_wvalid   (iydg6q2hl9i8dyd18x_01),
    .axi_wid      (eli2g_3s8txx4   ),
    .axi_wdata    (on8q6jgldwnfhnxl ),
    .axi_wstrb    (v2_7ykv6_69q6p5 ),
    .axi_wlast    (xxdd8qrecxg1h0_nwe ),


    .icb_wcmd_valid (icb_wcmd_valid),
    .icb_wcmd_ready (icb_wcmd_ready),
    .icb_wcmd_addr  (icb_wcmd_addr ), 
    .icb_wcmd_read  (icb_wcmd_read ), 
    .icb_wcmd_wdata (icb_wcmd_wdata),
    .icb_wcmd_wmask (icb_wcmd_wmask),
    .icb_wcmd_burst (icb_wcmd_burst),
    .icb_wcmd_beat  (icb_wcmd_beat ),
    .icb_wcmd_lock  (              ), 
    .icb_wcmd_excl  (icb_wcmd_excl ),
    .icb_wcmd_size  (icb_wcmd_size ),
    .icb_wcmd_usr   (icb_wcmd_usr  ), 

    .clk (clk),
    .rst_n (rst_n)
  );


    localparam yyi6c9dny1hxzp2 = ID_W+2;
    wire [ID_W-1:0]    i1jzyk_9b21dcj    ; 
    wire [1:0]                  xdqd89oa9qvwwg4sds  ; 


    wire [yyi6c9dny1hxzp2-1:0] sqnwox85n74r6s = {
                                             i1jzyk_9b21dcj  ,  
                                             xdqd89oa9qvwwg4sds        
                                            };
    wire [yyi6c9dny1hxzp2-1:0] h7vmjmxtagdl ;

    assign  { 
              axi_bid    , 
              axi_bresp    
            } = h7vmjmxtagdl ;

    wire qo210ozz3j4a489cqcm ;    
    wire vky5ebeqk89g3ku81m ; 

    wire n1fr6ji8a3j ; 
    vq28fpkbg0dxljs8bf0k # (
      .hejad2_b4dywimoxw5 (0),
      .evi4vkasjp742kf4 (1),
      .mhdlk  (BUFFER_DP),
      .onr7l  (yyi6c9dny1hxzp2)
    ) q037u7vw0lyuh8(
    .geml8twgru(1'b1),
    .bw6ftrau0(qo210ozz3j4a489cqcm), 
    .eef2g8(vky5ebeqk89g3ku81m), 
    .qbjvs30wtb(sqnwox85n74r6s    ),

    .td5hjljc_(axi_bus_clk_en),
    .wqljp(axi_bvalid  ), 
    .h9378(axi_bready  ), 
    .dqgck5s(h7vmjmxtagdl),

    .i0lklnhw28rc7dj(n1fr6ji8a3j),
    .gf33atgy  (clk  ),
    .ru_wi(rst_n)  
   );

  wire  mapugslkmxv351 ;
  wire  slggcmvgdj;
  dhou3hm297b56jmrnh31zua7 # (
    .nm_fj (AW),
    .onr7l (DW),
    .h1b (MW),
    .o7hawonznex2(ALLOW_BURST),
    .cibz (ID_W)
  ) ar26orka1ajeggs8o0dz9(
    .i5ydr9vb80xsvdjv2lm   (icb_wrsp_ready  ),
    .pimisco33wy7hvy   (icb_wrsp_valid  ),
    .nnqpeie69utf9y5h     (icb_wrsp_err    ),
    .o0d8x1ga2vq5_p_g__k (icb_wrsp_excl_ok),

    .nneek3ep5xykwl       (vky5ebeqk89g3ku81m),
    .g8khua4l0y77zjp       (qo210ozz3j4a489cqcm),
    .weop50xb_avne        (xdqd89oa9qvwwg4sds ),

    .mapugslkmxv351  (mapugslkmxv351),
    .slggcmvgdj (slggcmvgdj),

    .gf33atgy (clk),
    .ru_wi (rst_n)
  );

  wire r8aazdlqr6 = ((ixnmstf7hr62573gcwlidw == 2'b01) | (ixnmstf7hr62573gcwlidw == 2'b10)) & (~(vo3k0n9qzg9ph6m46 == 8'b0)) ;
  wire piygrateb  = hby4soro9kdqiigwkgo;

  wire qgbol4mpumx_qixqj72o3r;

  localparam nm9vgrzxtvpoz42 = 1+1+ID_W;
  ux607_gnrl_fifo # (
        .CUT_READY (1),
        .MSKO      (0),
        .DP  (FIFO_OUTS_NUM),
        .DW  (nm9vgrzxtvpoz42)
  ) isihu_4ctifhx (
        .i_vld(gut_a3vqb7tl6ve4jp1x0 && bkksqlu67uceqisenl ),
        .i_rdy(hgdqv2pzcv388wrnwbg),
        .i_dat({r8aazdlqr6,piygrateb, blcn1yvo8nt6t6xf}),
        .o_vld(qgbol4mpumx_qixqj72o3r),
        .o_rdy(qo210ozz3j4a489cqcm && vky5ebeqk89g3ku81m ),  
        .o_dat({slggcmvgdj,mapugslkmxv351, i1jzyk_9b21dcj}),  

        .clk  (clk),
        .rst_n(rst_n)
  );

   assign axi2icb_write_active = rsk12alll4cr | bjd0di16hl3k6r37 | n1fr6ji8a3j | qgbol4mpumx_qixqj72o3r;



endmodule








module  ux607_gnrl_axi2icb_read # (
  parameter BUFFER_DP = 2,
  parameter AW = 32,
  parameter DW = 32,
  parameter MW = 4,
  parameter ALLOW_BURST = 0,
  parameter FIFO_OUTS_NUM = 4,
  parameter ID_W = 4,
  parameter USR_W = 1
) (



  output                           axi_arready,
  input                            axi_arvalid,
  input [ID_W-1:0]        axi_arid,
  input [AW-1:0]      axi_araddr,
  input [7:0]                      axi_arlen,
  input [2:0]                      axi_arsize,
  input [1:0]                      axi_arburst,
  input                            axi_arlock,
  input [3:0]                      axi_arcache,
  input [2:0]                      axi_arprot,
  input [3:0]                      axi_arqos,
  input [3:0]                      axi_arregion,
  input [USR_W-1:0]          axi_aruser,


  input                            axi_rready,
  output                           axi_rvalid,
  output [ID_W-1:0]       axi_rid,
  output [DW-1:0]          axi_rdata,
  output [1:0]                     axi_rresp,
  output                           axi_rlast,


  output                           icb_rcmd_valid ,
  input                            icb_rcmd_ready ,
  output [AW-1:0]                  icb_rcmd_addr  ,
  output                           icb_rcmd_read  ,
  output [DW-1:0]                  icb_rcmd_wdata ,
  output [MW-1:0]                  icb_rcmd_wmask ,
  output [2:0]                     icb_rcmd_burst ,
  output [1:0]                     icb_rcmd_beat  ,
  output                           icb_rcmd_excl  ,             
  output [1:0]                     icb_rcmd_size  ,
  output [USR_W-1:0]               icb_rcmd_usr   ,

  output                           icb_rrsp_ready  , 
  input                            icb_rrsp_valid  , 
  input [DW-1:0]                   icb_rrsp_rdata  , 
  input                            icb_rrsp_err    , 
  input                            icb_rrsp_excl_ok, 

  input                            axi_bus_clk_en,

  output                           axi2icb_read_active,
  input clk  ,
  input rst_n  
  );




    localparam arybzlkhsez4dft4fc69 = ID_W+AW+8+3+2+1+4+3+4+4+USR_W;

    wire [arybzlkhsez4dft4fc69-1:0] a_3bnsvz8_htr = {
                                             axi_arid    ,  
                                             axi_araddr  ,
                                             axi_arlen   ,
                                             axi_arsize  ,
                                             axi_arburst ,
                                             axi_arlock  ,
                                             axi_arcache ,
                                             axi_arprot  ,
                                             axi_arqos   ,
                                             axi_arregion,
                                             axi_aruser   
                                            };
    wire [ID_W-1:0]    gcxgiwz42g2s_rurq    ; 
    wire [AW-1:0]  vda9tj7zj6kt6r_c  ; 
    wire [7:0]                  re7ej3htxwglcbr0a5   ; 
    wire [2:0]                  zphtb5ets8c3dkkn0l64t  ; 
    wire [1:0]                  ma8ggn0hb8nqcpgssh6 ; 
    wire                        utww_4dunp7eeoyx  ; 
    wire [3:0]                  luxzn6genvan6h9z9_y4kn ; 
    wire [2:0]                  sy4ydbfr_c26neik  ; 
    wire [3:0]                  st1clio7pqp88hlx01   ; 
    wire [3:0]                  wpadlaprzfxw8ph0ks1doh6;
    wire [USR_W-1:0]      kc5bx7zds9zvpnxu3  ; 

    wire [arybzlkhsez4dft4fc69-1:0] tfjmdd5q91e7pi ;

    assign  { 
              gcxgiwz42g2s_rurq    , 
              vda9tj7zj6kt6r_c  , 
              re7ej3htxwglcbr0a5   , 
              zphtb5ets8c3dkkn0l64t  , 
              ma8ggn0hb8nqcpgssh6 , 
              utww_4dunp7eeoyx  , 
              luxzn6genvan6h9z9_y4kn , 
              sy4ydbfr_c26neik  , 
              st1clio7pqp88hlx01   , 
              wpadlaprzfxw8ph0ks1doh6,
              kc5bx7zds9zvpnxu3    
            } = tfjmdd5q91e7pi ;

    wire fjgjb9yp3uixhp0ce ;    
    wire qr_6a5_o0x6yec2s5f ; 
    wire exqprj8_xrv3z ; 

    vq28fpkbg0dxljs8bf0k # (
      .hejad2_b4dywimoxw5 (1),
      .evi4vkasjp742kf4 (0),
      .mhdlk  (BUFFER_DP),
      .onr7l  (arybzlkhsez4dft4fc69)
    ) aprrbyg85wsud_3ri_(
    .geml8twgru(axi_bus_clk_en), 

    .bw6ftrau0(axi_arvalid      ), 
    .eef2g8(axi_arready      ), 
    .qbjvs30wtb(a_3bnsvz8_htr    ),

    .td5hjljc_(1'b1), 

    .wqljp(fjgjb9yp3uixhp0ce), 
    .h9378(qr_6a5_o0x6yec2s5f), 
    .dqgck5s(tfjmdd5q91e7pi    ),

    .i0lklnhw28rc7dj(exqprj8_xrv3z),
    .gf33atgy  (clk  ),
    .ru_wi(rst_n)  
   );


  wire m1rwfy550xbjnt651yvs5;
  wire t5c_79ikvtdn1cglfh5b_;
  wire bouo8ouss5ujfkm013;

  assign qr_6a5_o0x6yec2s5f     = bouo8ouss5ujfkm013 & m1rwfy550xbjnt651yvs5;
  assign t5c_79ikvtdn1cglfh5b_ = bouo8ouss5ujfkm013 & fjgjb9yp3uixhp0ce;

  ux607_gnrl_axi2icb_ar # (
    .AW (AW),
    .DW (DW),
    .MW (MW),
    .ALLOW_BURST(ALLOW_BURST),
    .ID_W (ID_W),
    .USR_W (USR_W)  
  ) iiwrcmvoh63ahvdljk(
     .axi_arready  (m1rwfy550xbjnt651yvs5 ),
     .axi_arvalid  (t5c_79ikvtdn1cglfh5b_ ),
     .axi_arid     (gcxgiwz42g2s_rurq    ),
     .axi_araddr   (vda9tj7zj6kt6r_c  ),
     .axi_arlen    (re7ej3htxwglcbr0a5   ),
     .axi_arsize   (zphtb5ets8c3dkkn0l64t  ),
     .axi_arburst  (ma8ggn0hb8nqcpgssh6 ),
     .axi_arlock   (utww_4dunp7eeoyx  ),
     .axi_arcache  (luxzn6genvan6h9z9_y4kn ),
     .axi_arprot   (sy4ydbfr_c26neik  ),
     .axi_arqos    (st1clio7pqp88hlx01   ),
     .axi_arregion (wpadlaprzfxw8ph0ks1doh6),
     .axi_aruser   (kc5bx7zds9zvpnxu3), 


     .icb_rcmd_valid (icb_rcmd_valid),
     .icb_rcmd_ready (icb_rcmd_ready),
     .icb_rcmd_addr  (icb_rcmd_addr ), 
     .icb_rcmd_read  (icb_rcmd_read ), 
     .icb_rcmd_wdata (icb_rcmd_wdata),
     .icb_rcmd_wmask (icb_rcmd_wmask),
     .icb_rcmd_burst (icb_rcmd_burst),
     .icb_rcmd_beat  (icb_rcmd_beat ),
     .icb_rcmd_lock  (              ), 
     .icb_rcmd_excl  (icb_rcmd_excl ),
     .icb_rcmd_size  (icb_rcmd_size ),
     .icb_rcmd_usr   (icb_rcmd_usr  ),

     .clk   (clk),
     .rst_n (rst_n)
  );


    localparam d4rf2qjcejeat0ug = ID_W+DW+2+1;
    wire [ID_W-1:0]    aqiu5iaab6p2ej    ; 
    wire [DW-1:0]       g32u54xok1emh7w  ; 
    wire [1:0]                  am6dug03mtmj5vrm5uuj  ; 
    wire                        bviecamw6kx251h0qee0  ; 

    wire [d4rf2qjcejeat0ug-1:0] wcx8l6zmds1l2z = {
                                             aqiu5iaab6p2ej    ,
                                             g32u54xok1emh7w  ,
                                             am6dug03mtmj5vrm5uuj  ,
                                             bviecamw6kx251h0qee0   
                                            };
    wire [d4rf2qjcejeat0ug-1:0] oyznb90rr_pu0l ;

    assign  { 
              axi_rid        ,  
              axi_rdata      ,  
              axi_rresp      ,  
              axi_rlast         
            } = oyznb90rr_pu0l ;

    wire z6i49kyfixjznjy19ki ;    
    wire qj3f7kzhtmxe8lyb ; 
    wire h__kt0wtrbia ; 

    vq28fpkbg0dxljs8bf0k # (
      .hejad2_b4dywimoxw5 (0),
      .evi4vkasjp742kf4 (1),
      .mhdlk  (BUFFER_DP),
      .onr7l  (d4rf2qjcejeat0ug)
    ) q35nsujqlr5e2ql(
    .geml8twgru(1'b1),
    .bw6ftrau0(z6i49kyfixjznjy19ki), 
    .eef2g8(qj3f7kzhtmxe8lyb), 
    .qbjvs30wtb(wcx8l6zmds1l2z    ),

    .td5hjljc_(axi_bus_clk_en),
    .wqljp(axi_rvalid  ), 
    .h9378(axi_rready  ), 
    .dqgck5s(oyznb90rr_pu0l),

    .i0lklnhw28rc7dj(h__kt0wtrbia),
    .gf33atgy  (clk  ),
    .ru_wi(rst_n)  
   );


  wire  rhakurg97nzjtd ;
  wire  wnegzux_m31q;
  fpg_i1rl2go50l8gnsv # (
    .nm_fj (AW),
    .onr7l (DW),
    .h1b (MW),
    .o7hawonznex2(ALLOW_BURST),
    .cibz (ID_W)
  ) dcvmc66_7ff3cw8120j(
    .ee0gaim_5o2cowj8cc   (icb_rrsp_ready  ),
    .iy0c52aia8jldt99i   (icb_rrsp_valid  ),
    .wtmpbfqxajai_cc   (icb_rrsp_rdata  ),
    .dt4m1v705h0fe     (icb_rrsp_err    ),
    .t_xyazag81f8t2zmg8b4 (icb_rrsp_excl_ok),

    .hjstsi51gm       (qj3f7kzhtmxe8lyb),
    .onpqhy0s69       (z6i49kyfixjznjy19ki),
    .aw7xjbi          (                ),
    .z0cc2y_uzoh_        (g32u54xok1emh7w ),
    .y8tc_vywu82ugn        (am6dug03mtmj5vrm5uuj ),
    .o2h9d51o6m6        (bviecamw6kx251h0qee0 ),

    .rhakurg97nzjtd        (rhakurg97nzjtd     ),
    .wnegzux_m31q       (wnegzux_m31q    ),

    .gf33atgy   (clk          ),
    .ru_wi (rst_n)
  );

  wire w3rlzdtdaan = ((ma8ggn0hb8nqcpgssh6 == 2'b01) | (ma8ggn0hb8nqcpgssh6 == 2'b10)) & (~(re7ej3htxwglcbr0a5 == 8'b0)) ;
  wire qe8p6_qys3vlb  = utww_4dunp7eeoyx;

  wire ciu5unao5uvd2mq6r7st83u;

  localparam jfjrr2q0m19ir7royv = 1+1+ID_W;
  ux607_gnrl_fifo # (
        .CUT_READY (1),
        .MSKO      (0),
        .DP  (FIFO_OUTS_NUM), 
        .DW  (jfjrr2q0m19ir7royv)
  ) wbz08fovrvbnwsq0 (
        .i_vld(fjgjb9yp3uixhp0ce && qr_6a5_o0x6yec2s5f ), 
        .i_rdy(bouo8ouss5ujfkm013),
        .i_dat({w3rlzdtdaan,qe8p6_qys3vlb, gcxgiwz42g2s_rurq}),
        .o_vld(ciu5unao5uvd2mq6r7st83u),
        .o_rdy(z6i49kyfixjznjy19ki && qj3f7kzhtmxe8lyb && bviecamw6kx251h0qee0 ),  
        .o_dat({wnegzux_m31q,rhakurg97nzjtd, aqiu5iaab6p2ej}),  

        .clk  (clk),
        .rst_n(rst_n)
  );


  assign axi2icb_read_active = exqprj8_xrv3z | h__kt0wtrbia | ciu5unao5uvd2mq6r7st83u;


endmodule








module ux607_gnrl_axi2icb_ar # (
  parameter AW = 32,
  parameter DW = 32,
  parameter MW = 4,
  parameter ALLOW_BURST = 0,
  parameter ID_W = 4, 
  parameter USR_W = 1
) (
  output                         axi_arready,
  input                          axi_arvalid,
  input [ID_W-1:0]               axi_arid,
  input [AW-1:0]                 axi_araddr,
  input [7:0]                    axi_arlen,
  input [2:0]                    axi_arsize,
  input [1:0]                    axi_arburst,
  input                          axi_arlock,
  input [3:0]                    axi_arcache,
  input [2:0]                    axi_arprot,
  input [3:0]                    axi_arqos,
  input [3:0]                    axi_arregion,
  input [USR_W-1:0]              axi_aruser,

  output                         icb_rcmd_valid,
  input                          icb_rcmd_ready,
  output [AW-1:0]                icb_rcmd_addr, 
  output                         icb_rcmd_read, 
  output [DW-1:0]                icb_rcmd_wdata,
  output [MW-1:0]                icb_rcmd_wmask,
  output [2:0]                   icb_rcmd_burst,
  output [1:0]                   icb_rcmd_beat,
  output                         icb_rcmd_lock,
  output                         icb_rcmd_excl,
  output [1:0]                   icb_rcmd_size,
  output [USR_W-1:0]             icb_rcmd_usr,

  input                         clk,
  input                         rst_n
  );

  wire       afkj5yhhtctg6s;
  wire [2:0] g85wmlhjsfg_;
  wire [2:0] qv6grfmv4g0b663;
  wire       d767w05jxusx0gx6;
  wire       w3rlzdtdaan;
  wire       bvx56ynjv2g4li;

  wire w_4lt6kv0fqfp1onbi;
  wire [1:0] teg4mq_q8o7732him0;
  wire [USR_W-1:0] cg17l88hjzg09y1n;
  wire [AW-1:0] kse881ijv015_p;
  wire jvzqm8i9b77;

  assign w3rlzdtdaan = axi_arvalid  & ((axi_arburst == 2'b01) | (axi_arburst == 2'b10)) & (~(axi_arlen == 8'b0)) ;
  assign bvx56ynjv2g4li = (g85wmlhjsfg_ != 3'b0);
  generate
    if (ALLOW_BURST == 0) begin :bd14fahfursl
  assign afkj5yhhtctg6s =1'b0;
  assign g85wmlhjsfg_ = 3'b0;
  assign qv6grfmv4g0b663 = 3'b0;
  assign d767w05jxusx0gx6 = 1'b0;
  assign jvzqm8i9b77       = 1'b0;
  assign w_4lt6kv0fqfp1onbi  = 1'b0;
  assign teg4mq_q8o7732him0  = 2'b0;
  assign cg17l88hjzg09y1n  = {USR_W{1'b0}};
  assign kse881ijv015_p  = {AW{1'b0}};
    end
    else begin :j_7fmjdgwqmy5
  assign qv6grfmv4g0b663 = afkj5yhhtctg6s ? 3'b0 : (g85wmlhjsfg_ + 3'b1);
  assign afkj5yhhtctg6s = ((DW==32) && (g85wmlhjsfg_==3'b111)) || ((DW==64) && (g85wmlhjsfg_==3'b011));

  assign d767w05jxusx0gx6 = (w3rlzdtdaan || bvx56ynjv2g4li) && icb_rcmd_valid && icb_rcmd_ready;
  assign jvzqm8i9b77 = w3rlzdtdaan && icb_rcmd_valid && icb_rcmd_ready && (g85wmlhjsfg_ == 3'b0);
  ux607_gnrl_dfflr #(3) azqo5a_gl8snymahf0 (d767w05jxusx0gx6, qv6grfmv4g0b663, g85wmlhjsfg_, clk, rst_n);
  ux607_gnrl_dffl #(1) f7kyai3p09je2 ( jvzqm8i9b77, axi_arlock, w_4lt6kv0fqfp1onbi, clk, rst_n); 
  ux607_gnrl_dffl #(2) zhxi0diz1cwc89d ( jvzqm8i9b77, axi_arsize[1:0], teg4mq_q8o7732him0, clk, rst_n); 
  ux607_gnrl_dffl #(USR_W) oqi5nue_c3jjqid4 ( jvzqm8i9b77, axi_aruser, cg17l88hjzg09y1n, clk, rst_n); 
  ux607_gnrl_dffl #(AW) vp0305x7ez6zpw_ ( jvzqm8i9b77, axi_araddr, kse881ijv015_p, clk, rst_n); 
    end
  endgenerate

  assign axi_arready   = icb_rcmd_ready && (!bvx56ynjv2g4li);

  assign icb_rcmd_valid   = axi_arvalid  || bvx56ynjv2g4li;
  assign icb_rcmd_read    = 1'b1; 
  assign icb_rcmd_wdata   = {DW{1'b0}};
  assign icb_rcmd_wmask   = {MW{1'b0}};

  assign icb_rcmd_lock    = 1'b0; 
  assign icb_rcmd_excl    = bvx56ynjv2g4li ? w_4lt6kv0fqfp1onbi : axi_arlock;
  assign icb_rcmd_size    = bvx56ynjv2g4li ? teg4mq_q8o7732him0[1:0] : axi_arsize[1:0];
  generate
    if (ALLOW_BURST == 0) begin :aqxqd0hfmq7dkb
  assign icb_rcmd_burst = 3'b0;
  assign icb_rcmd_beat  = 2'b0;
  assign icb_rcmd_addr  = axi_araddr;
    end
    else begin :ifts0ro55hlf5mzjq
  wire [2:0] ecgi_6q1ku_1o;
  wire       a0igv262zce64zbc3 = d767w05jxusx0gx6;


  wire [2:0] u32wwykc7v8xy898 = (!bvx56ynjv2g4li) ? (axi_araddr[4:2] + DW[7:5])
                                              : (ecgi_6q1ku_1o + DW[7:5]);
  ux607_gnrl_dfflr #(3) cwt2s31zb5t64mp1p3d (a0igv262zce64zbc3, u32wwykc7v8xy898, ecgi_6q1ku_1o, clk, rst_n);

  assign icb_rcmd_burst = (!w3rlzdtdaan && !bvx56ynjv2g4li) ? 3'b000 : 
                          (DW == 32)                     ? 3'b101 :
                                                           3'b010 ;
  assign icb_rcmd_beat  = (!w3rlzdtdaan && !bvx56ynjv2g4li) ? 2'b00 : 
                          (afkj5yhhtctg6s)                   ? 2'b10 :
                                                           2'b01 ;
  assign icb_rcmd_addr  = (!bvx56ynjv2g4li) ? axi_araddr                          : 
                          (DW == 32)     ? {kse881ijv015_p[AW-1:5],ecgi_6q1ku_1o,2'b0} :
                                           {kse881ijv015_p[AW-1:5],ecgi_6q1ku_1o,2'b0} ;
    end
  endgenerate
  assign icb_rcmd_usr   = bvx56ynjv2g4li ? cg17l88hjzg09y1n : axi_aruser;

endmodule







module ux607_gnrl_axi2icb_aw # (
  parameter AW = 32,
  parameter DW = 32,
  parameter MW = 4,
  parameter ALLOW_BURST = 0,
  parameter ID_W = 4,
  parameter USR_W = 1
) (
  output                         axi_awready,
  input                          axi_awvalid,
  input [ID_W-1:0]               axi_awid,
  input [AW-1:0]                 axi_awaddr,
  input [7:0]                    axi_awlen,
  input [2:0]                    axi_awsize,
  input [1:0]                    axi_awburst,
  input                          axi_awlock,
  input [3:0]                    axi_awcache,
  input [2:0]                    axi_awprot,
  input [3:0]                    axi_awqos,
  input [3:0]                    axi_awregion,
  input [USR_W-1:0]              axi_awuser,

  output                         axi_wready,
  input                          axi_wvalid,
  input [ID_W-1:0]               axi_wid,
  input [DW-1:0]                 axi_wdata,
  input [MW-1:0]                 axi_wstrb,
  input                          axi_wlast,

  output                         icb_wcmd_valid,
  input                          icb_wcmd_ready,
  output [AW-1:0]                icb_wcmd_addr, 
  output                         icb_wcmd_read, 
  output [DW-1:0]                icb_wcmd_wdata,
  output [MW-1:0]                icb_wcmd_wmask,
  output [2:0]                   icb_wcmd_burst,
  output [1:0]                   icb_wcmd_beat,
  output                         icb_wcmd_lock,
  output                         icb_wcmd_excl,
  output [1:0]                   icb_wcmd_size,
  output [USR_W-1:0]             icb_wcmd_usr,

  input                         clk,
  input                         rst_n
  );

  wire       afkj5yhhtctg6s;
  wire [2:0] g85wmlhjsfg_;
  wire [2:0] qv6grfmv4g0b663;
  wire       d767w05jxusx0gx6;
  wire       r8aazdlqr6;
  wire       vydagkrnnuoyq6j;

  wire p0gcuood618ubg;
  wire [2:0] lmn39rifwgsf99v22;
  wire [USR_W-1:0] jaxeeknuvin5uw;
  wire [AW-1:0] c__5jqkrm6qsue75x;
  wire jvzqm8i9b77;

  assign r8aazdlqr6 = axi_awvalid  & ((axi_awburst == 2'b01) | (axi_awburst == 2'b10)) & (~(axi_awlen == 8'b0)) ;
  assign vydagkrnnuoyq6j = (g85wmlhjsfg_ != 3'b0);
  generate
    if (ALLOW_BURST == 0) begin :n06sz1b1033n0489fq
  assign afkj5yhhtctg6s =1'b0;
  assign g85wmlhjsfg_ = 3'b0;
  assign qv6grfmv4g0b663 = 3'b0;
  assign d767w05jxusx0gx6 = 1'b0;
  assign jvzqm8i9b77       = 1'b0;
  assign p0gcuood618ubg  = 1'b0;
  assign lmn39rifwgsf99v22  = 3'b0;
  assign jaxeeknuvin5uw  = {USR_W{1'b0}};
  assign c__5jqkrm6qsue75x  = {AW{1'b0}};
    end
    else begin :eydxyrfp1w_48m1za
  assign qv6grfmv4g0b663 = afkj5yhhtctg6s ? 3'b0 : (g85wmlhjsfg_ + 3'b1);
  assign afkj5yhhtctg6s = ((DW==32) && (g85wmlhjsfg_==3'b111)) || ((DW==64) && (g85wmlhjsfg_==3'b011));

  assign d767w05jxusx0gx6 = (r8aazdlqr6 || vydagkrnnuoyq6j) && icb_wcmd_valid && icb_wcmd_ready;
  assign jvzqm8i9b77 = r8aazdlqr6 && icb_wcmd_valid && icb_wcmd_ready && (g85wmlhjsfg_ == 3'b0);
  ux607_gnrl_dfflr #(3) azqo5a_gl8snymahf0 (d767w05jxusx0gx6, qv6grfmv4g0b663, g85wmlhjsfg_, clk, rst_n);
  ux607_gnrl_dffl #(1) n4e9isv717t ( jvzqm8i9b77, axi_awlock, p0gcuood618ubg, clk, rst_n); 
  ux607_gnrl_dffl #(3) z69nt03um6lb ( jvzqm8i9b77, axi_awsize, lmn39rifwgsf99v22, clk, rst_n); 
  ux607_gnrl_dffl #(USR_W) zwipqefm4amkfrvd ( jvzqm8i9b77, axi_awuser, jaxeeknuvin5uw, clk, rst_n); 
  ux607_gnrl_dffl #(AW) drfd3kum8yt9b ( jvzqm8i9b77, axi_awaddr, c__5jqkrm6qsue75x, clk, rst_n); 
    end
  endgenerate


  assign axi_awready   = icb_wcmd_ready && (!vydagkrnnuoyq6j)  && axi_wvalid;
  assign axi_wready    = icb_wcmd_ready && (vydagkrnnuoyq6j || axi_awvalid);

  assign icb_wcmd_valid   = (axi_awvalid || vydagkrnnuoyq6j) && axi_wvalid ;

  assign icb_wcmd_read    = 1'b0; 
  assign icb_wcmd_wdata   = axi_wdata;
  assign icb_wcmd_wmask   = axi_wstrb;

  assign icb_wcmd_lock    = 1'b0;
  assign icb_wcmd_excl    = vydagkrnnuoyq6j ? p0gcuood618ubg : axi_awlock;
  assign icb_wcmd_size    = vydagkrnnuoyq6j ? lmn39rifwgsf99v22[1:0] : axi_awsize[1:0];
  generate
    if (ALLOW_BURST == 0) begin :uoqdh0j6lpgs754osq
  assign icb_wcmd_burst = 3'b0;
  assign icb_wcmd_beat  = 2'b0;
  assign icb_wcmd_addr  = axi_awaddr;
    end
    else begin :zcctv8k35m7uza7b8_
  wire [2:0] ecgi_6q1ku_1o;
  wire       a0igv262zce64zbc3 = d767w05jxusx0gx6;


  wire [2:0] u32wwykc7v8xy898 = (!vydagkrnnuoyq6j) ? (axi_awaddr[4:2] + DW[7:5])
                                              : (ecgi_6q1ku_1o + DW[7:5]);
  ux607_gnrl_dfflr #(3) cwt2s31zb5t64mp1p3d (a0igv262zce64zbc3, u32wwykc7v8xy898, ecgi_6q1ku_1o, clk, rst_n);
  assign icb_wcmd_burst = (!r8aazdlqr6 && !vydagkrnnuoyq6j) ? 3'b000 : 
                          (DW == 32)                     ? 3'b101 :
                                                           3'b010 ;
  assign icb_wcmd_beat  = (!r8aazdlqr6 && !vydagkrnnuoyq6j) ? 2'b00 : 
                          (afkj5yhhtctg6s)                   ? 2'b10 :
                                                           2'b01 ;
  assign icb_wcmd_addr  = (!vydagkrnnuoyq6j) ? axi_awaddr                          : 
                          (DW == 32)     ? {c__5jqkrm6qsue75x[AW-1:5],ecgi_6q1ku_1o,2'b0} :
                                           {c__5jqkrm6qsue75x[AW-1:5],ecgi_6q1ku_1o,2'b0} ;
    end
  endgenerate
  assign icb_wcmd_usr   = vydagkrnnuoyq6j ? jaxeeknuvin5uw : axi_awuser;

endmodule






module fpg_i1rl2go50l8gnsv # (
  parameter nm_fj = 32,
  parameter onr7l = 32,
  parameter h1b = 4,
  parameter o7hawonznex2 = 0,
  parameter cibz = 4
) (
  output                        ee0gaim_5o2cowj8cc,
  input                         iy0c52aia8jldt99i,
  input [onr7l-1:0]                wtmpbfqxajai_cc,
  input                         dt4m1v705h0fe,
  input                         t_xyazag81f8t2zmg8b4,

  input                         hjstsi51gm,
  output                        onpqhy0s69,
  output [cibz-1:0]             aw7xjbi,
  output [onr7l-1:0]               z0cc2y_uzoh_,
  output [1:0]                  y8tc_vywu82ugn,
  output                        o2h9d51o6m6,

  input                         rhakurg97nzjtd,
  input                         wnegzux_m31q,

  input                         gf33atgy,
  input                         ru_wi
  );

  wire       afkj5yhhtctg6s;
  wire [2:0] g85wmlhjsfg_;
  wire [2:0] qv6grfmv4g0b663;
  wire       d767w05jxusx0gx6;

  generate
    if (o7hawonznex2 == 0) begin :zxeaazldzfnvzriytwpy
  assign afkj5yhhtctg6s =1'b0;
  assign g85wmlhjsfg_ = 3'b0;
  assign qv6grfmv4g0b663 = 3'b0;
  assign d767w05jxusx0gx6 = 1'b0;
    end
    else begin :ih5kfdapc0zecu9n2
  assign qv6grfmv4g0b663 = afkj5yhhtctg6s ? 3'b0 : (g85wmlhjsfg_ + 3'b1);
  assign afkj5yhhtctg6s = ((onr7l==32) && (g85wmlhjsfg_==3'b111)) || ((onr7l==64) && (g85wmlhjsfg_==3'b011));
  assign d767w05jxusx0gx6 = wnegzux_m31q && iy0c52aia8jldt99i && ee0gaim_5o2cowj8cc;
  ux607_gnrl_dfflr #(3) azqo5a_gl8snymahf0 (d767w05jxusx0gx6, qv6grfmv4g0b663, g85wmlhjsfg_, gf33atgy, ru_wi);
    end
  endgenerate

  assign ee0gaim_5o2cowj8cc   = hjstsi51gm ;

  assign onpqhy0s69       = iy0c52aia8jldt99i ;
  assign aw7xjbi          = {cibz{1'b0}};
  assign z0cc2y_uzoh_        = wtmpbfqxajai_cc;
  assign y8tc_vywu82ugn        = {dt4m1v705h0fe,rhakurg97nzjtd};
  assign o2h9d51o6m6        = (!wnegzux_m31q) || (wnegzux_m31q && afkj5yhhtctg6s);
endmodule






module dhou3hm297b56jmrnh31zua7 # (
  parameter nm_fj = 32,
  parameter onr7l = 32,
  parameter h1b = 4,
  parameter o7hawonznex2 = 0,
  parameter cibz = 4
) (
  output                        i5ydr9vb80xsvdjv2lm,
  input                         pimisco33wy7hvy,
  input                         nnqpeie69utf9y5h,
  input                         o0d8x1ga2vq5_p_g__k,

  input                         nneek3ep5xykwl,
  output                        g8khua4l0y77zjp,
  output [1:0]                  weop50xb_avne,

  input                         mapugslkmxv351,
  input                         slggcmvgdj,

  input                         gf33atgy,
  input                         ru_wi
  );

  wire       afkj5yhhtctg6s;
  wire [2:0] g85wmlhjsfg_;
  wire [2:0] qv6grfmv4g0b663;
  wire       d767w05jxusx0gx6;

  generate
    if (o7hawonznex2 == 0) begin :j8ozrjobogznhspk8o0
  assign afkj5yhhtctg6s =1'b0;
  assign g85wmlhjsfg_ = 3'b0;
  assign qv6grfmv4g0b663 = 3'b0;
  assign d767w05jxusx0gx6 = 1'b0;
    end
    else begin :d01pprd7v58cqzbjyh8
  assign qv6grfmv4g0b663 = afkj5yhhtctg6s ? 3'b0 : (g85wmlhjsfg_ + 3'b1);
  assign afkj5yhhtctg6s = ((onr7l==32) && (g85wmlhjsfg_==3'b111)) || ((onr7l==64) && (g85wmlhjsfg_==3'b011));
  assign d767w05jxusx0gx6 = slggcmvgdj && pimisco33wy7hvy && i5ydr9vb80xsvdjv2lm;
  ux607_gnrl_dfflr #(3) azqo5a_gl8snymahf0 (d767w05jxusx0gx6, qv6grfmv4g0b663, g85wmlhjsfg_, gf33atgy, ru_wi);
    end
  endgenerate

  assign i5ydr9vb80xsvdjv2lm   = (slggcmvgdj && !afkj5yhhtctg6s) || (nneek3ep5xykwl);

  assign g8khua4l0y77zjp       = pimisco33wy7hvy && (!slggcmvgdj || (slggcmvgdj && afkj5yhhtctg6s));
  generate
    if (o7hawonznex2 == 0 ) begin :wn4_6f37wzih2huwlwsr
  assign weop50xb_avne        = {nnqpeie69utf9y5h,mapugslkmxv351};
    end
    else begin :q59bauebnu1gljw4h8w
  wire [1:0]  aroydyww3h7l5g;
  wire [1:0]  w9gci50qpvdyh3;
  wire        zzjze2gy_tyj9;
  assign zzjze2gy_tyj9 = slggcmvgdj && pimisco33wy7hvy && i5ydr9vb80xsvdjv2lm && !afkj5yhhtctg6s;
  assign aroydyww3h7l5g = (g85wmlhjsfg_ == 0) ? {nnqpeie69utf9y5h,mapugslkmxv351}
                                             : (w9gci50qpvdyh3 | {nnqpeie69utf9y5h,mapugslkmxv351})
                                             ;
  ux607_gnrl_dffl #(2) hny1pp8yq1d (zzjze2gy_tyj9, aroydyww3h7l5g, w9gci50qpvdyh3, gf33atgy, ru_wi);
  assign weop50xb_avne        = ({2{slggcmvgdj}} & w9gci50qpvdyh3) | {nnqpeie69utf9y5h,mapugslkmxv351};
    end
  endgenerate
endmodule
























module tnzq74jtghufc(

  output                         byiw0kxjclrie9tn3h,

  input                          ndsqg7zrec89ncrv9yu3k,
  input                          eth8quxx9hhjhxr4u9k2s77f,
  output                         zw6mbnvv_8hcztypnytp87v_vy,
  input  [16-1:0]   l_s_khzs83700pzjuq3_obo44, 
  input                          tcrjx_8vlmtrlqjvk3tu, 
  input  [64-1:0]        y0jaju01t8mqh2ycz05limpxfu,
  input  [8-1:0]     x88dy7qz1z117o2jmbslutlpm,
  input                          kykdx6vx9n3hm7k6oybv,
  input                          b59iokn7e2645ocyqifdk6sp1,
  input  [1:0]                   xs2l1_f3yynnrl_rw2zbe,
  input                          tmqgi_fx924f3bq8ms4u8t0,
  input                          kyvscpwy0vljnwysfxqxb,
  input                          sl5cpfvi658e8pl6nh2cm4,
  
  output                         hf8rqlrzsk0e9ho4orde_r,
  input                          opns8_xijy8grr0gygeszh,
  output                         hng3_y3ldjtyu4a9n45  ,
  output                         y1ovf4ea_l0kgs84_pwk6czrs,
  output [64-1:0]        n6fa00b9i708mtqu7yc9wjvxip,

  
  
  
  
  
  
  
  
  output                         rqf8b5xxbw0n1_qaw,
  input                          ocwcf75wgxfb1bawe,
  output [16-1:0]   holgl43_yucp7f7l,
  output                         gy2sgn_1bpkac7msq3,
  output                         oyev1ipmdflkvxygwr,
  output                         ihknw7_lm_572tv6s,
  output                         o31l03k34sdhwt4lkazfa5, 
  output                         k3x026c5w9wldgp0z07b_, 
  output [64-1:0]        r_1u6q2lzkfus3o9nfl,
  output [8-1:0]     yff7wf8wth2vjkdjpr,
  output [1:0]                   wt4e4tlh0u_4cljr2j5f9,

  
  input                          o4wuryrcvw13y2v5m6b6u,
  input                          vnqegbzme0jutvf  ,
  input  [64-1:0]        p9mcc6npaw32uigcp6,
  input                          jdj122rbumyogtin6xpg97,
  output                         bt4howrm5xnf6u4fuwrum6,

  input  gf33atgy,
  input  ru_wi
  );

  


  localparam egb08sh4q_5pj = 1;

  localparam msjfsjsyuq0_ = egb08sh4q_5pj;	  

  localparam tjt5wdq_mmk = msjfsjsyuq0_;


  localparam vqmyiw_o188k = 2;
  
  localparam s3xvyho = 4;
  localparam y61y499cunmtec  = 0;
  localparam a69a9ho1_kmpwc58n  = 1;
  localparam zxf2f6zwhhxrms0dvq1  = 2;
  localparam qn77zdua2lv05_  = 3;

  wire [s3xvyho-1:0] wd3zc6palghmam9to3v2;


  wire [s3xvyho-1:0] syd0rz5l9shsemv;

  assign wd3zc6palghmam9to3v2[y61y499cunmtec ] = tmqgi_fx924f3bq8ms4u8t0;
  assign wd3zc6palghmam9to3v2[a69a9ho1_kmpwc58n ] = kyvscpwy0vljnwysfxqxb;
  assign wd3zc6palghmam9to3v2[qn77zdua2lv05_ ] = sl5cpfvi658e8pl6nh2cm4;
  assign wd3zc6palghmam9to3v2[zxf2f6zwhhxrms0dvq1 ] = 1'b0;

  
  assign o31l03k34sdhwt4lkazfa5 = syd0rz5l9shsemv[y61y499cunmtec ];
  assign oyev1ipmdflkvxygwr = syd0rz5l9shsemv[a69a9ho1_kmpwc58n ];
  assign ihknw7_lm_572tv6s = syd0rz5l9shsemv[qn77zdua2lv05_ ];
  assign k3x026c5w9wldgp0z07b_ = syd0rz5l9shsemv[zxf2f6zwhhxrms0dvq1 ];


  wire [tjt5wdq_mmk*1-1:0] k1_j5ubhqqpfrl3p0bi186va9;
  wire [tjt5wdq_mmk*1-1:0] w0hjg2xow0ymilw7bcxpm2l;
  wire [tjt5wdq_mmk*16-1:0] xzpsiztjmn62eb967x1xkc6;
  wire [tjt5wdq_mmk*1-1:0] a_dm6kd_qbw2cv84wtboltif01;
  wire [tjt5wdq_mmk*64-1:0] ae00o9ay050qc5d5zxf18282b92;
  wire [tjt5wdq_mmk*8-1:0] puxr8jzij0m30qcwmdz2sufl51;
  wire [tjt5wdq_mmk*1-1:0] s6vj39lt1yt7f1ytk3pr3;
  wire [tjt5wdq_mmk*1-1:0] wspjbjcpf459zy17qhyz8jmqy7;
  wire [tjt5wdq_mmk*2-1:0] y7jg1o7n3jl52fxr0isdv8;
  wire [tjt5wdq_mmk*s3xvyho-1:0] w8o2oxw46tp1zf4rujrx4zyxw;

  wire [tjt5wdq_mmk*1-1:0] qkiytqsa_fo9x5ls7yb_x1k2;
  wire [tjt5wdq_mmk*1-1:0] idw2i93am7m9wy_5hzipgymj5k3;
  wire [tjt5wdq_mmk*1-1:0] wzmdtyq65i82w_tt0juwqle;
  wire [tjt5wdq_mmk*1-1:0] kz10yoaxkacgm38dwv37tl2ixfv;
  wire [tjt5wdq_mmk*64-1:0] fyvkbec2dn4rlcslyiyttfrx;

  
  assign k1_j5ubhqqpfrl3p0bi186va9 =
      
                           {
                             eth8quxx9hhjhxr4u9k2s77f
                           } ;

  wire[tjt5wdq_mmk-1:0] ccxw7l8izxzjj14ozqkgvvyd6 =
                           {
                             ndsqg7zrec89ncrv9yu3k
                           } ;

  assign xzpsiztjmn62eb967x1xkc6 =
                           {
                             l_s_khzs83700pzjuq3_obo44
                           } ;

  assign a_dm6kd_qbw2cv84wtboltif01 =
                           {
                             tcrjx_8vlmtrlqjvk3tu
                           } ;

  assign ae00o9ay050qc5d5zxf18282b92 =
                           {
                             y0jaju01t8mqh2ycz05limpxfu
                           } ;

  assign puxr8jzij0m30qcwmdz2sufl51 =
                           {
                             x88dy7qz1z117o2jmbslutlpm
                           } ;
                         
  assign s6vj39lt1yt7f1ytk3pr3 =
                           {
                             kykdx6vx9n3hm7k6oybv
                           } ;

  assign wspjbjcpf459zy17qhyz8jmqy7 =
                           {
                             b59iokn7e2645ocyqifdk6sp1
                           } ;
                           
  assign y7jg1o7n3jl52fxr0isdv8 =
                           {
                             xs2l1_f3yynnrl_rw2zbe
                           } ;

  assign w8o2oxw46tp1zf4rujrx4zyxw =
                           {
                             wd3zc6palghmam9to3v2
                           } ;


  assign                   {
                             zw6mbnvv_8hcztypnytp87v_vy
                           } = w0hjg2xow0ymilw7bcxpm2l;

  
  assign                   {
                             hf8rqlrzsk0e9ho4orde_r
                           } = qkiytqsa_fo9x5ls7yb_x1k2;

  assign                   {
                             hng3_y3ldjtyu4a9n45
                           } = wzmdtyq65i82w_tt0juwqle;

  assign                   {
                             y1ovf4ea_l0kgs84_pwk6czrs
                           } = kz10yoaxkacgm38dwv37tl2ixfv;
                           
  assign                   {
                             n6fa00b9i708mtqu7yc9wjvxip
                           } = fyvkbec2dn4rlcslyiyttfrx;

  assign idw2i93am7m9wy_5hzipgymj5k3 = {
                             opns8_xijy8grr0gygeszh
                           };


  ux607_gnrl_icb_arbt # (
  .ALLOW_BURST (0),
  .ARBT_SCHEME (3),
  .FIFO_CUT_READY  (0),
  .ALLOW_0CYCL_RSP (0),
                       
  .FIFO_OUTS_NUM   (8),
  .ARBT_NUM   (tjt5wdq_mmk),
  .ARBT_PTR_W (vqmyiw_o188k),
  .USR_W      (s3xvyho),
  .AW         (16),
  .DW         (64) 
  ) zdem0krmjsk2wo(
  .arbt_active            (byiw0kxjclrie9tn3h),

  .o_icb_cmd_valid        (rqf8b5xxbw0n1_qaw )     ,
  .o_icb_cmd_ready        (ocwcf75wgxfb1bawe )     ,
  .o_icb_cmd_read         (gy2sgn_1bpkac7msq3 )      ,
  .o_icb_cmd_addr         (holgl43_yucp7f7l )      ,
  .o_icb_cmd_size         (wt4e4tlh0u_4cljr2j5f9)     ,
  .o_icb_cmd_wdata        (r_1u6q2lzkfus3o9nfl )     ,
  .o_icb_cmd_wmask        (yff7wf8wth2vjkdjpr)      ,
  .o_icb_cmd_burst        ()     ,
  .o_icb_cmd_beat         ()     ,
  .o_icb_cmd_excl         ()     ,
  .o_icb_cmd_lock         ()     ,
  .o_icb_cmd_usr          (syd0rz5l9shsemv)     ,
                           
  .o_icb_rsp_valid        (o4wuryrcvw13y2v5m6b6u )     ,
  .o_icb_rsp_ready        (bt4howrm5xnf6u4fuwrum6)     ,
  .o_icb_rsp_err          (vnqegbzme0jutvf)        ,
  .o_icb_rsp_excl_ok      (jdj122rbumyogtin6xpg97)    ,
  .o_icb_rsp_rdata        (p9mcc6npaw32uigcp6 )     ,
  .o_icb_rsp_usr          ({s3xvyho{1'b0}}  )     ,
                               
  .i_bus_icb_cmd_sel_vec  (ccxw7l8izxzjj14ozqkgvvyd6) ,

  .i_bus_icb_cmd_ready    (w0hjg2xow0ymilw7bcxpm2l ) ,
  .i_bus_icb_cmd_valid    (k1_j5ubhqqpfrl3p0bi186va9 ) ,
  .i_bus_icb_cmd_read     (a_dm6kd_qbw2cv84wtboltif01 )  ,
  .i_bus_icb_cmd_addr     (xzpsiztjmn62eb967x1xkc6 )  ,
  .i_bus_icb_cmd_wdata    (ae00o9ay050qc5d5zxf18282b92 ) ,
  .i_bus_icb_cmd_wmask    (puxr8jzij0m30qcwmdz2sufl51)  ,
  .i_bus_icb_cmd_burst    ({tjt5wdq_mmk{3'b0}}),
  .i_bus_icb_cmd_beat     ({tjt5wdq_mmk{2'b0}}),
  .i_bus_icb_cmd_excl     (wspjbjcpf459zy17qhyz8jmqy7 ),
  .i_bus_icb_cmd_lock     (s6vj39lt1yt7f1ytk3pr3 ),
  .i_bus_icb_cmd_size     (y7jg1o7n3jl52fxr0isdv8 ),
  .i_bus_icb_cmd_usr      (w8o2oxw46tp1zf4rujrx4zyxw ),
                                
  .i_bus_icb_rsp_valid    (qkiytqsa_fo9x5ls7yb_x1k2 ) ,
  .i_bus_icb_rsp_ready    (idw2i93am7m9wy_5hzipgymj5k3 ) ,
  .i_bus_icb_rsp_err      (wzmdtyq65i82w_tt0juwqle)    ,
  .i_bus_icb_rsp_excl_ok  (kz10yoaxkacgm38dwv37tl2ixfv),
  .i_bus_icb_rsp_rdata    (fyvkbec2dn4rlcslyiyttfrx ) ,
  .i_bus_icb_rsp_usr      () ,
                             
  .clk                    (gf33atgy  )                     ,
  .rst_n                  (ru_wi)
  );



endmodule

























module ad3c301j_tm48vb7x3
 #(
    parameter nm_fj = 32,
    parameter onr7l = 32, 
    parameter h1b = 4, 
    parameter ktra3i = 2,
    parameter rm39njpb7w = 16,
    parameter wvmre88 = 32, 
    parameter bf0ngee0t = 1, 
    parameter xbpsp4_i = 4, 
    parameter k2qm7hpa_qinpd = 7,
    parameter quofpn_rylwqbg9 = 1
    )
  (
  output vlb2az38tbnj4,
  
  
      
  input  ujj9wb8hyzso,
  

  
  
  
  input                          eth8quxx9hhjhxr4u9k2s77f,
  output                         zw6mbnvv_8hcztypnytp87v_vy,
  input  [nm_fj-1:0]                l_s_khzs83700pzjuq3_obo44,
  input                          tcrjx_8vlmtrlqjvk3tu, 
  input  [onr7l-1:0]                y0jaju01t8mqh2ycz05limpxfu, 
  input  [h1b-1:0]                x88dy7qz1z117o2jmbslutlpm, 
  input  [2-1:0]                 xs2l1_f3yynnrl_rw2zbe, 
  input                          kyvscpwy0vljnwysfxqxb,
  input                          sl5cpfvi658e8pl6nh2cm4,
  input                          tmqgi_fx924f3bq8ms4u8t0,

  output                         hf8rqlrzsk0e9ho4orde_r, 
  input                          opns8_xijy8grr0gygeszh, 
  output                         hng3_y3ldjtyu4a9n45,   
  output [onr7l-1:0]                n6fa00b9i708mtqu7yc9wjvxip, 
  output                         y1ovf4ea_l0kgs84_pwk6czrs,

   

  output [bf0ngee0t-1:0] d53gmmeaj,  
  output [rm39njpb7w-1:0] coouz2jyj2n, 
  output [xbpsp4_i-1:0] dcmn368x8,
  output [wvmre88-1:0] opsl7g4,          
  input  [wvmre88-1:0] tn65z3ytg,
  output              wzor2kya,

  


  input  gc4b3kdcan6do88ta_,
  input  gf33atgy,
  input  ru_wi
  );




  wire aht5xalx865dt9ymg6t4;
  wire zjmbnwsbyle24ayly67;
  wire [nm_fj-1:0]   icfwo5l56zab795f;
  wire n78yvkhg0miifi58; 
  wire [onr7l-1:0] wu02k99r_ok2kjj4u119us; 
  wire [h1b-1:0] ccwk4o03vlem_hqcccf1g6; 
  wire [2-1:0] ltx9lurd9p2ivmnufrgrw; 
  wire z6ncd60zcel8m99zg6v;
  wire st9_is6howar7iysonyyhk;
  wire o8407eu9fhzcuymr2a4;

  wire s4dz24kz7cxir4hxtt; 
  wire epoc75xqnuvcqziu_9i55h; 
  wire w0vagcfu1v7wkym9f;   
  wire [onr7l-1:0] gxo5tf4bea2gsq4yyn; 
  wire sjx2nupt4_7eb6_metse;



  
  assign aht5xalx865dt9ymg6t4 = eth8quxx9hhjhxr4u9k2s77f;
  assign zw6mbnvv_8hcztypnytp87v_vy = zjmbnwsbyle24ayly67; 

  assign icfwo5l56zab795f   = l_s_khzs83700pzjuq3_obo44  ;
  assign n78yvkhg0miifi58   = tcrjx_8vlmtrlqjvk3tu  ;   
  assign wu02k99r_ok2kjj4u119us  = y0jaju01t8mqh2ycz05limpxfu ;   
  assign ccwk4o03vlem_hqcccf1g6  = x88dy7qz1z117o2jmbslutlpm ;   
  assign ltx9lurd9p2ivmnufrgrw   = xs2l1_f3yynnrl_rw2zbe  ;   
  assign z6ncd60zcel8m99zg6v  = kyvscpwy0vljnwysfxqxb ;   
  assign st9_is6howar7iysonyyhk  = sl5cpfvi658e8pl6nh2cm4 ;   
  assign o8407eu9fhzcuymr2a4  = tmqgi_fx924f3bq8ms4u8t0 ;   

  
  assign hf8rqlrzsk0e9ho4orde_r   = s4dz24kz7cxir4hxtt  ; 
  assign epoc75xqnuvcqziu_9i55h   = opns8_xijy8grr0gygeszh  ;
  assign hng3_y3ldjtyu4a9n45     = w0vagcfu1v7wkym9f    ;
  assign y1ovf4ea_l0kgs84_pwk6czrs = sjx2nupt4_7eb6_metse;
  assign n6fa00b9i708mtqu7yc9wjvxip   = gxo5tf4bea2gsq4yyn  ;



  wire nbvps3m_gx6i5a5a0hv; 
  wire p4_qmsjuqyw_lnh1era6; 
  wire xiymrsmu7uxfwu75glhy;   
  wire [onr7l-1:0] e7spu5mj4_9vdij31ii; 
  wire kj9_2o6_25ucmc4g8v2gk_;


  
  wire [onr7l+2-1:0]ziubvvomv2nddezv;
  wire [onr7l+2-1:0]kgh1znd6ahvjhj;

  assign ziubvvomv2nddezv = {
                          kj9_2o6_25ucmc4g8v2gk_,
                          xiymrsmu7uxfwu75glhy,
                          e7spu5mj4_9vdij31ii
                          };

  assign {
                          sjx2nupt4_7eb6_metse,
                          w0vagcfu1v7wkym9f,
                          gxo5tf4bea2gsq4yyn
                          } = kgh1znd6ahvjhj;

  wire o_gjp7hu_0ltcb0f0liqo1og2ggf = s4dz24kz7cxir4hxtt & epoc75xqnuvcqziu_9i55h;
  ux607_gnrl_pipe_stage # (
   .CUT_READY(0),                                                                                                                  
   .DP(1),                                                                                                                         
   .DW(onr7l + 2)
  ) cndjid07t9lpndtd (
    .i_vld(nbvps3m_gx6i5a5a0hv),
    .i_rdy(p4_qmsjuqyw_lnh1era6),
    .i_dat(ziubvvomv2nddezv),
    .o_vld(s4dz24kz7cxir4hxtt),
    .o_rdy(epoc75xqnuvcqziu_9i55h),
    .o_dat(kgh1znd6ahvjhj),

    .clk(gf33atgy),
    .rst_n(ru_wi)
  );
  
  
  
  
  
  

  
  

  
  
  
  
  
  







  vfqtyk384n562k49kg #(
      .l9r6r   (bf0ngee0t),
      .w4mvurd (0),
      .onr7l     (onr7l),
      .nm_fj     (nm_fj),
      .h1b     (h1b),
      .ktra3i (ktra3i)
  ) hr5w2qfg8xstcjpmp0f(
     .ujj9wb8hyzso       (ujj9wb8hyzso),
     
     .v9ov1b3vn5k4ctkb (aht5xalx865dt9ymg6t4),
     .ub9pjiu4juf6nuqoq2w6 (zjmbnwsbyle24ayly67),
     .ogvavqa7ta836s  (n78yvkhg0miifi58 ),
     .aw0a19a967dn7n0x25w  (icfwo5l56zab795f ), 
     .leieaos4fnc5s_81kr  (ltx9lurd9p2ivmnufrgrw ), 
     .ty6a2k41y0e9ir8_yzg (z6ncd60zcel8m99zg6v ),
     .s4_gwe0uskrbhp37ksb (st9_is6howar7iysonyyhk ),
     .cwkq4r6_upg_2884r (o8407eu9fhzcuymr2a4 ),
     .air1drtzqvyz1ydvdej (1'b0),
     .ba79qari93k2d1309g (1'b0),
     .sc169gxpr38lpe8 (wu02k99r_ok2kjj4u119us), 
     .hg1g2yh6yktfe_btdst7 (ccwk4o03vlem_hqcccf1g6), 
  
     .dy9ll1o6t6ytby71hf4 (nbvps3m_gx6i5a5a0hv),
     .ow4hbh48f0mt6le4o (p4_qmsjuqyw_lnh1era6),
     .dek0xt7q6guk2vf6 (e7spu5mj4_9vdij31ii),
     .uzwj715coelxmfqs   (xiymrsmu7uxfwu75glhy),
  
     .d53gmmeaj   (d53gmmeaj  ),  
     .coouz2jyj2n (coouz2jyj2n), 
     .dcmn368x8  (dcmn368x8 ),
     .opsl7g4  (opsl7g4 ),          
     .tn65z3ytg (tn65z3ytg),
     .wzor2kya  (wzor2kya ),

  
  
     .gc4b3kdcan6do88ta_(gc4b3kdcan6do88ta_  ),
     .gf33atgy  (gf33atgy  ),
     .ru_wi(ru_wi)  
    );


  


  wire p4polvlxij557_ai;

  ux607_gnrl_icb_active # (
    .OUTS_CNT_W(4)
  ) uo66ekv3mrchnvmc03zw( 
      
      .icb_active    (p4polvlxij557_ai),

      .icb_cmd_valid (aht5xalx865dt9ymg6t4), 
      .icb_cmd_ready (zjmbnwsbyle24ayly67), 

      .icb_rsp_valid (nbvps3m_gx6i5a5a0hv), 
      .icb_rsp_ready (p4_qmsjuqyw_lnh1era6), 
    
      .clk           (gf33atgy  ),
      .rst_n         (ru_wi)
  );




  assign vlb2az38tbnj4 = p4polvlxij557_ai 
                    | o_gjp7hu_0ltcb0f0liqo1og2ggf 
;

  assign kj9_2o6_25ucmc4g8v2gk_ = 1'b0;

endmodule





















module trhtyw9g0vmmg56x(

  output                         gapxosc6nar47nfpz8,

  input                          bm7mey1b6dibd5i6lfpukeue,

  input                          a8h5u6ohzhowdrvqrnlllzd70h,
  output                         pz92yc3xo60c49ayrztvq18a,
  input  [16-1:0]   pwzrcrecvxehn8htjdn3kv2d0, 
  input                          m5itqssum7ljklhpn5nvzvd93, 
  input  [64-1:0]        kkk0rwd1njowzq01nvxke,
  input  [8-1:0]     a2kttuidwhopy02uoajaf,
  input                          g4hx0dbyp7f7ou8x02a0,
  input                          zce_icdtm3r9hzeanwhlu3fv,
  input  [1:0]                   jkp1oke9n1q9ikytwx_7k,
  input                          njyud2m27xz7r6j0g0ieq17m,
  input                          ksa323b46ngmxwazg70t76,
  input                          bs4xe3ath5_4_iwylkfwppp,
  
  output                         mu3ut_ezr05qz2bbi7_vc_aod,
  input                          sk3bm3yc69h4ac84pc4killh,
  output                         b7g_hkjxumf964flze01v6p  ,
  output                         cmtnwdaxz9zk1858kalga2vt,
  output [64-1:0]        qjvmrd1013dapqkahq_f87b,

  
  
  
  
  
  input                          c52ldkop361ts52m0,
  output                         x88wat37r_vjsn57a,
  input  [16-1:0]   z3k8ps_o7osj4uosf_6i5,
  input                          rzon56p292pybf35mi_,
  input                          jn_zyepkhmn_mdbqe1,
  input                          w8k_3fawz__hfg4mk0mw7g, 
  input                          i88maxesdvq1fkint66,
  input                          nao0kbyh1yex0kg7uycyc,
  
  output                         ult8a6a0b4agydwsws,
  output                         gkbxrtlrxlk7_fk4  ,
  output [64-1:0]        d27a6w261um4big8wy8,
  output                         bwdpzndejgg3liwep6q_,


  
  
  
  
  
  
  
  output                         tw0yf9aln_vu06k8l,
  input                          q84eo09gg53r2jj5a5xn,
  output [16-1:0]   ss4cm882613f24kdjqsyl,
  output                         oefdpb9h9kx627r_0y5,
  output                         zm9uosdggg7ntkh97elw,
  output                         g_ahl2zik6mj75atnp_hej,
  output                         bjl40q8m35dwdn_mn9, 
  output                         w15kr9553b0c7034t3, 
  output                         x3zbwtak7e2z5ecil, 
  output [64-1:0]        fh1jm1za5zvqmvdloi,
  output [8-1:0]     sp_0hv_ae5rrl9vagusi,
  output [1:0]                   ssswxj_bpfx_ebsbj,

  
  input                          fsj22rallxmhdrvuwenpq,
  input                          hhlfu4md9k5v7naf1qt  ,
  input  [64-1:0]        aapsfpke41r7dyya4ah,
  input                          klw_a8tw9atjooozntm,
  output                         yign8d_dhrow0i5wjts4bd,

  input  gf33atgy,
  input  ru_wi
  );

  localparam mz57rd1hv60923ped3d63 = 1
            ;

  localparam egb08sh4q_5pj = 1;

  localparam msjfsjsyuq0_ = (egb08sh4q_5pj + 1);	  


  localparam xbyxn4rc3zjgf7rj3 = msjfsjsyuq0_;	  

  localparam tjt5wdq_mmk = xbyxn4rc3zjgf7rj3;

  localparam vqmyiw_o188k = 2;
  
  localparam s3xvyho = 5;
  localparam y61y499cunmtec  = 0;
  localparam a69a9ho1_kmpwc58n  = 1;
  localparam zxf2f6zwhhxrms0dvq1  = 2;
  localparam e4ffeu06r85bh8f1  = 3;
  localparam qn77zdua2lv05_  = 4;
  wire                         x0i6aykuzxn1t7_hyw9s7r4to;
  wire                         pbyudse8quydhisrzo9pbl4;
  wire [16-1:0]   vapgj050raiah87lnzt_a; 
  wire                         h3ja79v9nz27634fb0t1v0; 
  wire [64-1:0]        pan4gqh4n90vt5ya5374l;
  wire [8-1:0]     li0xl_bt9ldz9ytg3epkvvia;
  wire                         y7jy10ammgs97wz327hiqd60;
  wire                         pov96j_pauowws9r0r61pft;
  wire [1:0]                   crye2awvchg9tzjetea_;
  wire                         cvksl3f95u8b10a3rmr6qvom; 
  wire                         togorwkvhfveb6zwndvww; 
  wire                         i036i6j05gm5ht39aak7k; 
  wire                         xubhke6y45gk7d9bj7c1022icq;
 
  wire                         c8u60qjfyfel53grl6lmf5_3;
  wire                         jrzlu53zewh6pdohs96buh;
  wire                         vhl77l_vrkmhgbq9nx8p8ix  ;
  wire [s3xvyho-1:0]             tp3slxhiijptdvp_mvj  ;
  wire                         g_44fovc09leckknqa3lf1skd;
  wire [64-1:0]        sedkfhar7baq5_wmvydzjmit2;


  wire [s3xvyho-1:0]             u4lxgrzm51v7wy57nf9xgk7n  ;
  
  

  assign x0i6aykuzxn1t7_hyw9s7r4to = c52ldkop361ts52m0;
  assign x88wat37r_vjsn57a = pbyudse8quydhisrzo9pbl4; 

  assign vapgj050raiah87lnzt_a  = z3k8ps_o7osj4uosf_6i5 ;
  assign cvksl3f95u8b10a3rmr6qvom = rzon56p292pybf35mi_;
  assign togorwkvhfveb6zwndvww = jn_zyepkhmn_mdbqe1;
  assign i036i6j05gm5ht39aak7k = w8k_3fawz__hfg4mk0mw7g; 
  assign xubhke6y45gk7d9bj7c1022icq = i88maxesdvq1fkint66; 
  
  assign h3ja79v9nz27634fb0t1v0   = 1'b1;
  assign pan4gqh4n90vt5ya5374l  = {64{1'b0}};
  assign li0xl_bt9ldz9ytg3epkvvia  = {8{1'b0}};
  assign y7jy10ammgs97wz327hiqd60   = 1'b0;
  assign pov96j_pauowws9r0r61pft   = 1'b0;
  assign crye2awvchg9tzjetea_   = 2'b11;

  
  assign ult8a6a0b4agydwsws   = c8u60qjfyfel53grl6lmf5_3  ; 
  assign jrzlu53zewh6pdohs96buh   = 1'b1  ;
  assign gkbxrtlrxlk7_fk4     = vhl77l_vrkmhgbq9nx8p8ix    ;
  assign d27a6w261um4big8wy8   = sedkfhar7baq5_wmvydzjmit2  ;
  assign {bwdpzndejgg3liwep6q_ 
                                } = tp3slxhiijptdvp_mvj[mz57rd1hv60923ped3d63-1:0];
  wire [s3xvyho-1:0] e4jwo8izi2p0lam = {
                                        {s3xvyho-mz57rd1hv60923ped3d63{1'b0}},
                                        klw_a8tw9atjooozntm
                                     };


  wire [s3xvyho-1:0] w83156lngsir086yhuvfdn_2;

  wire [s3xvyho-1:0] enz6_e8c8fa3hrmevg12ih1;


  wire [s3xvyho-1:0] gwtmxtc4wx3iu0ji;

  wire   ch1vt4b75lwy52i7at2exlbwhl = ~xubhke6y45gk7d9bj7c1022icq;
  assign w83156lngsir086yhuvfdn_2[y61y499cunmtec ] = i036i6j05gm5ht39aak7k;
  assign w83156lngsir086yhuvfdn_2[a69a9ho1_kmpwc58n ] = cvksl3f95u8b10a3rmr6qvom;
  assign w83156lngsir086yhuvfdn_2[qn77zdua2lv05_ ] = togorwkvhfveb6zwndvww;
  assign w83156lngsir086yhuvfdn_2[zxf2f6zwhhxrms0dvq1 ] = xubhke6y45gk7d9bj7c1022icq;
  assign w83156lngsir086yhuvfdn_2[e4ffeu06r85bh8f1 ] = ch1vt4b75lwy52i7at2exlbwhl;

  assign enz6_e8c8fa3hrmevg12ih1[y61y499cunmtec ] = njyud2m27xz7r6j0g0ieq17m;
  assign enz6_e8c8fa3hrmevg12ih1[a69a9ho1_kmpwc58n ] = ksa323b46ngmxwazg70t76;
  assign enz6_e8c8fa3hrmevg12ih1[qn77zdua2lv05_ ] = bs4xe3ath5_4_iwylkfwppp;
  assign enz6_e8c8fa3hrmevg12ih1[zxf2f6zwhhxrms0dvq1 ] = 1'b0;
  assign enz6_e8c8fa3hrmevg12ih1[e4ffeu06r85bh8f1 ] = 1'b0;
  

  assign bjl40q8m35dwdn_mn9 = gwtmxtc4wx3iu0ji[y61y499cunmtec ];
  assign zm9uosdggg7ntkh97elw = gwtmxtc4wx3iu0ji[a69a9ho1_kmpwc58n ];
  assign g_ahl2zik6mj75atnp_hej = gwtmxtc4wx3iu0ji[qn77zdua2lv05_ ];
  assign w15kr9553b0c7034t3 = gwtmxtc4wx3iu0ji[zxf2f6zwhhxrms0dvq1 ];
  assign x3zbwtak7e2z5ecil = gwtmxtc4wx3iu0ji[e4ffeu06r85bh8f1 ];


  wire [tjt5wdq_mmk*1-1:0] k1_j5ubhqqpfrl3p0bi186va9;
  wire [tjt5wdq_mmk*1-1:0] w0hjg2xow0ymilw7bcxpm2l;
  wire [tjt5wdq_mmk*16-1:0] xzpsiztjmn62eb967x1xkc6;
  wire [tjt5wdq_mmk*1-1:0] a_dm6kd_qbw2cv84wtboltif01;
  wire [tjt5wdq_mmk*64-1:0] ae00o9ay050qc5d5zxf18282b92;
  wire [tjt5wdq_mmk*8-1:0] puxr8jzij0m30qcwmdz2sufl51;
  wire [tjt5wdq_mmk*1-1:0] s6vj39lt1yt7f1ytk3pr3;
  wire [tjt5wdq_mmk*1-1:0] wspjbjcpf459zy17qhyz8jmqy7;
  wire [tjt5wdq_mmk*2-1:0] y7jg1o7n3jl52fxr0isdv8;
  wire [tjt5wdq_mmk*s3xvyho-1:0] w8o2oxw46tp1zf4rujrx4zyxw;

  wire [tjt5wdq_mmk*1-1:0] qkiytqsa_fo9x5ls7yb_x1k2;
  wire [tjt5wdq_mmk*1-1:0] idw2i93am7m9wy_5hzipgymj5k3;
  wire [tjt5wdq_mmk*1-1:0] wzmdtyq65i82w_tt0juwqle;
  wire [tjt5wdq_mmk*s3xvyho-1:0] od5a1yudx9bmyqpwleexh4h9;
  wire [tjt5wdq_mmk*1-1:0] kz10yoaxkacgm38dwv37tl2ixfv;
  wire [tjt5wdq_mmk*64-1:0] fyvkbec2dn4rlcslyiyttfrx;

  
  assign k1_j5ubhqqpfrl3p0bi186va9 =
      
                           {
                             x0i6aykuzxn1t7_hyw9s7r4to
							 , a8h5u6ohzhowdrvqrnlllzd70h

                           } ;

  wire[tjt5wdq_mmk-1:0] ccxw7l8izxzjj14ozqkgvvyd6 =
                           {
								  nao0kbyh1yex0kg7uycyc
                                  ,bm7mey1b6dibd5i6lfpukeue

                           } ;

  assign xzpsiztjmn62eb967x1xkc6 =
                           {
                             vapgj050raiah87lnzt_a
							 ,pwzrcrecvxehn8htjdn3kv2d0
                           } ;

  assign a_dm6kd_qbw2cv84wtboltif01 =
                           {
                             h3ja79v9nz27634fb0t1v0
							 , m5itqssum7ljklhpn5nvzvd93

                           } ;

  assign ae00o9ay050qc5d5zxf18282b92 =
                           {
                             pan4gqh4n90vt5ya5374l
							 , kkk0rwd1njowzq01nvxke

                           } ;

  assign puxr8jzij0m30qcwmdz2sufl51 =
                           {
                             li0xl_bt9ldz9ytg3epkvvia
							 ,a2kttuidwhopy02uoajaf

                           } ;
                         
  assign s6vj39lt1yt7f1ytk3pr3 =
                           {
                             y7jy10ammgs97wz327hiqd60
							 ,g4hx0dbyp7f7ou8x02a0

                           } ;

  assign wspjbjcpf459zy17qhyz8jmqy7 =
                           {
                             pov96j_pauowws9r0r61pft
							 ,zce_icdtm3r9hzeanwhlu3fv

                           } ;
                           
  assign y7jg1o7n3jl52fxr0isdv8 =
                           {
                             crye2awvchg9tzjetea_
							 ,
                             jkp1oke9n1q9ikytwx_7k

                           } ;

  assign w8o2oxw46tp1zf4rujrx4zyxw =
                           {
                             w83156lngsir086yhuvfdn_2
							 , enz6_e8c8fa3hrmevg12ih1

                           } ;


  assign                   {
                             pbyudse8quydhisrzo9pbl4
							 , pz92yc3xo60c49ayrztvq18a

                           } = w0hjg2xow0ymilw7bcxpm2l;

  
  assign                   {
                             c8u60qjfyfel53grl6lmf5_3
							 ,
                             mu3ut_ezr05qz2bbi7_vc_aod

                           } = qkiytqsa_fo9x5ls7yb_x1k2;

  assign                   {
                             vhl77l_vrkmhgbq9nx8p8ix
							 ,
                             b7g_hkjxumf964flze01v6p

                           } = wzmdtyq65i82w_tt0juwqle;

  assign                   {
                             tp3slxhiijptdvp_mvj
							 ,
                             u4lxgrzm51v7wy57nf9xgk7n

                           } = od5a1yudx9bmyqpwleexh4h9;
  assign                   {
                             g_44fovc09leckknqa3lf1skd
							 ,
                             cmtnwdaxz9zk1858kalga2vt

                           } = kz10yoaxkacgm38dwv37tl2ixfv;
                           
  assign                   {
                             sedkfhar7baq5_wmvydzjmit2
							 ,
                             qjvmrd1013dapqkahq_f87b

                           } = fyvkbec2dn4rlcslyiyttfrx;

  assign idw2i93am7m9wy_5hzipgymj5k3 = {
                             jrzlu53zewh6pdohs96buh
							 ,
                             sk3bm3yc69h4ac84pc4killh

                           };


  ux607_gnrl_icb_arbt # (
  .ALLOW_BURST (0),
  .ARBT_SCHEME (3),
  .FIFO_CUT_READY  (0),
  .ALLOW_0CYCL_RSP (0),
                       
  .FIFO_OUTS_NUM   (3),
  .ARBT_NUM   (tjt5wdq_mmk),
  .ARBT_PTR_W (vqmyiw_o188k),
  .USR_W      (s3xvyho),
  .AW         (16),
  .DW         (64) 
  ) kcq1dt918_wrdfr3v(
  .arbt_active            (gapxosc6nar47nfpz8),

  .o_icb_cmd_valid        (tw0yf9aln_vu06k8l )     ,
  .o_icb_cmd_ready        (q84eo09gg53r2jj5a5xn )     ,
  .o_icb_cmd_read         (oefdpb9h9kx627r_0y5 )      ,
  .o_icb_cmd_addr         (ss4cm882613f24kdjqsyl )      ,
  .o_icb_cmd_size         (ssswxj_bpfx_ebsbj)     ,
  .o_icb_cmd_wdata        (fh1jm1za5zvqmvdloi )     ,
  .o_icb_cmd_wmask        (sp_0hv_ae5rrl9vagusi)      ,
  .o_icb_cmd_burst        ()     ,
  .o_icb_cmd_beat         ()     ,
  .o_icb_cmd_excl         ()     ,
  .o_icb_cmd_lock         ()     ,
  .o_icb_cmd_usr          (gwtmxtc4wx3iu0ji)     ,
                           
  .o_icb_rsp_valid        (fsj22rallxmhdrvuwenpq )     ,
  .o_icb_rsp_ready        (yign8d_dhrow0i5wjts4bd)     ,
  .o_icb_rsp_err          (hhlfu4md9k5v7naf1qt)        ,
  .o_icb_rsp_excl_ok      (1'b0)    ,
  .o_icb_rsp_rdata        (aapsfpke41r7dyya4ah )     ,
  .o_icb_rsp_usr          (e4jwo8izi2p0lam)     ,
                               
  .i_bus_icb_cmd_sel_vec  (ccxw7l8izxzjj14ozqkgvvyd6) ,

  .i_bus_icb_cmd_ready    (w0hjg2xow0ymilw7bcxpm2l ) ,
  .i_bus_icb_cmd_valid    (k1_j5ubhqqpfrl3p0bi186va9 ) ,
  .i_bus_icb_cmd_read     (a_dm6kd_qbw2cv84wtboltif01 )  ,
  .i_bus_icb_cmd_addr     (xzpsiztjmn62eb967x1xkc6 )  ,
  .i_bus_icb_cmd_wdata    (ae00o9ay050qc5d5zxf18282b92 ) ,
  .i_bus_icb_cmd_wmask    (puxr8jzij0m30qcwmdz2sufl51)  ,
  .i_bus_icb_cmd_burst    ({tjt5wdq_mmk{3'b0}}),
  .i_bus_icb_cmd_beat     ({tjt5wdq_mmk{2'b0}}),
  .i_bus_icb_cmd_excl     (wspjbjcpf459zy17qhyz8jmqy7 ),
  .i_bus_icb_cmd_lock     (s6vj39lt1yt7f1ytk3pr3 ),
  .i_bus_icb_cmd_size     (y7jg1o7n3jl52fxr0isdv8 ),
  .i_bus_icb_cmd_usr      (w8o2oxw46tp1zf4rujrx4zyxw ),
                                
  .i_bus_icb_rsp_valid    (qkiytqsa_fo9x5ls7yb_x1k2 ) ,
  .i_bus_icb_rsp_ready    (idw2i93am7m9wy_5hzipgymj5k3 ) ,
  .i_bus_icb_rsp_err      (wzmdtyq65i82w_tt0juwqle)    ,
  .i_bus_icb_rsp_excl_ok  (kz10yoaxkacgm38dwv37tl2ixfv),
  .i_bus_icb_rsp_rdata    (fyvkbec2dn4rlcslyiyttfrx ) ,
  .i_bus_icb_rsp_usr      (od5a1yudx9bmyqpwleexh4h9 ) ,
                             
  .clk                    (gf33atgy  )                     ,
  .rst_n                  (ru_wi)
  );

endmodule

























module odg9yeykg220ymcco
 #(
    parameter nm_fj = 32,
    parameter onr7l = 32, 
    parameter h1b = 4, 
    parameter ktra3i =2,
    parameter rm39njpb7w = 16,
    parameter wvmre88 = 32, 
    parameter bf0ngee0t = 1, 
    parameter xbpsp4_i = 4, 
    parameter k2qm7hpa_qinpd = 7,
    parameter quofpn_rylwqbg9 = 1
    )
  (
  output qz0hhqemjh,
  
  
      
  input  ujj9wb8hyzso,
  
  
  input  ndsqg7zrec89ncrv9yu3k,

  input                          bm7mey1b6dibd5i6lfpukeue,

  input                          a8h5u6ohzhowdrvqrnlllzd70h,
  output                         pz92yc3xo60c49ayrztvq18a,
  input  [16-1:0]   pwzrcrecvxehn8htjdn3kv2d0, 
  input                          m5itqssum7ljklhpn5nvzvd93, 
  input  [64-1:0]        kkk0rwd1njowzq01nvxke,
  input  [8-1:0]     a2kttuidwhopy02uoajaf,
  input                          g4hx0dbyp7f7ou8x02a0,
  input                          zce_icdtm3r9hzeanwhlu3fv,
  input  [1:0]                   jkp1oke9n1q9ikytwx_7k,
  input                          njyud2m27xz7r6j0g0ieq17m,
  input                          ksa323b46ngmxwazg70t76,
  input                          bs4xe3ath5_4_iwylkfwppp,
  
  output                         mu3ut_ezr05qz2bbi7_vc_aod,
  input                          sk3bm3yc69h4ac84pc4killh,
  output                         b7g_hkjxumf964flze01v6p  ,
  output                         cmtnwdaxz9zk1858kalga2vt,
  output [64-1:0]        qjvmrd1013dapqkahq_f87b,
  
  
  
  
  
  
  
  input  c52ldkop361ts52m0,
  output x88wat37r_vjsn57a,
  input  [nm_fj-1:0] z3k8ps_o7osj4uosf_6i5,
  input  rzon56p292pybf35mi_,
  input  jn_zyepkhmn_mdbqe1,
  input  w8k_3fawz__hfg4mk0mw7g,
  input  i88maxesdvq1fkint66,
  input  nao0kbyh1yex0kg7uycyc,

  output ult8a6a0b4agydwsws, 
  output gkbxrtlrxlk7_fk4,   
  output [onr7l-1:0] d27a6w261um4big8wy8, 
  output bwdpzndejgg3liwep6q_, 
  

  output [bf0ngee0t-1:0] d53gmmeaj,  
  output [rm39njpb7w-1:0] coouz2jyj2n, 
  output [xbpsp4_i-1:0] dcmn368x8,
  output [wvmre88-1:0] opsl7g4,          
  input  [wvmre88-1:0] tn65z3ytg,
  output              wzor2kya,

  

  input [8*32-1:0] pcr4upio7_tx37, 
  input [8*1-1:0] uzklqlncpqqm1rav,
  input [8*1-1:0] ortueunvnkx_l5m_j,
  input [8*1-1:0] hwuhtb7ucto_utk56,
  input [8*2-1:0] i1env2kmns7qvvuuc,
  input [8*1-1:0] g3s3vpafvy3i,


  input  gc4b3kdcan6do88ta_,
  input  gf33atgy,
  input  ru_wi
  );

  localparam e5uali4u800wo_y_vg0 = 0;
  localparam ki03am94rna_vw1j = e5uali4u800wo_y_vg0;
  localparam xy2bbpcor078mpqxrm = ki03am94rna_vw1j; 
  localparam s3xvyho = xy2bbpcor078mpqxrm + 1;



  wire th06du2c8e2_b7k;
  wire irjoi8wvo25u209f_5;
  wire zxe59xihintdqfy9d;
  wire [nm_fj-1:0] zvk11dhgg2s67mkq;
  wire fbzs0o4ysyuzeg_qdj;
  wire me1n4pvwxa7n3u8l05;
  wire qaidts35dk5jcji0n;
  wire r8nzx6_1no31zeloft;
  wire vo0q_cm1x8dbf97fd;
  wire [onr7l-1:0] u4r4b_6kp09q767q;
  wire [h1b-1:0] lhibcc3xwm6cy;
  wire [2-1:0] r19ik0uppwcr;

  wire klkflmsyyf5w7ar; 
  wire wy36iirxspfw56864; 
  wire lkjqs6kiuyj;   
  wire [onr7l-1:0] h7f6k_ims_9p3; 
  wire sxxoah7zbvh8noti;

  wire zs89k7qgupd1xlvx63l2r; 
  wire iaaolhc_afh_9est07sqv; 
  wire u6w9b_jfa7l3hw7mrgi;   
  wire [onr7l-1:0] k2vp4nzypxpjqeoddj5a; 
  wire kbw6te9rg57czki5bi_qw;

  wire gapxosc6nar47nfpz8;

  trhtyw9g0vmmg56x r4kicw0ojal14fl(

     .gapxosc6nar47nfpz8(gapxosc6nar47nfpz8),

     .bm7mey1b6dibd5i6lfpukeue (bm7mey1b6dibd5i6lfpukeue),
     .a8h5u6ohzhowdrvqrnlllzd70h(a8h5u6ohzhowdrvqrnlllzd70h),
     .pz92yc3xo60c49ayrztvq18a(pz92yc3xo60c49ayrztvq18a),
     .pwzrcrecvxehn8htjdn3kv2d0 (pwzrcrecvxehn8htjdn3kv2d0 ), 
     .m5itqssum7ljklhpn5nvzvd93 (m5itqssum7ljklhpn5nvzvd93 ), 
     .kkk0rwd1njowzq01nvxke(kkk0rwd1njowzq01nvxke),
     .a2kttuidwhopy02uoajaf(a2kttuidwhopy02uoajaf),
     .g4hx0dbyp7f7ou8x02a0 (g4hx0dbyp7f7ou8x02a0 ),
     .zce_icdtm3r9hzeanwhlu3fv (zce_icdtm3r9hzeanwhlu3fv ),
     .jkp1oke9n1q9ikytwx_7k (jkp1oke9n1q9ikytwx_7k ),
     .njyud2m27xz7r6j0g0ieq17m (njyud2m27xz7r6j0g0ieq17m ),
     .ksa323b46ngmxwazg70t76 (ksa323b46ngmxwazg70t76 ),
     .bs4xe3ath5_4_iwylkfwppp (bs4xe3ath5_4_iwylkfwppp ),
     .mu3ut_ezr05qz2bbi7_vc_aod  (mu3ut_ezr05qz2bbi7_vc_aod  ),
     .sk3bm3yc69h4ac84pc4killh  (sk3bm3yc69h4ac84pc4killh  ),
     .b7g_hkjxumf964flze01v6p    (b7g_hkjxumf964flze01v6p    ),
     .cmtnwdaxz9zk1858kalga2vt(cmtnwdaxz9zk1858kalga2vt),
     .qjvmrd1013dapqkahq_f87b  (qjvmrd1013dapqkahq_f87b  ),

     .c52ldkop361ts52m0 (c52ldkop361ts52m0),
     .x88wat37r_vjsn57a (x88wat37r_vjsn57a),
     .z3k8ps_o7osj4uosf_6i5  (z3k8ps_o7osj4uosf_6i5 ),
     .rzon56p292pybf35mi_ (rzon56p292pybf35mi_),
     .jn_zyepkhmn_mdbqe1 (jn_zyepkhmn_mdbqe1),
     .w8k_3fawz__hfg4mk0mw7g (w8k_3fawz__hfg4mk0mw7g), 
     .i88maxesdvq1fkint66 (i88maxesdvq1fkint66),
	 .nao0kbyh1yex0kg7uycyc(nao0kbyh1yex0kg7uycyc),
                                          
     .ult8a6a0b4agydwsws (ult8a6a0b4agydwsws),
     .gkbxrtlrxlk7_fk4   (gkbxrtlrxlk7_fk4  ),
     .bwdpzndejgg3liwep6q_   (bwdpzndejgg3liwep6q_  ),
     .d27a6w261um4big8wy8 (d27a6w261um4big8wy8),


     .tw0yf9aln_vu06k8l (th06du2c8e2_b7k),
     .q84eo09gg53r2jj5a5xn (irjoi8wvo25u209f_5),
     .ss4cm882613f24kdjqsyl  (zvk11dhgg2s67mkq ),
     .oefdpb9h9kx627r_0y5  (zxe59xihintdqfy9d ),
     .zm9uosdggg7ntkh97elw (fbzs0o4ysyuzeg_qdj),
     .g_ahl2zik6mj75atnp_hej (me1n4pvwxa7n3u8l05),
     .bjl40q8m35dwdn_mn9 (qaidts35dk5jcji0n), 
     .w15kr9553b0c7034t3 (r8nzx6_1no31zeloft),
     .x3zbwtak7e2z5ecil (vo0q_cm1x8dbf97fd),
     .fh1jm1za5zvqmvdloi (u4r4b_6kp09q767q),
     .sp_0hv_ae5rrl9vagusi (lhibcc3xwm6cy),
     .ssswxj_bpfx_ebsbj  (r19ik0uppwcr ),
                                      
     .fsj22rallxmhdrvuwenpq (zs89k7qgupd1xlvx63l2r),
     .hhlfu4md9k5v7naf1qt   (u6w9b_jfa7l3hw7mrgi  ),
     .aapsfpke41r7dyya4ah (k2vp4nzypxpjqeoddj5a),
     .klw_a8tw9atjooozntm(kbw6te9rg57czki5bi_qw  ),
     .yign8d_dhrow0i5wjts4bd (iaaolhc_afh_9est07sqv),
     .gf33atgy  (gf33atgy  ),
     .ru_wi(ru_wi)  
  );





  wire v9ov1b3vn5k4ctkb;
  wire ub9pjiu4juf6nuqoq2w6;

  assign v9ov1b3vn5k4ctkb = th06du2c8e2_b7k;
  assign irjoi8wvo25u209f_5   = ub9pjiu4juf6nuqoq2w6;



  localparam csmadmx55manue7x3eepi = nm_fj + 4;
  wire [csmadmx55manue7x3eepi-1:0] uq8r9oikrd0fwx7;
  wire [csmadmx55manue7x3eepi-1:0] fqvk0uqonsuwykg8x;
  wire [nm_fj-1:0] v7q8td8d2htgx9l;
  wire ry6skqfxztdifqh4;
  wire zlxk8g_divsy1l;
  wire jtdssyaup2rfsui;
  wire oswjjcaw60mj0nu5;

  wire mil2qez5yypky6y3w97t = th06du2c8e2_b7k & irjoi8wvo25u209f_5;
  wire gkcxjf8pd9icfo9m; 
  wire k61r7muvzx7ha_fj3a = klkflmsyyf5w7ar & wy36iirxspfw56864;
  assign  uq8r9oikrd0fwx7 = {    zvk11dhgg2s67mkq
                               ,fbzs0o4ysyuzeg_qdj
                               ,qaidts35dk5jcji0n
                               ,r8nzx6_1no31zeloft
                               ,me1n4pvwxa7n3u8l05
                               };
  assign {  v7q8td8d2htgx9l
           ,ry6skqfxztdifqh4
           ,zlxk8g_divsy1l
           ,jtdssyaup2rfsui
           ,oswjjcaw60mj0nu5
           } = fqvk0uqonsuwykg8x;

  ux607_gnrl_fifo # (
   .CUT_READY(0),
   .MSKO(0),
   .DP(1),
   .DW(csmadmx55manue7x3eepi)
  ) t5jy7vqhrnq (
    .i_vld(mil2qez5yypky6y3w97t), 
    .i_rdy(),
    .i_dat(uq8r9oikrd0fwx7  ),
    .o_vld(gkcxjf8pd9icfo9m), 
    .o_rdy(k61r7muvzx7ha_fj3a), 
    .o_dat(fqvk0uqonsuwykg8x  ),
  
    .clk  (gf33atgy  ),
    .rst_n(ru_wi)  
   );

  localparam bfe8r_4hym5e4k = 32'h80000000;
  wire [32-1:0] eqvm7s0ujyq_yg4qw9e = {bfe8r_4hym5e4k[32-1:nm_fj], v7q8td8d2htgx9l};

  wire exot1hcpkxp3es = ~jtdssyaup2rfsui;
  wire c1rvv8xwiji7k = jtdssyaup2rfsui;
  wire ml9067zkhuig = 1'b0;
  wire qvjpb9kw9ae1dxuoz2tqwqp;
  
  assign sxxoah7zbvh8noti = qvjpb9kw9ae1dxuoz2tqwqp;

  d7stl61zflp21cls1tg kjnw8nf8sd_5ajjyn3x0 (
      .pcr4upio7_tx37     (pcr4upio7_tx37   ), 
      .uzklqlncpqqm1rav  (uzklqlncpqqm1rav),
      .ortueunvnkx_l5m_j  (ortueunvnkx_l5m_j),
      .hwuhtb7ucto_utk56  (hwuhtb7ucto_utk56),
      .i1env2kmns7qvvuuc  (i1env2kmns7qvvuuc),
      .g3s3vpafvy3i  (g3s3vpafvy3i),

      .sxvvsxtbhyvt    (1'b0),
      .rm1dxjejhq7dh3q5m  (1'b0 ),
      .xatytj_r0fv14q  (1'b0 ),

      .oily7    (c1rvv8xwiji7k),
      .ly3dor8    (ml9067zkhuig),
      .p1m    (exot1hcpkxp3es),

      .u2k4dyp52s_m(ry6skqfxztdifqh4),
      .bktu0z1mk56(zlxk8g_divsy1l),
      .e98zc_xde8d (eqvm7s0ujyq_yg4qw9e),
      .foj6m18  (qvjpb9kw9ae1dxuoz2tqwqp) 
  );

  



  vfqtyk384n562k49kg #(
      .l9r6r   (bf0ngee0t),
      .w4mvurd (1),
      .onr7l     (onr7l),
      .nm_fj     (nm_fj),
      .h1b     (h1b),
      .ktra3i (ktra3i)
  ) dg23xv64_tlt8qhf0f2d(
     .ujj9wb8hyzso       (ujj9wb8hyzso),
     
     .v9ov1b3vn5k4ctkb (v9ov1b3vn5k4ctkb),
     .ub9pjiu4juf6nuqoq2w6 (ub9pjiu4juf6nuqoq2w6),
     .ogvavqa7ta836s  (zxe59xihintdqfy9d ),
     .aw0a19a967dn7n0x25w  (zvk11dhgg2s67mkq ), 
     .leieaos4fnc5s_81kr  (r19ik0uppwcr ), 
     .ty6a2k41y0e9ir8_yzg (fbzs0o4ysyuzeg_qdj),
     .s4_gwe0uskrbhp37ksb (me1n4pvwxa7n3u8l05),
     .cwkq4r6_upg_2884r (qaidts35dk5jcji0n),
     .air1drtzqvyz1ydvdej (r8nzx6_1no31zeloft),
     .ba79qari93k2d1309g (vo0q_cm1x8dbf97fd),
     .sc169gxpr38lpe8 (u4r4b_6kp09q767q), 
     .hg1g2yh6yktfe_btdst7 (lhibcc3xwm6cy), 
  
     .dy9ll1o6t6ytby71hf4 (klkflmsyyf5w7ar),
     .ow4hbh48f0mt6le4o (wy36iirxspfw56864),
     .dek0xt7q6guk2vf6 (h7f6k_ims_9p3),
     .uzwj715coelxmfqs   (lkjqs6kiuyj),
  
     .d53gmmeaj   (d53gmmeaj  ),  
     .coouz2jyj2n (coouz2jyj2n), 
     .dcmn368x8  (dcmn368x8 ),
     .opsl7g4  (opsl7g4 ),          
     .tn65z3ytg (tn65z3ytg),
     .wzor2kya  (wzor2kya ),

  
  
     .gc4b3kdcan6do88ta_(gc4b3kdcan6do88ta_  ),
     .gf33atgy  (gf33atgy  ),
     .ru_wi(ru_wi)  
    );


  

  wire ygjpyr2srt2fpb7a;
  wire k0p07wax7i8qs4irfw = klkflmsyyf5w7ar;
  assign wy36iirxspfw56864 =  ygjpyr2srt2fpb7a;
  wire [s3xvyho-1:0] iwxu78sftoab_xrp = { sxxoah7zbvh8noti 
                                  };
  wire [64+s3xvyho:0] r194g36kplm5e5jwt = {
                                        h7f6k_ims_9p3
                                       ,lkjqs6kiuyj 
                                       ,iwxu78sftoab_xrp 
                                        };
  wire [64+s3xvyho:0] d7jq9fe2dpeqo396iig;
  assign {
            kbw6te9rg57czki5bi_qw
                          } = d7jq9fe2dpeqo396iig[s3xvyho-1:0]; 

  assign u6w9b_jfa7l3hw7mrgi = d7jq9fe2dpeqo396iig[s3xvyho]; 
  assign k2vp4nzypxpjqeoddj5a = d7jq9fe2dpeqo396iig[64+s3xvyho:s3xvyho+1]; 

  ux607_gnrl_pipe_stage # (
   .CUT_READY(0),                                                                                                                  
   .DP(1),                                                                                                                         
   .DW(64 + s3xvyho + 1)
  ) zulv5xxzsl9148lyi (
    .i_vld(k0p07wax7i8qs4irfw),
    .i_rdy(ygjpyr2srt2fpb7a),
    .i_dat(r194g36kplm5e5jwt),
    .o_vld(zs89k7qgupd1xlvx63l2r),
    .o_rdy(iaaolhc_afh_9est07sqv),
    .o_dat(d7jq9fe2dpeqo396iig),

    .clk(gf33atgy),
    .rst_n(ru_wi)
  );



  wire xi__l8hr5qqzazk;

  ux607_gnrl_icb_active # (
    .OUTS_CNT_W(3)
  ) enli1omqm5gvim( 
      
      .icb_active    (xi__l8hr5qqzazk),

      .icb_cmd_valid (v9ov1b3vn5k4ctkb), 
      .icb_cmd_ready (ub9pjiu4juf6nuqoq2w6), 

      .icb_rsp_valid (klkflmsyyf5w7ar), 
      .icb_rsp_ready (wy36iirxspfw56864), 
    
      .clk           (gf33atgy  ),
      .rst_n         (ru_wi)
  );


  assign qz0hhqemjh = xi__l8hr5qqzazk 
                    | gapxosc6nar47nfpz8
                    | zs89k7qgupd1xlvx63l2r
                    | gkcxjf8pd9icfo9m
                    ;


endmodule





















module vfqtyk384n562k49kg #(
    parameter w4mvurd = 0,
    parameter l9r6r = 1,
    parameter onr7l = 32,
    parameter h1b = 4,
    parameter nm_fj = 32,
    parameter ktra3i = 2 
)(
  
  
      
  input  ujj9wb8hyzso,
  
  
  
  
  input  v9ov1b3vn5k4ctkb, 
  output ub9pjiu4juf6nuqoq2w6, 
  input  ogvavqa7ta836s,  
  input  [nm_fj-1:0] aw0a19a967dn7n0x25w, 
  input  [onr7l-1:0] sc169gxpr38lpe8, 
  input  [h1b-1:0] hg1g2yh6yktfe_btdst7, 
  input  [2-1:0] leieaos4fnc5s_81kr, 
  input  ty6a2k41y0e9ir8_yzg,
  input  s4_gwe0uskrbhp37ksb,
  input  cwkq4r6_upg_2884r,
  input  air1drtzqvyz1ydvdej,
  input  ba79qari93k2d1309g,

  
  output dy9ll1o6t6ytby71hf4, 
  input  ow4hbh48f0mt6le4o, 
  output [onr7l-1:0] dek0xt7q6guk2vf6, 
  output uzwj715coelxmfqs, 

  output [l9r6r-1:0]      d53gmmeaj,  
  output [nm_fj-ktra3i-1:0] coouz2jyj2n, 
  output [h1b-1:0] dcmn368x8,
  output [onr7l-1:0] opsl7g4,          
  input  [onr7l-1:0] tn65z3ytg,
  output          wzor2kya,

  

  input  gc4b3kdcan6do88ta_,
  input  gf33atgy,
  input  ru_wi
  );
















































  
  
  
  

  ic0yi2sqfgf91w_hnsr #(
      .l9r6r   (l9r6r),
      .w4mvurd (w4mvurd),
      .onr7l     (onr7l),
      .nm_fj     (nm_fj),
      .h1b     (h1b),
      .ktra3i (ktra3i) 
  ) xo3ak26m3c1lfa5fb1g839x(
     .ujj9wb8hyzso       (ujj9wb8hyzso),
     
     
     
     
     
     
     
     
     
 
     .rknesgym0iijlr1u3v (v9ov1b3vn5k4ctkb),
     .vti6vqnpltrn64t39k (ub9pjiu4juf6nuqoq2w6),
     .z6n982dyua9x0eqp  (ogvavqa7ta836s ),
     .mddf4pbndy0oc4d4  (aw0a19a967dn7n0x25w ), 
     .u1ka1mgouppse (sc169gxpr38lpe8), 
     .nzj8jq9gceaf4a (hg1g2yh6yktfe_btdst7), 
     .mcipb0j9a8xv_j  (leieaos4fnc5s_81kr ),
     .e2kmvafoxxb7npnxu (ty6a2k41y0e9ir8_yzg),
     .ih2telexpjpi0ehern (s4_gwe0uskrbhp37ksb),
     .lea00ldnngihbv (cwkq4r6_upg_2884r),
     .x8ib2e59xcbcw (air1drtzqvyz1ydvdej),
     .pqqc8ir4ioesu (ba79qari93k2d1309g),

     .rjw47ts8n04ixvk (dy9ll1o6t6ytby71hf4),
     .t57z5g7wnk77b (ow4hbh48f0mt6le4o),
     .yome33f3f3s_p8j (dek0xt7q6guk2vf6),
     .mnzp2sek_cf9u   (uzwj715coelxmfqs  ),
  
     .d53gmmeaj   (d53gmmeaj  ),  
     .coouz2jyj2n (coouz2jyj2n), 
     .dcmn368x8  (dcmn368x8 ),
     .opsl7g4  (opsl7g4 ),          
     .tn65z3ytg (tn65z3ytg),
     .wzor2kya  (wzor2kya ),

  

     .gc4b3kdcan6do88ta_(gc4b3kdcan6do88ta_  ),
     .gf33atgy  (gf33atgy  ),
     .ru_wi(ru_wi)  
    );


endmodule









































module ic0yi2sqfgf91w_hnsr #(
    parameter w4mvurd = 0,
    parameter l9r6r = 1,
    parameter onr7l = 32,
    parameter h1b = 4,
    parameter nm_fj = 32,
    parameter ktra3i = 3 
)(
  
  
  
      
  input  ujj9wb8hyzso,
  
  
  
  
  input  rknesgym0iijlr1u3v, 
  output vti6vqnpltrn64t39k, 
  input  z6n982dyua9x0eqp,  
  input  [nm_fj-1:0] mddf4pbndy0oc4d4, 
  input  [onr7l-1:0] u1ka1mgouppse, 
  input  [h1b-1:0] nzj8jq9gceaf4a, 
  input  [1:0]    mcipb0j9a8xv_j,
  input  e2kmvafoxxb7npnxu,
  input  ih2telexpjpi0ehern,
  input  lea00ldnngihbv,
  input  x8ib2e59xcbcw,
  input  pqqc8ir4ioesu,

  
  output rjw47ts8n04ixvk, 
  input  t57z5g7wnk77b, 
  output [onr7l-1:0] yome33f3f3s_p8j, 
  output mnzp2sek_cf9u,

  output [l9r6r-1:0]      d53gmmeaj,  
  output [nm_fj-ktra3i-1:0] coouz2jyj2n, 
  output [h1b-1:0] dcmn368x8,
  output [onr7l-1:0] opsl7g4,          
  input  [onr7l-1:0] tn65z3ytg,
  output          wzor2kya,

  

  input  gc4b3kdcan6do88ta_,
  input  gf33atgy,
  input  ru_wi
  );


  ux607_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(1)
  ) vsmkuuhmv71me (
    .i_vld(rknesgym0iijlr1u3v), 
    .i_rdy(vti6vqnpltrn64t39k), 
    .i_dat(1'b0),
    .o_vld(rjw47ts8n04ixvk), 
    .o_rdy(t57z5g7wnk77b), 
    .o_dat(),
  
    .clk  (gf33atgy  ),
    .rst_n(ru_wi)  
   );
   generate
   if (l9r6r == 1) begin :spufqwrxip7qm
   assign d53gmmeaj = rknesgym0iijlr1u3v & vti6vqnpltrn64t39k;  
   end
   else begin :mk075oglayw
   assign d53gmmeaj[0] = rknesgym0iijlr1u3v && vti6vqnpltrn64t39k && ((&mcipb0j9a8xv_j) || !mddf4pbndy0oc4d4[ktra3i-1]);  
   assign d53gmmeaj[1] = rknesgym0iijlr1u3v && vti6vqnpltrn64t39k && ((&mcipb0j9a8xv_j) ||  mddf4pbndy0oc4d4[ktra3i-1]);  
   end
   endgenerate
   wire t2ziluu62w = (~z6n982dyua9x0eqp);  
   assign coouz2jyj2n= mddf4pbndy0oc4d4 [nm_fj-1:ktra3i];          
   assign dcmn368x8 = {h1b{t2ziluu62w}} & nzj8jq9gceaf4a[h1b-1:0];          
   assign opsl7g4 = u1ka1mgouppse[onr7l-1:0];          

   wire k12_lh2q7xhw = |d53gmmeaj | ujj9wb8hyzso;

   ux607_clkgate d_1aogp4xlh5z(
     .clk_in   (gf33atgy        ),
     .clkgate_bypass(gc4b3kdcan6do88ta_  ),
     .clock_en (k12_lh2q7xhw),
     .clk_out  (wzor2kya)
   );

   assign yome33f3f3s_p8j = tn65z3ytg;
   assign mnzp2sek_cf9u   = 1'b0;

   



endmodule




















module suzytsmnh3c_jk3y2hekvvubgi(
  input   vhqr9jgt5,

  input [6-1:0] u4amtcbhq_6g6rx9,
  input [5-1:0] sm0ktbr6as2sl7ho,

  output  rl_3d1m7gcc0,
  output  tsdapc3y0fh,
  output  mohep6fqp67x,
  output  mmmu7pm6e_uqx,

  output [8-1:0] e_9jhaby2__46fj,
  output [8-1:0] lpcj6ymxsst2n,
  output [8-1:0] wdb90nca460cp,
  output [8-1:0] rin3amuhzyhjgg 
);

  
  
  
  
  
  
  
  
  
  
  
  wire xjgw_pgn3zvvj81kjr = (sm0ktbr6as2sl7ho[3] == 1'b0);
  wire xcs9mpv5oxv3cqcwp63 = (sm0ktbr6as2sl7ho[3] == 1'b0);
  wire rissmhpk44xeppv2nnb = (sm0ktbr6as2sl7ho[3] == 1'b1);
  wire swmawuezj2sw5zqm = (sm0ktbr6as2sl7ho[3] == 1'b1);

  
  assign rl_3d1m7gcc0 = vhqr9jgt5;
  assign tsdapc3y0fh = vhqr9jgt5;
  assign mohep6fqp67x = vhqr9jgt5;
  assign mmmu7pm6e_uqx = vhqr9jgt5;

  wire hg7uzxj8k2t = xjgw_pgn3zvvj81kjr;
  wire tznbcmcotat8_j5 = xcs9mpv5oxv3cqcwp63;
  wire em0_90yhe07 = rissmhpk44xeppv2nnb;
  wire xe614yrxpmu = swmawuezj2sw5zqm;

  
  assign e_9jhaby2__46fj = {u4amtcbhq_6g6rx9, sm0ktbr6as2sl7ho[5-1:4], ~hg7uzxj8k2t};
  assign lpcj6ymxsst2n = {u4amtcbhq_6g6rx9, sm0ktbr6as2sl7ho[5-1:4], ~tznbcmcotat8_j5};
  assign wdb90nca460cp = {u4amtcbhq_6g6rx9, sm0ktbr6as2sl7ho[5-1:4], ~em0_90yhe07};
  assign rin3amuhzyhjgg = {u4amtcbhq_6g6rx9, sm0ktbr6as2sl7ho[5-1:4], ~xe614yrxpmu};

endmodule

module uy3gep77czajwdyrmq3ed7su(
  input   s71tjwwz,
  input   vhqr9jgt5,
  input [64-1:0] mm89bcd_zxeoe1y,
  input [8-1:0] amz4453y8nx6q,

  input [6-1:0] u4amtcbhq_6g6rx9,
  input [5-1:0] sm0ktbr6as2sl7ho,

  output  rl_3d1m7gcc0,
  output  tsdapc3y0fh,
  output  mohep6fqp67x,
  output  mmmu7pm6e_uqx,

  
  output [8-1:0] e_9jhaby2__46fj,
  output [8-1:0] lpcj6ymxsst2n,
  output [8-1:0] wdb90nca460cp,
  output [8-1:0] rin3amuhzyhjgg,
  
  output [32-1:0] e6rwnjewsq6s6oro,
  output [32-1:0] u74ed5k2tobo,
  output [32-1:0] cthiem_1bgmj,
  output [32-1:0] dg5w1zgjmlq1a4n,

  output [4-1:0] ft2vjq7oh7l1hzqu,
  output [4-1:0] wbr3gkcxil8f_hgq,
  output [4-1:0] t1ncj092lli,
  output [4-1:0] vhh7ujoe4fwn_8
);


  
  
  
  
  
  
  
  
  
  
  wire xjgw_pgn3zvvj81kjr = (sm0ktbr6as2sl7ho[3] == 1'b0);
  wire xcs9mpv5oxv3cqcwp63 = (sm0ktbr6as2sl7ho[3] == 1'b0);
  wire rissmhpk44xeppv2nnb = (sm0ktbr6as2sl7ho[3] == 1'b1);
  wire swmawuezj2sw5zqm = (sm0ktbr6as2sl7ho[3] == 1'b1);

  wire p7rmbur0xccjwdnk5 = (sm0ktbr6as2sl7ho[3] == 1'b1);
  wire ur1vxspyie29kpc = (sm0ktbr6as2sl7ho[3] == 1'b1);
  wire bslwrjopzc87oi4bsrv = (sm0ktbr6as2sl7ho[3] == 1'b0);
  wire go7d4ugf170bue27d = (sm0ktbr6as2sl7ho[3] == 1'b0);

  wire biipajw18_fl = s71tjwwz ? xjgw_pgn3zvvj81kjr : p7rmbur0xccjwdnk5; 
  wire jf_rufxm5ekxf = s71tjwwz ? xcs9mpv5oxv3cqcwp63 : ur1vxspyie29kpc;  
  wire yftvtx4ubo4h = s71tjwwz ? rissmhpk44xeppv2nnb : bslwrjopzc87oi4bsrv;  
  wire qqsaiabm1mheei = s71tjwwz ? swmawuezj2sw5zqm : go7d4ugf170bue27d; 

  assign rl_3d1m7gcc0 = vhqr9jgt5 & biipajw18_fl;
  assign tsdapc3y0fh = vhqr9jgt5 & jf_rufxm5ekxf; 
  assign mohep6fqp67x = vhqr9jgt5 & yftvtx4ubo4h; 
  assign mmmu7pm6e_uqx = vhqr9jgt5 & qqsaiabm1mheei;

  
  assign e_9jhaby2__46fj = {u4amtcbhq_6g6rx9, sm0ktbr6as2sl7ho[5-1:4], ~s71tjwwz};
  assign lpcj6ymxsst2n = {u4amtcbhq_6g6rx9, sm0ktbr6as2sl7ho[5-1:4], ~s71tjwwz};
  assign wdb90nca460cp = {u4amtcbhq_6g6rx9, sm0ktbr6as2sl7ho[5-1:4], ~s71tjwwz};
  assign rin3amuhzyhjgg = {u4amtcbhq_6g6rx9, sm0ktbr6as2sl7ho[5-1:4], ~s71tjwwz};

  assign e6rwnjewsq6s6oro = mm89bcd_zxeoe1y[31:00];
  assign u74ed5k2tobo = mm89bcd_zxeoe1y[63:32];
  assign cthiem_1bgmj = mm89bcd_zxeoe1y[31:00];
  assign dg5w1zgjmlq1a4n = mm89bcd_zxeoe1y[63:32];

  assign ft2vjq7oh7l1hzqu = amz4453y8nx6q[3:0];
  assign wbr3gkcxil8f_hgq = amz4453y8nx6q[7:4];
  assign t1ncj092lli = amz4453y8nx6q[3:0];
  assign vhh7ujoe4fwn_8 = amz4453y8nx6q[7:4];


endmodule

module y5gz1t0e4pyw9jr0abfow4_gfn1kng3(
  input   dpjdlj8bv4q,
  input   vhqr9jgt5,

  input [6-1:0] u4amtcbhq_6g6rx9,
  input [5-1:0] sm0ktbr6as2sl7ho,

  input  vpfe1f6au,
  input  g7u0q4_wwj_,

  input  [64-1:0] xduvlstjiiwj,
  input  [64-1:0] pbu6py7mm4i,

  output  rl_3d1m7gcc0,
  output  tsdapc3y0fh,
  output  mohep6fqp67x,
  output  mmmu7pm6e_uqx,

  output [32-1:0] e6rwnjewsq6s6oro,          
  output [32-1:0] u74ed5k2tobo,          
  output [32-1:0] cthiem_1bgmj,          
  output [32-1:0] dg5w1zgjmlq1a4n,          

  output [4-1:0] ft2vjq7oh7l1hzqu,          
  output [4-1:0] wbr3gkcxil8f_hgq,          
  output [4-1:0] t1ncj092lli,          
  output [4-1:0] vhh7ujoe4fwn_8,          

  output [8-1:0] e_9jhaby2__46fj,
  output [8-1:0] lpcj6ymxsst2n,
  output [8-1:0] wdb90nca460cp,
  output [8-1:0] rin3amuhzyhjgg
);

  
  
  
  
  
  
  
  

  
  assign rl_3d1m7gcc0 = vhqr9jgt5;
  assign tsdapc3y0fh = vhqr9jgt5; 
  assign mohep6fqp67x = vhqr9jgt5; 
  assign mmmu7pm6e_uqx = vhqr9jgt5; 

  wire tfxy7_r0ativro0 = vpfe1f6au;

  assign e_9jhaby2__46fj = {u4amtcbhq_6g6rx9, tfxy7_r0ativro0, ~dpjdlj8bv4q};
  assign lpcj6ymxsst2n = {u4amtcbhq_6g6rx9, tfxy7_r0ativro0, ~dpjdlj8bv4q};
  assign wdb90nca460cp = {u4amtcbhq_6g6rx9, tfxy7_r0ativro0, ~dpjdlj8bv4q};
  assign rin3amuhzyhjgg = {u4amtcbhq_6g6rx9, tfxy7_r0ativro0, ~dpjdlj8bv4q};


  
  assign e6rwnjewsq6s6oro = dpjdlj8bv4q ? xduvlstjiiwj[31:00] : pbu6py7mm4i[31:00] ;          
  assign u74ed5k2tobo = dpjdlj8bv4q ? xduvlstjiiwj[63:32] : pbu6py7mm4i[63:32] ;          
  assign cthiem_1bgmj = dpjdlj8bv4q ? pbu6py7mm4i[31:00] : xduvlstjiiwj[31:00] ;          
  assign dg5w1zgjmlq1a4n = dpjdlj8bv4q ? pbu6py7mm4i[63:32] : xduvlstjiiwj[63:32] ;          



  assign ft2vjq7oh7l1hzqu = g7u0q4_wwj_ ? {4{1'b1}} : {4{1'b0}};
  assign wbr3gkcxil8f_hgq = g7u0q4_wwj_ ? {4{1'b1}} : {4{1'b0}};
  assign t1ncj092lli = g7u0q4_wwj_ ? {4{1'b1}} : {4{1'b0}};
  assign vhh7ujoe4fwn_8 = g7u0q4_wwj_ ? {4{1'b1}} : {4{1'b0}};

endmodule

module p7k2hwgr9tazox9ivj695zpxhajkb(
  input   e5uheiss35t1,

  input [32-1:0] i6_p95sqjet02,          
  input [32-1:0] g8qh7ytfxpof4e_,          
  input [32-1:0] wt5ewwuq7uqf,          
  input [32-1:0] vxikm1a46oon,          

  output  [64-1:0] iw6t1cm4o67qw1,
  output  [64-1:0] mggrpeuiih45,
  output  [64-1:0] n9lrm5b8dl_r2gg,
  output  [64-1:0] xq_xgf70o0nt0zy 

);

  
  
  
  
  
  
  
  


  assign iw6t1cm4o67qw1 = e5uheiss35t1 ? {g8qh7ytfxpof4e_[31:0], i6_p95sqjet02[31:0]} : {vxikm1a46oon[31:0], wt5ewwuq7uqf[31:0]};
  assign mggrpeuiih45 = e5uheiss35t1 ? {vxikm1a46oon[31:0], wt5ewwuq7uqf[31:0]} : {g8qh7ytfxpof4e_[31:0], i6_p95sqjet02[31:0]};
  assign n9lrm5b8dl_r2gg = e5uheiss35t1 ? {g8qh7ytfxpof4e_[31:0], i6_p95sqjet02[31:0]} : {vxikm1a46oon[31:0], wt5ewwuq7uqf[31:0]}; 
  assign xq_xgf70o0nt0zy = e5uheiss35t1 ? {vxikm1a46oon[31:0], wt5ewwuq7uqf[31:0]} : {g8qh7ytfxpof4e_[31:0], i6_p95sqjet02[31:0]}; 



endmodule

module f2w7478x4kvdp7gsxub2tls31 #(
  parameter f16zrowg1s1f5 = 4,
  parameter mp26klefy4v2f = 4,
  parameter cu7ihzi5k8 = 4,
  parameter cqf2oxizzealhe = 1 
) (

  input  ffckqqivts0p,
  input  yseo05ez9cr0r,

  input  g5ptjmebcoo5nwcg,
  output pjmu7ih6ul43bacz,
  input  [f16zrowg1s1f5-1:0] s6tktwbreyy7r,
  input  h014w4n6dlj78fr3,
  input  jf6zw884wuj,

  output l1mjv4a3o1i7qxeru,
  input  vmc_730ubm6z6mit,
  output [mp26klefy4v2f-1:0] ok1b1b_3nv0,

  input  sgk1y63o9l50k3,
  output gqhewm9l9lvfgkbf7,
  input  [f16zrowg1s1f5-1:0] mchi632scfby1t0n,
  input  ofjszjvfai0r49q,
  input  mlewhkn_ph,

  output eapg2epq1a388t4,
  input  osuxnyc17r3xf,
  output [mp26klefy4v2f-1:0] sy8hpqbz5umprdog,

  output nk9dw9ied4zd2h,
  input  czec2uuagggq,
  output [f16zrowg1s1f5-1:0] d5xonxqryf7,

  input  qegs8svpsb6wzol,
  output k0csx0ynvoz54fjx,
  input  [mp26klefy4v2f-1:0] c20li_6i3x,

  output f5lbzfpsc02anbqy,

  input  gf33atgy,
  input  ru_wi
);

  wire ha_v037qx159m5 = nk9dw9ied4zd2h & czec2uuagggq;
  wire t572txr8fwwpm = qegs8svpsb6wzol & k0csx0ynvoz54fjx;

  wire ryk02bb42dwyksg;
  wire avdigyddrs6k4ffgtmr;
  wire n1aghvm5tz2vw1j0;
  wire gmdp1f22yjbki2pb;

  wire   ziu97huopy1h1whc = (~ryk02bb42dwyksg) & g5ptjmebcoo5nwcg;
  assign pjmu7ih6ul43bacz     = (~ryk02bb42dwyksg) & n1aghvm5tz2vw1j0;

  wire   ioul1ae6r946c3030 = (~avdigyddrs6k4ffgtmr) & sgk1y63o9l50k3;
  assign gqhewm9l9lvfgkbf7     = (~avdigyddrs6k4ffgtmr) & gmdp1f22yjbki2pb;

  wire qz2x37lhg63diy5fg1c6n = (yseo05ez9cr0r & 1'b1) | (ffckqqivts0p & 1'b0);
  wire e32w__6okfhy9dy = ryk02bb42dwyksg ? 1'b1 : avdigyddrs6k4ffgtmr ? 1'b0 : qz2x37lhg63diy5fg1c6n;

  wire sx9c860hj2s0m0ath;

  ux607_gnrl_fifo # (
   .CUT_READY(0),
   .DP(cu7ihzi5k8),
   .DW(cqf2oxizzealhe)
  ) jlqdbsky6gz6rpzbb8ps (
   .i_vld(ha_v037qx159m5),
   .i_rdy(sx9c860hj2s0m0ath), 
   .i_dat(e32w__6okfhy9dy),
   .o_vld(), 
   .o_rdy(t572txr8fwwpm), 
   .o_dat(f5lbzfpsc02anbqy),
 
   .clk  (gf33atgy  ),
   .rst_n(ru_wi)  
  );


  assign nk9dw9ied4zd2h  = (sx9c860hj2s0m0ath) & (ziu97huopy1h1whc | ioul1ae6r946c3030);
  assign n1aghvm5tz2vw1j0 = (sx9c860hj2s0m0ath) & czec2uuagggq & (~e32w__6okfhy9dy);
  assign gmdp1f22yjbki2pb = (sx9c860hj2s0m0ath) & czec2uuagggq & e32w__6okfhy9dy;

  assign d5xonxqryf7  = e32w__6okfhy9dy ? mchi632scfby1t0n  : s6tktwbreyy7r; 
  wire   s6ihn1xv9mba = e32w__6okfhy9dy ? ofjszjvfai0r49q : h014w4n6dlj78fr3; 
  wire   f_u78kx0t   = e32w__6okfhy9dy ? mlewhkn_ph   : jf6zw884wuj; 


  assign ok1b1b_3nv0 = c20li_6i3x;
  assign sy8hpqbz5umprdog = c20li_6i3x;
  assign k0csx0ynvoz54fjx = f5lbzfpsc02anbqy ? osuxnyc17r3xf : vmc_730ubm6z6mit; 
  assign l1mjv4a3o1i7qxeru = qegs8svpsb6wzol & (~f5lbzfpsc02anbqy);
  assign eapg2epq1a388t4 = qegs8svpsb6wzol &   f5lbzfpsc02anbqy ;

  
  
  wire ddvybufy77nvxthjk = (e32w__6okfhy9dy == 1'b1) & s6ihn1xv9mba & ha_v037qx159m5;
  
  wire sb3rvg4skymhquoxv = ryk02bb42dwyksg & f_u78kx0t & ha_v037qx159m5;
  wire zrlioy37cygj3_90z0a = ddvybufy77nvxthjk |   sb3rvg4skymhquoxv;
  wire pzzk1f38lzaxj5f17gw9qt = ddvybufy77nvxthjk & (~sb3rvg4skymhquoxv);
  
  ux607_gnrl_dfflr #(1) eo5fygmvyej8_swlydi5b (zrlioy37cygj3_90z0a, pzzk1f38lzaxj5f17gw9qt, ryk02bb42dwyksg, gf33atgy, ru_wi);

  
  
  wire w6nb6r3ciafkq6wph67 = (e32w__6okfhy9dy == 1'b0) & s6ihn1xv9mba & ha_v037qx159m5;
  
  wire ojnqigg33_6piae7ku50k = avdigyddrs6k4ffgtmr & f_u78kx0t & ha_v037qx159m5;
  wire zoyzrzgnbetmeb2qh4 = w6nb6r3ciafkq6wph67 |   ojnqigg33_6piae7ku50k;
  wire gud41sx2s2zj28zdl = w6nb6r3ciafkq6wph67 & (~ojnqigg33_6piae7ku50k);
  
  ux607_gnrl_dfflr #(1) u9nonitew587hemj32dj (zoyzrzgnbetmeb2qh4, gud41sx2s2zj28zdl, avdigyddrs6k4ffgtmr, gf33atgy, ru_wi);




endmodule


















module k7eqwfmolitp9my9g4(
  output zpdvh58o0evhzt,
  output q0duv6epk3ccff620vhhx2,
  output rpkosm9pbcpggwup90_ge9,
  output xwmkl_9n7oehwe7hh_a6aompojzukuik,
 
  output                               hv39pppvbmeqy8b6,
  input                                dukd0zozp1ektzmt7f,
  output[32-1:0]          t6l88yqbe4wokkhiso9t,
  output                               hyec__ebnw8lbcssd81,
  output                               vs2610q9_on1r996p,
  output                               coy3buxdw6yq3duh21azuwflk,
  output                               r_8h5lxb39ug57zli04e_o,
  output                               pv7q0ikpayogkay57rgyr,
  input                                dsq8f3rhmb7yc876v8,
  input                                enu_vumk17eoj1fma5ilz0,

  output                               ou74jmm5p6th0y0kcdwpqv2ey,
  output                               adwzzx09c_s_x1seh,
  input                                zp0aylmm0k4yw4w561bgzh,


  output kd96ha16hcj4wyo0,
  output j9kszxa35hle0cl9,
  output [6-1:0] myqlprv648_pqf92vvj,


  input  [32-1:0] z8alxhlwgz117, 
  input  [32-1:0] q4j831gvqooep12, 
  output tyg8z9t16af4e8xtdiw,
  output qkl9_olndwlohzaurunzkg,

  output                        fpihselr34pn79, 
  output                        jm4__y98e00ukvb4hiw_f, 

  input                         w4sit6hoc28giqb51t3n6,
  output                        tbli88os0gfvjlfl6ttv1,

  input  [32-1:0]  hxvldlso5zpp81, 
  input                         ahhi0t6w86wbz891shq, 
  input                         zkqavy8j9jzdikz_29v7am, 
  input                         ibt51xz_a6yo4yknr5mx1, 
  input  [64-1:0]       bl79n71wkynirgcs3,
  input  [8-1:0]    o8smcfmzt25hxpwcn,
  input                         y4tsxz4rprpynubw3rvm, 
  input                         n7jh1zclcr_s0l4bgd, 
  input                         wunjscg6om1d0yu8o, 
  input                         f24hbj6y6nq5sy45lqzm5s, 
  input                         od57enqth4m5g9lpdduxdx, 
  input                         vqfoysp81h8x_kvfv1sg56, 
  input                         l03z9wtep77xkwohwq0e_1lm, 
  input                         eymxkl1knoowfwizivwrzpsi, 
  input                         rbrj5qqhjrxh023fhy4v2ce, 
  input                         e4wqef4o71wrrp_crj0dw8, 
  input                         xdyys2soinatq_bm7r2g35ie, 

  output                        yp6atu2uzbb053onf7h7j_g3,
  output                        gl9dazcghkmei56i8tlb  ,
  output                        k7x2rdsdsxkmoiyluje7bf2aa  ,
  output[64-1:0]        j1utgrdwzlhqppb8rev5pbh55, 
 

  

  output                          rinamilgle00i5xmx_vt,
  input                           j8wlfupbw25hdmohz5q0,
  output  [32-1:0]   z64bwdr23steb7s9y9j, 
  output                          bg1spy6_v2kbo75pz1d6, 
  output  [64-1:0]        xyeq7c6icdac80_y0jup,
  output  [8-1:0]     za5ms2soyuucfxo_jbn,
  output  [2:0]                   b7aet1zp_fcfxn8h7rw0u1,
  output  [1:0]                   t3szwnvfo2nj3wk6r5kvt,
  output                          m4x1_gvw8v_sc8h7c8_6,
  output                          hpeqnhpztp9l_d3yx16l,
  output  [1:0]                   bngbyv57e7juc0vkk2y8i,
  output                          cneu8a119tg3vmie6zr2h_, 
  output                          jw2dzv9gi7gygudyqql6fz, 
  output                          o_7kpry6inkqpqi1bf1nd, 
  output                          f97tgz_qybmvln6nz5dqt458, 
  output                          znotwr53pu47f5m1agm, 

  output                          zf_v02okbs8_euhd64,
  input                           wq4r8m45isqp8_o4pdtitz,
  output  [32-1:0]   qpzo6lin6brrytho7, 
  output                          k7j6g0757jovg8xstgrvwf, 
  output  [64-1:0]      nwx86gohbrn08nvh60789,
  output  [8-1:0]      bebhplbk2k43sfoehvt66w,
  output  [2:0]                   ljk3q52m5tirt6shbcwbf,
  output  [1:0]                   ucj9poqgl683ej1pihkh,
  output                          u9hi0xtx8u0mn0l_7p,
  output                          rm04yhu6ondli9u0g6din,
  output  [1:0]                   o5fmtstd7kef7z4m7jefm,
  output                          vvadj6ew1h5wq9z5askkzr9, 
  output                          lop06h0_z_4tt1s04up, 
  output                          ivllgcn1kiix2iamzwf0u, 
  output                          rnmvpk356vfgxd_045g, 
  output                          a46c4xo4texvc9o, 
  
  
  
  input                           ze2bfnigu62i9937pcxnjc,
  output                          c86b14qr2qo45_qw2ns,
  input                           dm5b92mx0redfbuhs1u3d  ,
  input                           c4cb28s8l8rdx2e53vww,
  input [64-1:0]        c3vtv1izxu7rm5646jsmmke, 
  
  input                           mm70cenjp_1wmcs135nh4wl,
  output                          p4dpiqc4w_g42ni5jsaj,
  input                           ezntrtg3q1must0tfcgn  ,
  input                           h99vs7dtnw2w96vts56dhc2,
  input [64-1:0]        glqyhrpm6zzwddhsd6mcd1u, 

  output                          c9oejgc5s6_v8ooyy8c0x1, 
  output [64-1:0]    sktjnm1h7yu59cy6lnbf0gx40e_,  
  output                          izozgg91hphikoatw0xsa,  

  output                          m7rpuph0hm25ukmyralijiy, 
  output [64-1:0]    r_13gm13ck84al5d7ty5lf_m,  
  output                          ck7dirv94s9jkefjfed0h0mp,  
  
  

  output                          jkq984ky8fozrzq,
  output                          g3_8p4g7w5grnl62xy,
  input                           vqwqaofc8sz_yjccd,

  input                           tyxs3jzhr2i2gq9dt7,
  output                          zti98n829owa2p,
  input  [24-1:0]  ye256knohacnaakiw2nqck6,
  input  [24-1:0]  hyxeikuobvxjumz2hibay,
  input  [32-1:0]  zkojor8433oflab2kpvtzi1z9,
  input  [32-1:0]  nx6i4o0_cbqmlan1ylpodj9y,
  input  [32-1:0]  tgfv2w2s7qhwkl0pdpf_79v4e,
  input  [32-1:0]  qfjl6250hpfb57pxl0t53q6fd,
 
  
  output                          j2kcz1faqhvh1ler6j,  
  output [6-1:0]  a6gdkt5h77dh0mcj8t4gq,
  output                          wixbtbeqlhzelg4t ,
  output [24-1:0]  uh_ekyw7cw8c3d3xj1,          
   
  output                          uf44audysjgtvdnua67,  
  output [6-1:0]  qtcasxm90cy0bwaqaxz, 
  output                          y38seii6ja77q2jy08 ,
  output [24-1:0]  f42g8ulc2y43ntmai5,          

 


  input                            cgnsvvj7srbljqst,          
  
  
  output                          rgf8pa4kn20jusruz,  
  output [8-1:0] wjwjffxr_4lulivwz, 
  output [4-1:0] z6udkjbx164gh9yo1o,
  output [32-1:0] frkunk72hlttw0ar0np,          
                                  
  output                          r2tvaf8px0p9vlw4we,  
  output [8-1:0] srfn4smswwo6hbyaa, 
  output [4-1:0] a_u2kfmgv2ho357c,
  output [32-1:0] svj88sv2u56fepzmg,          
                                 
  output                          rzf167thmprvps0tm62i,  
  output [8-1:0] lv7fu0hif2n2zhmgtcc, 
  output [4-1:0] oj5t3f0lq1n9ae82x,
  output [32-1:0] hat38salswlktk821,          
                                
  output                          caxkrdjq0tjnnne9,  
  output [8-1:0] qpuk8ry0w9_r7ur4gcnx, 
  output [4-1:0] v8jl1eh8o0n5g765,
  output [32-1:0] c0xnu9p8he2hw10h,          

  input gf33atgy,
  input ru_wi
  );



     
  wire qhkxw_0dnntylavbxym4jh6kdq5;
  wire eq6xz7m5lnl9uvy2 = qhkxw_0dnntylavbxym4jh6kdq5 ? 1'b1 : (vqfoysp81h8x_kvfv1sg56 & l03z9wtep77xkwohwq0e_1lm);
  wire behhrrdejekhg_3v4ju = (vqfoysp81h8x_kvfv1sg56 & eymxkl1knoowfwizivwrzpsi);
  wire p2kqppuunqlu40r = (vqfoysp81h8x_kvfv1sg56 & rbrj5qqhjrxh023fhy4v2ce);
  wire ong4xrs8cubfol     = xdyys2soinatq_bm7r2g35ie;

  wire ldgy0gmteitowu43nw5 = (vqfoysp81h8x_kvfv1sg56 & eymxkl1knoowfwizivwrzpsi & (~l03z9wtep77xkwohwq0e_1lm));
  wire reffh2y56n2410r_6a54c  = eq6xz7m5lnl9uvy2 & e4wqef4o71wrrp_crj0dw8;
  wire lkkimoh3n0l0cploih  = behhrrdejekhg_3v4ju & e4wqef4o71wrrp_crj0dw8;

  wire s8iygpzng_5v9083x1skh1xq00434b6_ = vqfoysp81h8x_kvfv1sg56 & (~rbrj5qqhjrxh023fhy4v2ce);
  
  
  
  
  localparam rmrgua6tlcyvz6q9e  = 3;
  
  localparam x3l7iptxd_0o4qa66  = 3'd0;
  
  localparam upuj82vcjn7bivcb1q  = 3'd1;
  
  localparam vaakncgdsx0fhzn1  = 3'd2;
  
  localparam du5mug53rvo4exdqvb  = 3'd3;
  
  localparam g8al00jhg6lk0rm_54u  = 3'd4;
  
  localparam u4bfs29wpxrhgi2r  = 3'd5;
  
  localparam iq46j_jt063p5es7p  = 3'd6;
  
  localparam ozrbgq56cf8gpvw3  = 3'd7;
  
  wire [rmrgua6tlcyvz6q9e-1:0] uwn2_an5cnlum12v;
  wire [rmrgua6tlcyvz6q9e-1:0] i1doij84r9a3_;
  wire bm460sko0qpzmueg5;

  wire [rmrgua6tlcyvz6q9e-1:0] u99tnldu986760c5;
  wire [rmrgua6tlcyvz6q9e-1:0] htn58z08fvzcwm13x4z;
  wire [rmrgua6tlcyvz6q9e-1:0] nb3914w6z5nmnlsmou;
  wire [rmrgua6tlcyvz6q9e-1:0] ox24gqid_5st2md2nzm;
  wire [rmrgua6tlcyvz6q9e-1:0] s37i5yerdn69n2;
  wire [rmrgua6tlcyvz6q9e-1:0] y5ramxcxkrqsz12gk;
  wire [rmrgua6tlcyvz6q9e-1:0] f1o45m2wg79no44n5d;
  wire [rmrgua6tlcyvz6q9e-1:0] gyiivu76k6m_fi;
  wire wfoen161d4r42bkqp34lj;
  wire l_0ukthd8bmvihg5o40mjg2;
  wire ar7ss7g0h7o9d58_adekeyg;
  wire w326dccv5z3q6ww691lf;
  wire hayqsfattzuc50458bllmr;
  wire hln5byq3t_zxwy8c51dq;
  wire i1iwskvd2cedxy_x32z926u;
  wire j98f_s869qm5bv_dhgbcim3;


  
  wire m2nk0s7zuy2ivs6gx = (i1doij84r9a3_ == x3l7iptxd_0o4qa66);
  wire myiw_93cf76tua4vp2x = (i1doij84r9a3_ == upuj82vcjn7bivcb1q);
  wire hcnuxviddm5zvn0cyzv7m = (i1doij84r9a3_ == vaakncgdsx0fhzn1);
  wire g1evvi19a50ju8wyn5 = (i1doij84r9a3_ == du5mug53rvo4exdqvb);
  wire gjxds3mwzdpqkwxketiaa = (i1doij84r9a3_ == g8al00jhg6lk0rm_54u);
  wire mxk6xl0c64kzkrplmm = (i1doij84r9a3_ == u4bfs29wpxrhgi2r);
  wire uafmsty4hif2k4iobx = (i1doij84r9a3_ == iq46j_jt063p5es7p);
  wire r2dy3qdfqfohba22hlsf5 = (i1doij84r9a3_ == ozrbgq56cf8gpvw3);

  wire ue54sje856um8518nhjen;
  wire s9hgy6syn2arl9fxs8kb0;
  wire zqa26f3l044pht447ti8x_r8rmh;

      
          
  assign wfoen161d4r42bkqp34lj = m2nk0s7zuy2ivs6gx & ue54sje856um8518nhjen;
  assign u99tnldu986760c5      = upuj82vcjn7bivcb1q; 

          
  assign l_0ukthd8bmvihg5o40mjg2 = myiw_93cf76tua4vp2x & (hv39pppvbmeqy8b6 ? dukd0zozp1ektzmt7f : 1'b1);
  assign htn58z08fvzcwm13x4z      = 
                             (s8iygpzng_5v9083x1skh1xq00434b6_) ? (
                               
                                   du5mug53rvo4exdqvb
                         ) : vaakncgdsx0fhzn1;

      
          
  wire dkox2mp78q58i66;
  assign ar7ss7g0h7o9d58_adekeyg  = hcnuxviddm5zvn0cyzv7m & zqa26f3l044pht447ti8x_r8rmh ;
             
  assign nb3914w6z5nmnlsmou     = dkox2mp78q58i66 ? x3l7iptxd_0o4qa66 : du5mug53rvo4exdqvb; 
  
      
          
  wire imzw3o6xtgdmikumc;
  assign w326dccv5z3q6ww691lf  = g1evvi19a50ju8wyn5 & imzw3o6xtgdmikumc;
  assign ox24gqid_5st2md2nzm     = g8al00jhg6lk0rm_54u; 
  
      
          
  wire yhwk19tompbv5zx;
  assign hayqsfattzuc50458bllmr  = gjxds3mwzdpqkwxketiaa & yhwk19tompbv5zx;
  assign s37i5yerdn69n2     = u4bfs29wpxrhgi2r;
  
      
          
  wire o_0q4jefxhht9mcddirs7; 
  assign hln5byq3t_zxwy8c51dq  = mxk6xl0c64kzkrplmm & o_0q4jefxhht9mcddirs7;
  assign y5ramxcxkrqsz12gk     = iq46j_jt063p5es7p;
  
      
          
  wire jzytexqffyvv5d75cjxbqox8; 
  wire l88go20t1nggrq383;
  assign i1iwskvd2cedxy_x32z926u  = uafmsty4hif2k4iobx & jzytexqffyvv5d75cjxbqox8;
  assign f1o45m2wg79no44n5d     = l88go20t1nggrq383 ? ozrbgq56cf8gpvw3 : x3l7iptxd_0o4qa66; 
  
      
          
  wire zxz6ihlgme0sknfg8ncdly9z;
  assign j98f_s869qm5bv_dhgbcim3  = r2dy3qdfqfohba22hlsf5 & zxz6ihlgme0sknfg8ncdly9z ;
  assign gyiivu76k6m_fi     = x3l7iptxd_0o4qa66;
  

  
  assign bm460sko0qpzmueg5 = 
        wfoen161d4r42bkqp34lj |
        l_0ukthd8bmvihg5o40mjg2 |
        ar7ss7g0h7o9d58_adekeyg |
        w326dccv5z3q6ww691lf |
        hayqsfattzuc50458bllmr |
        hln5byq3t_zxwy8c51dq |
        i1iwskvd2cedxy_x32z926u |
        j98f_s869qm5bv_dhgbcim3;

  
  assign uwn2_an5cnlum12v = 
              ({rmrgua6tlcyvz6q9e{wfoen161d4r42bkqp34lj}} & u99tnldu986760c5)
            | ({rmrgua6tlcyvz6q9e{l_0ukthd8bmvihg5o40mjg2}} & htn58z08fvzcwm13x4z)
            | ({rmrgua6tlcyvz6q9e{ar7ss7g0h7o9d58_adekeyg}} & nb3914w6z5nmnlsmou)
            | ({rmrgua6tlcyvz6q9e{w326dccv5z3q6ww691lf}} & ox24gqid_5st2md2nzm)
            | ({rmrgua6tlcyvz6q9e{hayqsfattzuc50458bllmr}} & s37i5yerdn69n2)
            | ({rmrgua6tlcyvz6q9e{hln5byq3t_zxwy8c51dq}} & y5ramxcxkrqsz12gk)
            | ({rmrgua6tlcyvz6q9e{i1iwskvd2cedxy_x32z926u}} & f1o45m2wg79no44n5d)
            | ({rmrgua6tlcyvz6q9e{j98f_s869qm5bv_dhgbcim3}} & gyiivu76k6m_fi)
              ;

  ux607_gnrl_dfflr #(rmrgua6tlcyvz6q9e) zbc0vitfiyt3m9r3g (bm460sko0qpzmueg5, uwn2_an5cnlum12v, i1doij84r9a3_, gf33atgy, ru_wi);

  wire c2q6lda5ak6w6cr45iz_q4 = bm460sko0qpzmueg5 & (uwn2_an5cnlum12v == ozrbgq56cf8gpvw3); 
  wire tvalp2jhv5332aqhj12i = bm460sko0qpzmueg5 & (uwn2_an5cnlum12v == x3l7iptxd_0o4qa66); 

  assign jm4__y98e00ukvb4hiw_f = tvalp2jhv5332aqhj12i;


  assign fpihselr34pn79 = (~m2nk0s7zuy2ivs6gx); 
  assign tbli88os0gfvjlfl6ttv1 = m2nk0s7zuy2ivs6gx;




  wire rtfuf_qdpdfw3yf7b0xae = 1'b0
                           | dsq8f3rhmb7yc876v8
                           | enu_vumk17eoj1fma5ilz0
                           ;

  wire tt_8kztvw6mmh5kxjnrmef6dom = hv39pppvbmeqy8b6 & dukd0zozp1ektzmt7f & rtfuf_qdpdfw3yf7b0xae;
  wire mq15b0rzwjb5dc_b054jgqsk14s = jm4__y98e00ukvb4hiw_f;
  wire zpt2wiw4web6uqeqlyall52phd = tt_8kztvw6mmh5kxjnrmef6dom | mq15b0rzwjb5dc_b054jgqsk14s;
  wire l3smhdkp7na3d_o4i60mmnt_5kp = tt_8kztvw6mmh5kxjnrmef6dom;

  ux607_gnrl_dfflr #(1) u_kelrp2gw0aihdkcg_6jmir17wg (zpt2wiw4web6uqeqlyall52phd, l3smhdkp7na3d_o4i60mmnt_5kp, qhkxw_0dnntylavbxym4jh6kdq5, gf33atgy, ru_wi);

  assign hv39pppvbmeqy8b6  = myiw_93cf76tua4vp2x & ldgy0gmteitowu43nw5;
  assign t6l88yqbe4wokkhiso9t = hxvldlso5zpp81; 
  assign hyec__ebnw8lbcssd81 = 1'b0;
  assign vs2610q9_on1r996p= 1'b1;
  assign coy3buxdw6yq3duh21azuwflk = f24hbj6y6nq5sy45lqzm5s;
  assign r_8h5lxb39ug57zli04e_o = y4tsxz4rprpynubw3rvm;
  assign pv7q0ikpayogkay57rgyr = wunjscg6om1d0yu8o;

  assign ou74jmm5p6th0y0kcdwpqv2ey = 1'b0;
  assign adwzzx09c_s_x1seh = 1'b0;


  
  
  
  wire [3-1:0] o0td_p0x46d9jh72w4l1g4;
  wire [3-1:0] drjpx3qgvtravae6qzchne;
  wire d2i8ojpp6nmcemv = hayqsfattzuc50458bllmr;

  wire [3-1:0] pukmc1wrlg05lh7ua = ye256knohacnaakiw2nqck6[(24-1):21];
  wire [3-1:0] atzysb0ixj_b2ly3jzp = hyxeikuobvxjumz2hibay[(24-1):21];

  ux607_gnrl_dfflr #(3) eq42v57ewfzt5op (d2i8ojpp6nmcemv, pukmc1wrlg05lh7ua, o0td_p0x46d9jh72w4l1g4, gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(3) dl0k9v__dd7bn (d2i8ojpp6nmcemv, atzysb0ixj_b2ly3jzp, drjpx3qgvtravae6qzchne, gf33atgy, ru_wi);

  wire x7jix80161slp;
  ux607_gnrl_dfflr #(1) uk0h39gxuqwobgah_ (d2i8ojpp6nmcemv, cgnsvvj7srbljqst, x7jix80161slp, gf33atgy, ru_wi);


  wire tg3c0ha5844xz = o0td_p0x46d9jh72w4l1g4[0] & o0td_p0x46d9jh72w4l1g4[1] ;
  wire dvn3st2c0wavqa6 = drjpx3qgvtravae6qzchne[0] & drjpx3qgvtravae6qzchne[1] ;

  wire e0ny5yl0v2ik890te  = o0td_p0x46d9jh72w4l1g4[0] & o0td_p0x46d9jh72w4l1g4[2];
  wire uhrfddgw6k1clj2oc  = drjpx3qgvtravae6qzchne[0] & drjpx3qgvtravae6qzchne[2];

  
  
  
  
  wire tqiycgs52p5ubxsuyib_v1zt7;
      
           
           
  wire xb8j0rrc_88sw9m1_7ximu1sj = l_0ukthd8bmvihg5o40mjg2 & (~eq6xz7m5lnl9uvy2) & (~behhrrdejekhg_3v4ju);
      
  wire jxpj6_9tx5iktrgs;
  wire ydasmvx5h2ezeqd8nzjocww = tqiycgs52p5ubxsuyib_v1zt7 & jxpj6_9tx5iktrgs;
  wire u27qjkb5zqe12szsltsn84e = xb8j0rrc_88sw9m1_7ximu1sj |   ydasmvx5h2ezeqd8nzjocww;
  wire oy67t8p1b1as7_r4qp4hek3jt = (~ydasmvx5h2ezeqd8nzjocww);
  ux607_gnrl_dfflr #(1) v3tueeign88vdxdo7qvw12ytrgj (u27qjkb5zqe12szsltsn84e, oy67t8p1b1as7_r4qp4hek3jt, tqiycgs52p5ubxsuyib_v1zt7, gf33atgy, ru_wi);

  assign  rinamilgle00i5xmx_vt = tqiycgs52p5ubxsuyib_v1zt7; 

  assign s9hgy6syn2arl9fxs8kb0 = rinamilgle00i5xmx_vt & j8wlfupbw25hdmohz5q0;
  assign ue54sje856um8518nhjen = w4sit6hoc28giqb51t3n6 & tbli88os0gfvjlfl6ttv1;

  
  
  localparam ku4rkdvsjrgvr70b8i1e7dj7t7qedj = (4-1);
  
  wire [2-1:0] kwbmlmwj_ec;
    
  wire d2jsegrkoa154kuy = s9hgy6syn2arl9fxs8kb0;
    
  wire bxc0qc1hr_cb1a4x1zadth = (kwbmlmwj_ec == 2'b0);
  wire nlfdn3rz3118m7vvwo = (kwbmlmwj_ec == ku4rkdvsjrgvr70b8i1e7dj7t7qedj[2-1:0]);
  assign jxpj6_9tx5iktrgs = s9hgy6syn2arl9fxs8kb0 & nlfdn3rz3118m7vvwo;
  wire v0t2k69nbehh = d2jsegrkoa154kuy | jxpj6_9tx5iktrgs;
  wire [2-1:0] ox18q467wzh8vsuj = 
                                   jxpj6_9tx5iktrgs ? {2{1'b0}}
                                 : d2jsegrkoa154kuy ? (kwbmlmwj_ec + {{2-1{1'b0}},1'b1})
                                 : kwbmlmwj_ec;
  
  ux607_gnrl_dfflr #(2) opyi12br8u9_35k_ni (v0t2k69nbehh, ox18q467wzh8vsuj, kwbmlmwj_ec, gf33atgy, ru_wi);


  wire [5-1:0]      p_ikh0oqv24akv2uf7x1fjl    = hxvldlso5zpp81[4:0];
  wire [27-1:0]   iua4w9ohhqap05m4cd13br = hxvldlso5zpp81[(32-1):5];
  
  wire [6-1:0] f7igcfdxvo4ze3scv1f56l = iua4w9ohhqap05m4cd13br[6-1:0];
  wire [21-1:0]        x2i9sijf_tn1es8efcjsap3 = iua4w9ohhqap05m4cd13br[27-1:6];

  wire [2-1:0] kethvb4xg0vo30bsrgzwhhu = kwbmlmwj_ec + p_ikh0oqv24akv2uf7x1fjl[5-1:3];

  assign  z64bwdr23steb7s9y9j  = {iua4w9ohhqap05m4cd13br,kethvb4xg0vo30bsrgzwhhu,3'b0}; 
  assign  b7aet1zp_fcfxn8h7rw0u1 = 3'b010;

  assign  cneu8a119tg3vmie6zr2h_  = y4tsxz4rprpynubw3rvm;
  assign  jw2dzv9gi7gygudyqql6fz  = n7jh1zclcr_s0l4bgd;
  assign  o_7kpry6inkqpqi1bf1nd  = wunjscg6om1d0yu8o;
  assign  bg1spy6_v2kbo75pz1d6  = 1'b1;
  wire  q7k1vzcndghghxtpbf = bxc0qc1hr_cb1a4x1zadth;
  wire  cu9wchz0hcex50o2m_yx   = nlfdn3rz3118m7vvwo;
  assign  t3szwnvfo2nj3wk6r5kvt = {cu9wchz0hcex50o2m_yx,q7k1vzcndghghxtpbf};
  assign  xyeq7c6icdac80_y0jup = 64'b0;
  assign  za5ms2soyuucfxo_jbn = 8'b0;
  assign m4x1_gvw8v_sc8h7c8_6 = 1'b0;
  assign hpeqnhpztp9l_d3yx16l = 1'b0;
  assign bngbyv57e7juc0vkk2y8i = 2'b11;
  assign f97tgz_qybmvln6nz5dqt458 = 1'b0;
  assign znotwr53pu47f5m1agm = 1'b0;

  
  
  
  wire [2-1:0] m8e4y5p5zfei0w;
    
  wire bh0_09jdv_nabkpizd8n;
  wire rzjjndlw_np7otl63 = bh0_09jdv_nabkpizd8n;
    
  wire xp_8ug3xaxvs1hzjo4ime = (m8e4y5p5zfei0w == 2'b0);
  wire pcfm3_o_60ze1zpucjl = (m8e4y5p5zfei0w == ku4rkdvsjrgvr70b8i1e7dj7t7qedj[2-1:0]);
  wire xzheht9iavqj32dq7zx = bh0_09jdv_nabkpizd8n & pcfm3_o_60ze1zpucjl;
  wire ddht2k_7yytr_fa5yogp = rzjjndlw_np7otl63 | xzheht9iavqj32dq7zx;
  wire [2-1:0] csy24t9fh7gacp9f = 
                                   xzheht9iavqj32dq7zx ? {2{1'b0}}
                                 : rzjjndlw_np7otl63 ? (m8e4y5p5zfei0w + {{2-1{1'b0}},1'b1})
                                 : m8e4y5p5zfei0w;
  
  ux607_gnrl_dfflr #(2) ui0nyss5vsvizbzfh0s (ddht2k_7yytr_fa5yogp, csy24t9fh7gacp9f, m8e4y5p5zfei0w, gf33atgy, ru_wi);

  assign bh0_09jdv_nabkpizd8n = ze2bfnigu62i9937pcxnjc & c86b14qr2qo45_qw2ns;
  assign zqa26f3l044pht447ti8x_r8rmh = xzheht9iavqj32dq7zx;


  
  
  
  wire [2-1:0] abkco79gja8ucsoev2ubkpk2 = m8e4y5p5zfei0w + p_ikh0oqv24akv2uf7x1fjl[5-1:3];
  assign yp6atu2uzbb053onf7h7j_g3 = (zkqavy8j9jzdikz_29v7am & ze2bfnigu62i9937pcxnjc & xp_8ug3xaxvs1hzjo4ime);

  
  
  
  

  assign  c86b14qr2qo45_qw2ns = 1'b1;
  assign  p4dpiqc4w_g42ni5jsaj = 1'b1;

  wire [64-1:0] htccp96oizuk1a;
  wire [64-1:0] q0kf3wejj2ljn;
  wire [64-1:0] tw4im4bn8pi1ufhxz;
  wire [64-1:0] d6lpoh_00tk5e;

  wire gcz9x4cwo29b0qf36pij8;
  wire ubzlvoihm1c1uqa3t8;
  wire qk8lkfqbo_y1wy4gxq_;
  wire qudwatuvrp5y9d0nvgcrwp;

  wire k08eg8pj4df464__j0ipg_ = bh0_09jdv_nabkpizd8n & (abkco79gja8ucsoev2ubkpk2 == 2'd0);
  wire lp8b8bvgaau52roriib2d358s = bh0_09jdv_nabkpizd8n & (abkco79gja8ucsoev2ubkpk2 == 2'd1);
  wire b8aoll1aq0pcny4p8p3vchqa = bh0_09jdv_nabkpizd8n & (abkco79gja8ucsoev2ubkpk2 == 2'd2);
  wire v_6jdjelrr5zab3dksxlc6 = bh0_09jdv_nabkpizd8n & (abkco79gja8ucsoev2ubkpk2 == 2'd3);

  wire x4isgx7oe0184agqzzjmlr0y8m ;
  wire tb5ry0377l4br2og796q6b4vdwb;

  wire mhohb0lw3mcvzmi2ujll49x = tb5ry0377l4br2og796q6b4vdwb ;
  wire hs_j3lgya4fdwkg4a0sw = tb5ry0377l4br2og796q6b4vdwb;
  wire f22p64375noi3g4804r56smqf = x4isgx7oe0184agqzzjmlr0y8m ;  
  wire dwhsf5xpc4pie944568l5 = x4isgx7oe0184agqzzjmlr0y8m;

  wire[64-1:0] gpk4vhwx1y9syp2f87;
  wire[64-1:0] p_e7sa6_osd_xum1695xa;
  wire[64-1:0] d71p0fs4x5n9ihzq8ei4;
  wire[64-1:0] bul4dyiq6rmukxrz0;

  wire nj3n5yvnbk6y_p;
  wire xjfk40rs7og5b;

  p7k2hwgr9tazox9ivj695zpxhajkb x8e0k4tp6fo4g5t6psflu(
     .e5uheiss35t1 (nj3n5yvnbk6y_p),
   
     .i6_p95sqjet02(zkojor8433oflab2kpvtzi1z9),          
     .g8qh7ytfxpof4e_(nx6i4o0_cbqmlan1ylpodj9y),          
     .wt5ewwuq7uqf(tgfv2w2s7qhwkl0pdpf_79v4e),          
     .vxikm1a46oon(qfjl6250hpfb57pxl0t53q6fd),          
   
     .iw6t1cm4o67qw1(gpk4vhwx1y9syp2f87),
     .mggrpeuiih45(p_e7sa6_osd_xum1695xa),
     .n9lrm5b8dl_r2gg(d71p0fs4x5n9ihzq8ei4),
     .xq_xgf70o0nt0zy(bul4dyiq6rmukxrz0) 
   );

  wire jfsin5gv7n8szn0k7 = k08eg8pj4df464__j0ipg_ | mhohb0lw3mcvzmi2ujll49x;
  wire ouokwtt3n_xb7ylgueiz = lp8b8bvgaau52roriib2d358s | hs_j3lgya4fdwkg4a0sw;
  wire tvj67o0l_dwlcr85a = b8aoll1aq0pcny4p8p3vchqa | f22p64375noi3g4804r56smqf;
  wire gwwlucljdvaidu05z1c = v_6jdjelrr5zab3dksxlc6 | dwhsf5xpc4pie944568l5;

  wire  [64-1:0]    wrskvdxy06p_m2cq0zbb9a6k = {
                           {8{o8smcfmzt25hxpwcn[7]}},
                           {8{o8smcfmzt25hxpwcn[6]}},
                           {8{o8smcfmzt25hxpwcn[5]}},
                           {8{o8smcfmzt25hxpwcn[4]}},
                           {8{o8smcfmzt25hxpwcn[3]}},
                           {8{o8smcfmzt25hxpwcn[2]}},
                           {8{o8smcfmzt25hxpwcn[1]}},
                           {8{o8smcfmzt25hxpwcn[0]}}
                                      };

  wire [64-1:0] u_ciwfo83llp0rxtv555pm4sf0g = 
       (c3vtv1izxu7rm5646jsmmke & (~wrskvdxy06p_m2cq0zbb9a6k)) | (bl79n71wkynirgcs3 & wrskvdxy06p_m2cq0zbb9a6k);

  wire [64-1:0] tk7w6dok4ea3weblj6k65yczvj  = (ibt51xz_a6yo4yknr5mx1 & ze2bfnigu62i9937pcxnjc & xp_8ug3xaxvs1hzjo4ime) ? u_ciwfo83llp0rxtv555pm4sf0g : c3vtv1izxu7rm5646jsmmke;  

  wire[64-1:0] ctdf7z4eixqhewqg = k08eg8pj4df464__j0ipg_ ? tk7w6dok4ea3weblj6k65yczvj : gpk4vhwx1y9syp2f87;
  wire[64-1:0] bhaa9fd3j02i0yp2chs = lp8b8bvgaau52roriib2d358s ? tk7w6dok4ea3weblj6k65yczvj : p_e7sa6_osd_xum1695xa;
  wire[64-1:0] c4c5q97zhvs65kzi = b8aoll1aq0pcny4p8p3vchqa ? tk7w6dok4ea3weblj6k65yczvj : d71p0fs4x5n9ihzq8ei4;
  wire[64-1:0] vaocl_eo5fq1hbx = v_6jdjelrr5zab3dksxlc6 ? tk7w6dok4ea3weblj6k65yczvj : bul4dyiq6rmukxrz0;

  ux607_gnrl_dfflr #(64) jp7j25mzv137ltv_bj (jfsin5gv7n8szn0k7, ctdf7z4eixqhewqg, htccp96oizuk1a, gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(64) ewsdr009wlxsba3emmoh (ouokwtt3n_xb7ylgueiz, bhaa9fd3j02i0yp2chs, q0kf3wejj2ljn, gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(64) kg3ftodfsq5up58in (tvj67o0l_dwlcr85a, c4c5q97zhvs65kzi, tw4im4bn8pi1ufhxz, gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(64) ny94i35gumms2ahp38io (gwwlucljdvaidu05z1c, vaocl_eo5fq1hbx, d6lpoh_00tk5e, gf33atgy, ru_wi);

  wire bs0ils61i1jf336hjbfj0 = ue54sje856um8518nhjen;
  wire k6cw0tvmrjgoe4vr8d5l = bs0ils61i1jf336hjbfj0 | jfsin5gv7n8szn0k7;
  wire n6_95ppa9lyud2x2yky = bs0ils61i1jf336hjbfj0 | ouokwtt3n_xb7ylgueiz;
  wire a32zyyl0c1kzg5rixhrqdg4m = bs0ils61i1jf336hjbfj0 | tvj67o0l_dwlcr85a;
  wire dehb90ig_3bh4q6o81mcp = bs0ils61i1jf336hjbfj0 | gwwlucljdvaidu05z1c;

  wire lnla2rsa02zjg38nlyduu0u = bs0ils61i1jf336hjbfj0 ? 1'b0 : dm5b92mx0redfbuhs1u3d;
  wire lx6qt27bbez_a1wkg_ow489 = bs0ils61i1jf336hjbfj0 ? 1'b0 : dm5b92mx0redfbuhs1u3d;
  wire a57_4x81d8dt37c4vuc0hyn = bs0ils61i1jf336hjbfj0 ? 1'b0 : dm5b92mx0redfbuhs1u3d;
  wire wdr8jor7f52ovdvcmfdeovr = bs0ils61i1jf336hjbfj0 ? 1'b0 : dm5b92mx0redfbuhs1u3d;

  ux607_gnrl_dfflr #(1) f9el_6gkcy6rh2fdahjjd (k6cw0tvmrjgoe4vr8d5l, lnla2rsa02zjg38nlyduu0u, gcz9x4cwo29b0qf36pij8, gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1) dttu5ha0o2p28bjdm2r73i (n6_95ppa9lyud2x2yky, lx6qt27bbez_a1wkg_ow489, ubzlvoihm1c1uqa3t8, gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1) m3x17e4ogmdfndbpea2c1o9anl (a32zyyl0c1kzg5rixhrqdg4m, a57_4x81d8dt37c4vuc0hyn, qk8lkfqbo_y1wy4gxq_, gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1) xmztdiwvt3lv68asnv4vwdi1 (dehb90ig_3bh4q6o81mcp, wdr8jor7f52ovdvcmfdeovr, qudwatuvrp5y9d0nvgcrwp, gf33atgy, ru_wi);

  assign dkox2mp78q58i66 = | {dm5b92mx0redfbuhs1u3d,
                           qudwatuvrp5y9d0nvgcrwp,
                           qk8lkfqbo_y1wy4gxq_, ubzlvoihm1c1uqa3t8, gcz9x4cwo29b0qf36pij8}; 

  assign gl9dazcghkmei56i8tlb     = dm5b92mx0redfbuhs1u3d;
  assign k7x2rdsdsxkmoiyluje7bf2aa = c4cb28s8l8rdx2e53vww;
  assign j1utgrdwzlhqppb8rev5pbh55   = c3vtv1izxu7rm5646jsmmke;

  wire ocq75bq28525mfnvv3 = x4isgx7oe0184agqzzjmlr0y8m &   nj3n5yvnbk6y_p; 
  wire y9s3aw4yqt2n96ozqlle3 = x4isgx7oe0184agqzzjmlr0y8m & (~nj3n5yvnbk6y_p); 
  wire[21-1:0] ubap4so8ss9fe62gkt = ye256knohacnaakiw2nqck6[21-1:0];
  wire[21-1:0] r6bf4f_q4xmws67zfq2 = hyxeikuobvxjumz2hibay[21-1:0];
  wire[21-1:0] vt2imvvskb5o8v;
  wire[21-1:0] tpk635xyt5_b98sb5;

  ux607_gnrl_dfflr #(21) o86g1mbu5s38n6lt96fsl0a (ocq75bq28525mfnvv3, ubap4so8ss9fe62gkt, vt2imvvskb5o8v, gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(21) m5x9iq4mzo9th2fklrpqfi (y9s3aw4yqt2n96ozqlle3, r6bf4f_q4xmws67zfq2, tpk635xyt5_b98sb5, gf33atgy, ru_wi);

  
  
  
  wire euc0hml8qo;
    
  wire qewkz_tphc72x4 = imzw3o6xtgdmikumc & mxk6xl0c64kzkrplmm;
    
  wire ia2lrypcba = (euc0hml8qo == 1'b1);
  wire urnnwq3exu732b_7 = imzw3o6xtgdmikumc & mxk6xl0c64kzkrplmm & ia2lrypcba;
  wire lu3_mdbpbwqk = qewkz_tphc72x4 | urnnwq3exu732b_7;
  wire wucd_zlrkttqq7tt = urnnwq3exu732b_7 ? 1'b0
                    : qewkz_tphc72x4 ? (euc0hml8qo + 1'b1)
                    : euc0hml8qo;
  
  ux607_gnrl_dfflr #(1) dukvhgkkxbhmzupmq6 (lu3_mdbpbwqk, wucd_zlrkttqq7tt, euc0hml8qo, gf33atgy, ru_wi);

  wire   c5q77wvcrg77lxzfadlscie = mxk6xl0c64kzkrplmm & imzw3o6xtgdmikumc & (~ia2lrypcba);
  assign o_0q4jefxhht9mcddirs7  = mxk6xl0c64kzkrplmm & imzw3o6xtgdmikumc & ia2lrypcba;
  

  
  
  
  assign yhwk19tompbv5zx = tyxs3jzhr2i2gq9dt7 & zti98n829owa2p;

  wire vuspkrmkr7ac6f3f;
    
  wire ca7n91ul4ydrfr6y = yhwk19tompbv5zx & uafmsty4hif2k4iobx;
    
  wire fd5rrv7ic6cdoqs_w = (vuspkrmkr7ac6f3f == 1'b1);
  wire mudxg2vrnwn8hmfw = yhwk19tompbv5zx & uafmsty4hif2k4iobx & fd5rrv7ic6cdoqs_w;
  wire w3he0mrqvm0lhje8 = ca7n91ul4ydrfr6y | mudxg2vrnwn8hmfw;
  wire q1_gk1ih6ipf1zujs = mudxg2vrnwn8hmfw ? 1'b0
                    : ca7n91ul4ydrfr6y ? (vuspkrmkr7ac6f3f + 1'b1)
                    : vuspkrmkr7ac6f3f;
  
  ux607_gnrl_dfflr #(1) e_0v3l0ed44el9uxzp2ql4 (w3he0mrqvm0lhje8, q1_gk1ih6ipf1zujs, vuspkrmkr7ac6f3f, gf33atgy, ru_wi);

  wire ru6h4chgeola28s10mngd05o = yhwk19tompbv5zx & uafmsty4hif2k4iobx & l88go20t1nggrq383;
  wire xazv45h8k8zfgrzyfv7_lo = yhwk19tompbv5zx & uafmsty4hif2k4iobx & (~fd5rrv7ic6cdoqs_w);
  assign jzytexqffyvv5d75cjxbqox8  = yhwk19tompbv5zx & uafmsty4hif2k4iobx & fd5rrv7ic6cdoqs_w;

  assign x4isgx7oe0184agqzzjmlr0y8m  = ru6h4chgeola28s10mngd05o &   fd5rrv7ic6cdoqs_w ;
  assign tb5ry0377l4br2og796q6b4vdwb = ru6h4chgeola28s10mngd05o & (~fd5rrv7ic6cdoqs_w);

  
  
  
  wire srrihnqfodnx68_8p;
      
  wire op1lty0w05u47_ue = 
                         (imzw3o6xtgdmikumc & g1evvi19a50ju8wyn5) |
                         (imzw3o6xtgdmikumc & mxk6xl0c64kzkrplmm) 
                       ;
      
  wire eskn4dwrn91ydr6v7 = 
                         (jzytexqffyvv5d75cjxbqox8 & uafmsty4hif2k4iobx) 
                       ;
  wire w6_2112jo6slz0nwi = op1lty0w05u47_ue |   eskn4dwrn91ydr6v7;
  wire ihrglgkb_oiec80gz8 = op1lty0w05u47_ue;
  ux607_gnrl_dfflr #(1) tevelzi0q72gecaq_e (w6_2112jo6slz0nwi, ihrglgkb_oiec80gz8, srrihnqfodnx68_8p, gf33atgy, ru_wi);

  assign  jkq984ky8fozrzq = srrihnqfodnx68_8p; 



  
  
  
  
  wire moqwwz55ay2mifynbhha;
      
  wire lc2p52hlxbo03s74chc2h3by_7x = x4isgx7oe0184agqzzjmlr0y8m;
      
  wire iczcb7jh0plgt;
  wire bnctold1_kpqu9ty7uvqvu1 = moqwwz55ay2mifynbhha & iczcb7jh0plgt;
  wire dv3y_brlz73wxsp_qr80feq95 = lc2p52hlxbo03s74chc2h3by_7x | bnctold1_kpqu9ty7uvqvu1;
  wire cyrk1ifx52yk80i1agzm_rgfwo = (~bnctold1_kpqu9ty7uvqvu1);
  ux607_gnrl_dfflr #(1) e87f75bpb8_24b3quia3nonkmzony (dv3y_brlz73wxsp_qr80feq95, cyrk1ifx52yk80i1agzm_rgfwo, moqwwz55ay2mifynbhha, gf33atgy, ru_wi);

  assign  zf_v02okbs8_euhd64 = moqwwz55ay2mifynbhha; 

  wire i1n4qg6dqh8js3m3q4 = zf_v02okbs8_euhd64 & wq4r8m45isqp8_o4pdtitz;

  
  
  
  wire [2-1:0] xoyv6g81ld;
    
  wire o2baujz9fy9lp04n9 = i1n4qg6dqh8js3m3q4;
    
  wire wn8dn28ep04qnynezff = (xoyv6g81ld == 2'b0);
  wire z82owypbst_uwwtrgboq6 = (xoyv6g81ld == ku4rkdvsjrgvr70b8i1e7dj7t7qedj[2-1:0]);
  assign iczcb7jh0plgt = i1n4qg6dqh8js3m3q4 & z82owypbst_uwwtrgboq6;
  wire kedzfu6gdlxf1oze9 = o2baujz9fy9lp04n9 | iczcb7jh0plgt;
  wire [2-1:0] pkp2xtnc70_uvbb_v = 
                                   iczcb7jh0plgt ? {2{1'b0}}
                                 : o2baujz9fy9lp04n9 ? (xoyv6g81ld + {{2-1{1'b0}},1'b1})
                                 : xoyv6g81ld;
  
  ux607_gnrl_dfflr #(2) v110hc04afautx (kedzfu6gdlxf1oze9, pkp2xtnc70_uvbb_v, xoyv6g81ld, gf33atgy, ru_wi);


  wire[21-1:0] oxfs9oldqrys1nr = nj3n5yvnbk6y_p ? vt2imvvskb5o8v : tpk635xyt5_b98sb5;

  wire [6-1:0] clke8uwxp_988e = f7igcfdxvo4ze3scv1f56l;
  assign  qpzo6lin6brrytho7  = {oxfs9oldqrys1nr, clke8uwxp_988e, xoyv6g81ld,3'b0}; 
  wire [32-1:0] gkfif1c6_keasol5_mo2xgqdsa  = {oxfs9oldqrys1nr, clke8uwxp_988e, 2'b0,3'b0}; 
  wire [32-1:0] rlq163wp2nwj9ogopvjrznngih  = {iua4w9ohhqap05m4cd13br, 2'b0,3'b0}; 

  assign  ljk3q52m5tirt6shbcwbf = 3'b001; 

  assign  vvadj6ew1h5wq9z5askkzr9  = y4tsxz4rprpynubw3rvm;
  assign  lop06h0_z_4tt1s04up  = n7jh1zclcr_s0l4bgd;
  assign  ivllgcn1kiix2iamzwf0u  = wunjscg6om1d0yu8o;
  assign  k7j6g0757jovg8xstgrvwf  = 1'b0;
  wire  hvmgtgcbbqpzrp1a53bwy8 = wn8dn28ep04qnynezff;
  wire  vyjwuz8o2dx_1ja3nuy   = z82owypbst_uwwtrgboq6;
  assign  ucj9poqgl683ej1pihkh = {vyjwuz8o2dx_1ja3nuy,hvmgtgcbbqpzrp1a53bwy8};
  wire rpwi300et2o9udps5 = (xoyv6g81ld == 2'd0);
  wire cvfbtpik0hlvnec = (xoyv6g81ld == 2'd1);
  wire ikythk__cph6woz = (xoyv6g81ld == 2'd2);
  wire ca4ir_y7n32ykoj = (xoyv6g81ld == 2'd3);
  assign nwx86gohbrn08nvh60789 = (
                                (htccp96oizuk1a & {64{rpwi300et2o9udps5}}) 
                              | (q0kf3wejj2ljn & {64{cvfbtpik0hlvnec}}) 
                              | (tw4im4bn8pi1ufhxz & {64{ikythk__cph6woz}}) 
                              | (d6lpoh_00tk5e & {64{ca4ir_y7n32ykoj}}) 
                            );
  assign bebhplbk2k43sfoehvt66w = {8{1'b1}};
  assign u9hi0xtx8u0mn0l_7p = 1'b0;
  assign rm04yhu6ondli9u0g6din = 1'b0;
  assign o5fmtstd7kef7z4m7jefm = 2'b11;
  assign rnmvpk356vfgxd_045g = 1'b0;
  assign a46c4xo4texvc9o = 1'b0;

  
  
  
  wire [2-1:0] oq_1magiy3ybgw_8b;
    
  wire l82p7_8fgxootq8noll30l;
  wire m7fcspo0llkc4rmn = l82p7_8fgxootq8noll30l;
    
  wire ttondh96wgwhj24yho_jw9x = (oq_1magiy3ybgw_8b == 2'b0);
  wire bqnj6agg0tk79y19_k = (oq_1magiy3ybgw_8b == ku4rkdvsjrgvr70b8i1e7dj7t7qedj[2-1:0]);
  wire nq2p9gxwh3u7jn7fnzzr = l82p7_8fgxootq8noll30l & bqnj6agg0tk79y19_k;
  wire cnv2yd7kqjo_d6hk9q = m7fcspo0llkc4rmn | nq2p9gxwh3u7jn7fnzzr;
  wire [2-1:0] jw_c6fo4ptxemngzuyqa = 
                                   nq2p9gxwh3u7jn7fnzzr ? {2{1'b0}}
                                 : m7fcspo0llkc4rmn ? (oq_1magiy3ybgw_8b + {{2-1{1'b0}},1'b1})
                                 : oq_1magiy3ybgw_8b;
  
  ux607_gnrl_dfflr #(2) eou8lz8iryrj0ta64ecs (cnv2yd7kqjo_d6hk9q, jw_c6fo4ptxemngzuyqa, oq_1magiy3ybgw_8b, gf33atgy, ru_wi);

  assign l82p7_8fgxootq8noll30l = mm70cenjp_1wmcs135nh4wl & p4dpiqc4w_g42ni5jsaj;
  assign zxz6ihlgme0sknfg8ncdly9z = l82p7_8fgxootq8noll30l & bqnj6agg0tk79y19_k;


  
  

  wire ntw_ioifg95pt88xriadvf = ue54sje856um8518nhjen;

  wire h2hmhs04kszw1e73fudw = ntw_ioifg95pt88xriadvf | (l82p7_8fgxootq8noll30l & (oq_1magiy3ybgw_8b == 2'd0));
  wire yf13otuvp7gi4pr6lmxvz = ntw_ioifg95pt88xriadvf | (l82p7_8fgxootq8noll30l & (oq_1magiy3ybgw_8b == 2'd1));
  wire sk91b88y65v4roxq6h6_f6c3 = ntw_ioifg95pt88xriadvf | (l82p7_8fgxootq8noll30l & (oq_1magiy3ybgw_8b == 2'd2));
  wire qvez3_qw6ccuayii2re = ntw_ioifg95pt88xriadvf | (l82p7_8fgxootq8noll30l & (oq_1magiy3ybgw_8b == 2'd3));

  wire p659o1x0buon58ou4zgay = ntw_ioifg95pt88xriadvf ? 1'b0 : ezntrtg3q1must0tfcgn;
  wire pa24i69v4p8y_n3miq6pzuw = ntw_ioifg95pt88xriadvf ? 1'b0 : ezntrtg3q1must0tfcgn;
  wire u3lmyxkn_d10kigq23ck1v = ntw_ioifg95pt88xriadvf ? 1'b0 : ezntrtg3q1must0tfcgn;
  wire l3tdjf0opdq5k90mqusdg = ntw_ioifg95pt88xriadvf ? 1'b0 : ezntrtg3q1must0tfcgn;

  wire x1xuv11gx00j0evs7t6ry1;
  wire v1qdoewhc0q6k75k1ifk;
  wire av584m1rz376o0jdpg4n;
  wire o1y9e6yjncsm3t80m0eejc;

  ux607_gnrl_dfflr #(1) ts5i95hhj_pyifpgod758a1olx (h2hmhs04kszw1e73fudw, p659o1x0buon58ou4zgay, x1xuv11gx00j0evs7t6ry1, gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1) q51lx38s7w_pw_s6u9lcfb (yf13otuvp7gi4pr6lmxvz, pa24i69v4p8y_n3miq6pzuw, v1qdoewhc0q6k75k1ifk, gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1) iainlkizqkkauulv33586wh (sk91b88y65v4roxq6h6_f6c3, u3lmyxkn_d10kigq23ck1v, av584m1rz376o0jdpg4n, gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1) bm5j895aiwteuzafrdqb_2 (qvez3_qw6ccuayii2re, l3tdjf0opdq5k90mqusdg, o1y9e6yjncsm3t80m0eejc, gf33atgy, ru_wi);

  wire h9rwhx3dvgc9nc3h8o = | {ezntrtg3q1must0tfcgn,
                          o1y9e6yjncsm3t80m0eejc,
                          av584m1rz376o0jdpg4n, v1qdoewhc0q6k75k1ifk, x1xuv11gx00j0evs7t6ry1}; 

  assign g3_8p4g7w5grnl62xy = mxk6xl0c64kzkrplmm
                        | g1evvi19a50ju8wyn5 
                          ;

  assign imzw3o6xtgdmikumc = g3_8p4g7w5grnl62xy & vqwqaofc8sz_yjccd;

    
    
    
    
  wire yknrmk1dwifymi51 = ~ong4xrs8cubfol;
  wire hr4h3z6hojvm8hxfc7k =  ong4xrs8cubfol;
  wire q0kqweouhqcu2g_2 = (~e0ny5yl0v2ik890te) & (uhrfddgw6k1clj2oc |   x7jix80161slp ); 
  wire ew9_u8s1q6gmcuq1 = (~uhrfddgw6k1clj2oc) & (e0ny5yl0v2ik890te | (~x7jix80161slp));
  assign nj3n5yvnbk6y_p = s8iygpzng_5v9083x1skh1xq00434b6_ ? yknrmk1dwifymi51 : q0kqweouhqcu2g_2;
  assign xjfk40rs7og5b = s8iygpzng_5v9083x1skh1xq00434b6_ ? hr4h3z6hojvm8hxfc7k : ew9_u8s1q6gmcuq1;

  wire dcj2an8gay608_myt = (nj3n5yvnbk6y_p & tg3c0ha5844xz) | (xjfk40rs7og5b & dvn3st2c0wavqa6); 
  wire d_m5wnahz6811rvt3y  = (nj3n5yvnbk6y_p & e0ny5yl0v2ik890te)  | (xjfk40rs7og5b & uhrfddgw6k1clj2oc); 


    
  assign l88go20t1nggrq383 = s8iygpzng_5v9083x1skh1xq00434b6_ ? (eq6xz7m5lnl9uvy2 ? dcj2an8gay608_myt : 1'b0) : dcj2an8gay608_myt; 

  
      
  wire bklaemmjtx2y4kwclft = (j98f_s869qm5bv_dhgbcim3 & h9rwhx3dvgc9nc3h8o);
      
  wire kk81r9ixfaj5h3svk_3wifjjfne5 = (ibt51xz_a6yo4yknr5mx1 & ar7ss7g0h7o9d58_adekeyg & dkox2mp78q58i66);

  assign c9oejgc5s6_v8ooyy8c0x1 = bklaemmjtx2y4kwclft;
  assign m7rpuph0hm25ukmyralijiy = kk81r9ixfaj5h3svk_3wifjjfne5;

  assign izozgg91hphikoatw0xsa = 1'b0;  
  assign ck7dirv94s9jkefjfed0h0mp = 1'b0;  

  assign sktjnm1h7yu59cy6lnbf0gx40e_ = {{64-32{1'b0}},gkfif1c6_keasol5_mo2xgqdsa};  
  assign r_13gm13ck84al5d7ty5lf_m = {{64-32{1'b0}},rlq163wp2nwj9ogopvjrznngih};  

  
  
      
  wire l1nzgi1fse3cafcr2yi = imzw3o6xtgdmikumc & g1evvi19a50ju8wyn5;
  wire a35bayxb4ukd9rmpxf46q = l1nzgi1fse3cafcr2yi;  
  wire ts8s4jr4ph0f55rftwoqdz3va = l1nzgi1fse3cafcr2yi;  



  
  wire pxznrfv19o5tm3l = behhrrdejekhg_3v4ju ? 1'b0 : 1'b1;
  
  
  wire ix64b9ofahmqk31_ = pxznrfv19o5tm3l & (eq6xz7m5lnl9uvy2 ? 1'b0 : ibt51xz_a6yo4yknr5mx1 ? 1'b1 : 1'b0);

  
  
  
  wire b2fn0b6b_98odte = pxznrfv19o5tm3l & (p2kqppuunqlu40r ? 1'b1 : eq6xz7m5lnl9uvy2 ? d_m5wnahz6811rvt3y : 1'b0);


  
  

  assign a6gdkt5h77dh0mcj8t4gq = f7igcfdxvo4ze3scv1f56l;
  assign qtcasxm90cy0bwaqaxz = f7igcfdxvo4ze3scv1f56l;

  wire [3-1:0] arwn3azytv2k;
  assign arwn3azytv2k [2]  = b2fn0b6b_98odte;
  assign arwn3azytv2k [1] = ix64b9ofahmqk31_;
  assign arwn3azytv2k [0] = pxznrfv19o5tm3l;
  assign uh_ekyw7cw8c3d3xj1 = {arwn3azytv2k, x2i9sijf_tn1es8efcjsap3}; 
  assign f42g8ulc2y43ntmai5 = {arwn3azytv2k, x2i9sijf_tn1es8efcjsap3};          

  
  
  
  wire [64-1:0] yxa9r0cr3smxr383cjacv = (~fd5rrv7ic6cdoqs_w) ? htccp96oizuk1a : tw4im4bn8pi1ufhxz; 
  wire [64-1:0] je52cr2irpjui5zk7f_c4m = (~fd5rrv7ic6cdoqs_w) ? q0kf3wejj2ljn : d6lpoh_00tk5e;  

  wire vpfe1f6au = g3_8p4g7w5grnl62xy ? ia2lrypcba : fd5rrv7ic6cdoqs_w;

  wire e3bo9qay_vlwu2e6v = (
                         (l88go20t1nggrq383 & imzw3o6xtgdmikumc & mxk6xl0c64kzkrplmm) | 
                          (yhwk19tompbv5zx & uafmsty4hif2k4iobx & (s8iygpzng_5v9083x1skh1xq00434b6_ ? 1'b0 : 1'b1))
                      );

  wire vf99c0pc80jq7is8g67q = (
                         (l88go20t1nggrq383 & o_0q4jefxhht9mcddirs7) | 
                          jzytexqffyvv5d75cjxbqox8 
                  );


  assign j2kcz1faqhvh1ler6j = a35bayxb4ukd9rmpxf46q | (nj3n5yvnbk6y_p & vf99c0pc80jq7is8g67q);
  assign uf44audysjgtvdnua67 = ts8s4jr4ph0f55rftwoqdz3va | (xjfk40rs7og5b & vf99c0pc80jq7is8g67q);


      
      
  wire g7u0q4_wwj_ = (tyxs3jzhr2i2gq9dt7 & uafmsty4hif2k4iobx) ? 1'b1 : 1'b0;
  assign wixbtbeqlhzelg4t  = g7u0q4_wwj_;
  assign y38seii6ja77q2jy08  = g7u0q4_wwj_;





   y5gz1t0e4pyw9jr0abfow4_gfn1kng3 mzfkek7zy3821ly5v5(
    .dpjdlj8bv4q  (nj3n5yvnbk6y_p),
    .vhqr9jgt5  (e3bo9qay_vlwu2e6v),


    .vpfe1f6au (vpfe1f6au),
    .g7u0q4_wwj_ (g7u0q4_wwj_),

    .u4amtcbhq_6g6rx9 (f7igcfdxvo4ze3scv1f56l),
    .sm0ktbr6as2sl7ho(p_ikh0oqv24akv2uf7x1fjl),

    .xduvlstjiiwj (yxa9r0cr3smxr383cjacv),
    .pbu6py7mm4i (je52cr2irpjui5zk7f_c4m),

    .rl_3d1m7gcc0  (rgf8pa4kn20jusruz),
    .tsdapc3y0fh  (r2tvaf8px0p9vlw4we),
    .mohep6fqp67x  (rzf167thmprvps0tm62i),
    .mmmu7pm6e_uqx  (caxkrdjq0tjnnne9),

    .e6rwnjewsq6s6oro (frkunk72hlttw0ar0np),          
    .u74ed5k2tobo (svj88sv2u56fepzmg),          
    .cthiem_1bgmj (hat38salswlktk821),          
    .dg5w1zgjmlq1a4n (c0xnu9p8he2hw10h),          

    .ft2vjq7oh7l1hzqu (z6udkjbx164gh9yo1o),          
    .wbr3gkcxil8f_hgq (a_u2kfmgv2ho357c),          
    .t1ncj092lli (oj5t3f0lq1n9ae82x),          
    .vhh7ujoe4fwn_8 (v8jl1eh8o0n5g765),          

    .e_9jhaby2__46fj(wjwjffxr_4lulivwz),
    .lpcj6ymxsst2n(srfn4smswwo6hbyaa),
    .wdb90nca460cp(lv7fu0hif2n2zhmgtcc),
    .rin3amuhzyhjgg(qpuk8ry0w9_r7ur4gcnx)
);


  assign zti98n829owa2p = 1'b1;


  assign tyg8z9t16af4e8xtdiw = r2dy3qdfqfohba22hlsf5 & (z8alxhlwgz117[32-1:5] == qpzo6lin6brrytho7[32-1:5]);
  assign qkl9_olndwlohzaurunzkg = r2dy3qdfqfohba22hlsf5 & (q4j831gvqooep12[32-1:5] == qpzo6lin6brrytho7[32-1:5]);

  assign kd96ha16hcj4wyo0 = xjfk40rs7og5b;
  assign j9kszxa35hle0cl9 = (~s8iygpzng_5v9083x1skh1xq00434b6_) & jzytexqffyvv5d75cjxbqox8;
  assign myqlprv648_pqf92vvj = f7igcfdxvo4ze3scv1f56l;

  assign zpdvh58o0evhzt            = p2kqppuunqlu40r & jm4__y98e00ukvb4hiw_f;
      
  assign q0duv6epk3ccff620vhhx2     = zpdvh58o0evhzt  & hcnuxviddm5zvn0cyzv7m & dkox2mp78q58i66; 

  assign rpkosm9pbcpggwup90_ge9     = (reffh2y56n2410r_6a54c | lkkimoh3n0l0cploih) & jm4__y98e00ukvb4hiw_f;
      
  assign xwmkl_9n7oehwe7hh_a6aompojzukuik = reffh2y56n2410r_6a54c & h9rwhx3dvgc9nc3h8o;

endmodule





















module gsmnxrg40o2b1e4gc(
  output a03er8qo6p0zpb           ,
  output z8uuyp_3l6aqut86nkd__vvwgs    ,
  output bzsjo5unerpy5i0e_q_6eqn       ,
  output ctfhepdgvm53k59kbbe0s0924he0ijd,

  output                               hv39pppvbmeqy8b6,
  output[32-1:0]          t6l88yqbe4wokkhiso9t,
  output                               hyec__ebnw8lbcssd81,
  output                               vs2610q9_on1r996p,
  output                               coy3buxdw6yq3duh21azuwflk,
  output                               r_8h5lxb39ug57zli04e_o,
  output                               pv7q0ikpayogkay57rgyr,
  input                                dsq8f3rhmb7yc876v8,
  input                                enu_vumk17eoj1fma5ilz0,

  output                               ou74jmm5p6th0y0kcdwpqv2ey,
  output                               adwzzx09c_s_x1seh,
  input                                zp0aylmm0k4yw4w561bgzh,


  output tq5w2fd0flcywep677l,
  output juwj_oo3r8yt2a4hg,
  output k6_e3_saw0oup16pudov,
  output pzfb_24lrjd770iigjx4sm,
  output [6-1:0] zpq6nysk8b654ynyt4zj9k,
  output [6-1:0] d2lstp52x9w9900ioarrtfk,
  input                            cgnsvvj7srbljqst,


  input                           sej7ti3911672ok72k,
  output                          z2s7c4x2upx2k94,
  input  [32-1:0]    hdwldkfk3vetnqg3us, 
  input                           kix9_o92mst68vescu79v, 
  input                           ihkz9tebg3jd5f47z, 
  input                           tu1v8ryo2rv95crsvz, 
  input                           ghikvq604upn2v,
  input                           t4leke6w3uzo3gxu3yhk, 
  input                           oodqv7hv99boddj3kk48j, 
  input                           g2x5gi27ly4aw24, 
  input                           g16len3w2wk22u, 
  input                           vx_fynrmojs7gx, 
  input                           xpd4oma8mrw21r9b0mc8c, 
  input                           ytx0p13ahjuk751e8crl_0, 
  input  [64-1:0]       uacpumgrbwt0fmb,
  input  [8-1:0]       v0uq3fcdfb8eatt3,
  input                           c4otadutq6rav14ed2,     
  input                           mw8uaelv0i5zfav,     
  input  [1:0]                    uq0oocqz_ys0no4o_t,
  input                           ohprpkw231g_f2qqzmq,
  input                           e3l8n6__k56uw5o7jujwibr,
  input                           rwmac6nity_ikz7xbj_ta1nce,
  input                           en9ogfq6nx_uirma3y2jiigbh,
  input                           t9otq6y33fc5qs21p9d2rc3zn,
  input                           xpbzeko14yty79dehft9e2l,


  output                          r57mgw9ntmg26lxok,
  input                           cac59gne730vqiq,
  output                          ypuolenm4dvdg,
  output                          yu5m552dobcb8gbsq,
  output [64-1:0]         bo_q_t246zgg3q, 
  output [32-1:0]    d4k4iwwrjuzjqt, 



  output                          ktkt_7t0wo1gkg8gormhm,

  output                          rjy1ysvx9590bpklijsn0ucgaga,
  input                           d_933icutbtk8nknxip5t1ds,
  output  [32-1:0]   a45qubts5uovcopirpl9jxs7uia, 
  output                          kwbu6olmnnt53fot6kfntm2q7t, 
  output  [64-1:0]        kq9lkjt85jst7fa5smg1nud,
  output  [8-1:0]     mekhipn8vmxn5adno3jrpek8nkm,
  output  [2:0]                   wbwviedmyjzfiwi2t1yh0ibf7wv3,
  output  [1:0]                   h99v8xeu9gkycpsn1wl3lrow7,
  output                          jvloelo3plm6zwbisesi7fwa,
  output                          ecz8u30wtuyonhyfwfrfrc30g,
  output  [1:0]                   vxwea8jbxv6m5tu7nkqtf6,
  output                          jsswxoezxjsdw154f5xt1omqrup, 
  output                          e5cyxxxkg4061gq3_ksqdax_7op, 
  output                          m3pduyvpfh4ximuy0dl6k_wjuc, 
  output                          xhts19tgn12c186fduss6cfjyz, 
  output                          zt7xddfgq3m2nsc8s_3a48r8, 

  output                          s9lcmqjp282zoimy_nw6kv2u,

  output                          pkm6vgcr8iz_el5103gzwdew0hki,
  input                           vdbkch1krpijvuukam8k5_9g6h4d,
  output  [32-1:0]   gi8g2jgc5r69ozgg2517f4, 
  output                          nqq4y60r7eh5lbir_nzlqf2q7k, 
  output  [64-1:0]        rf_rtoowzj9m6zi6taqyqn6ku,
  output  [8-1:0]     kqa4ro7t84z342uqr2plzmi1,
  output  [2:0]                   d50l6nnxdfj7iuhnqe9gjobewaj4,
  output  [1:0]                   ziqf65e93q9kc_6bj_n4gd2op,
  output                          lkflakila483fdjdz1hrtobjiz,
  output                          zg0qkr8fhe1v0eku3at17q,
  output  [1:0]                   gu2ufdscjjb3hvpwrwu6c8h,
  output                          pn9rf9nl21n4t8clpsygzbo72n, 
  output                          u6t2h_hm580phvwuvdedyagaqg, 
  output                          h1p8zhyrvirdo9c78wx8cmal83, 
  output                          d11v3v5k967aul6l7_up53azs, 
  output                          tnfd_mhtdr0hw58lveup8w8, 



  input                           fp_qm6eq7380_uydc6pb2sw7,
  output                          z9eviza6dmjc6u7jbuzirzh8z1ce,
  input                           gz2qngl9towiwc_nk48gu38p9  ,
  input                           saolr4xnpfm570snrsqk7hazshkz,
  input [64-1:0]          b85cqul2sjbg0c5ta0bcpgpluvma, 

  input                           me8sa0hl_2m6xmtdm4r_1tn7cer4,
  output                          gv_wy8qy9rm50mn4yg66yvagb60l,
  input                           byn2o0bi_9ggzegrnvskn  ,
  input                           m12x1nn4kvsdeqofo9rqi8aawa,
  input [64-1:0]          e0xiuuzhk1qbwdjlub9o_cca5, 


  output                          tjzl_75hfxv6m,
  output [64-1:0]    ay20xnz1tx3gv1k,  
  output                          fyo0ut7e82c,  


  output                          jkq984ky8fozrzq,
  output                          g3_8p4g7w5grnl62xy,
  input                           vqwqaofc8sz_yjccd,

     
  input                           tyxs3jzhr2i2gq9dt7,
  output                          zti98n829owa2p,
  input  [24-1:0]  ye256knohacnaakiw2nqck6,
  input  [24-1:0]  hyxeikuobvxjumz2hibay,
  input  [32-1:0]  zkojor8433oflab2kpvtzi1z9,
  input  [32-1:0]  nx6i4o0_cbqmlan1ylpodj9y,
  input  [32-1:0]  tgfv2w2s7qhwkl0pdpf_79v4e,
  input  [32-1:0]  qfjl6250hpfb57pxl0t53q6fd,
     
  
  output                          j2kcz1faqhvh1ler6j,  
  output [6-1:0]  a6gdkt5h77dh0mcj8t4gq,
  output                          wixbtbeqlhzelg4t ,
  output [24-1:0]  uh_ekyw7cw8c3d3xj1,          
   
  output                          uf44audysjgtvdnua67,  
  output [6-1:0]  qtcasxm90cy0bwaqaxz, 
  output                          y38seii6ja77q2jy08 ,
  output [24-1:0]  f42g8ulc2y43ntmai5,          

  
  output                           rgf8pa4kn20jusruz,  
  output [8-1:0]  wjwjffxr_4lulivwz, 
  output [4-1:0]  z6udkjbx164gh9yo1o,
  output [32-1:0]  frkunk72hlttw0ar0np,          
                                   
  output                           r2tvaf8px0p9vlw4we,  
  output [8-1:0]  srfn4smswwo6hbyaa, 
  output [4-1:0]  a_u2kfmgv2ho357c,
  output [32-1:0]  svj88sv2u56fepzmg,          
                                  
  output                           rzf167thmprvps0tm62i,  
  output [8-1:0]  lv7fu0hif2n2zhmgtcc, 
  output [4-1:0]  oj5t3f0lq1n9ae82x,
  output [32-1:0]  hat38salswlktk821,          
                     
  output                           caxkrdjq0tjnnne9,  
  output [8-1:0]  qpuk8ry0w9_r7ur4gcnx, 
  output [4-1:0]  v8jl1eh8o0n5g765,
  output [32-1:0]  c0xnu9p8he2hw10h,          



  input  [32-1:0] z8alxhlwgz117, 
  input  [32-1:0] q4j831gvqooep12, 
  output yafkacaefbdmi3hm6rvuao, 
  output u4frf_hcy8c0dh_aqkgsrp, 
  

  output bda77mp8zde61a_,
  output tlwo81ky1a6b8,
  output l9x1ubg9wznb6ixv1i,
  output y5otpn351odm3mnpnfdshm,
  output rnlnwebfnqcg8g5oq_2gv0,

  input  gf33atgy,
  input  ru_wi
);

  localparam nsy582liduihtlix7j5       = 9;

  localparam d8ba36mdzefszkfe3pwmzqxhwx  = 3;
  localparam fumremxmy8mtkpij650zgfe79i  = 1;
  localparam yy567yahzg = 2;
  localparam yjbrpsqyidt47leh_ = (2-1);


  localparam qrt6p0l7zsi7heuq = (8 + 1);
  localparam ynlkel_xoan9ow       = 3;




  wire  [3-1:0]  pwi4opocymgcqmwe_vq4sm0; 
  wire  [3-1:0]  tq4o19u3oc43c2v2sc9hsityj; 

  wire  [3-1:0]  nc91g6pv91sa5ofkv6oqrzywy; 
  wire  [3-1:0]  p738fnhowqrqokqjpa0a748b; 

  wire                          zfu2vonacwweg65jwl5h;
  wire                          ecc0pa6dsujd5fk_ztk1odty;
  wire  [32-1:0]   t60xfh0jvayj7nnp_3swk1v; 
  wire                          p2m0mydv1zb_6iqetg5; 
  wire  [64-1:0]        a01toa5fu8pmct9z1qeb;
  wire  [8-1:0]     ex_5rp8vtq6iwx6hm_w;
  wire  [2:0]                   m_zge7ydxw1me0bp66_b;
  wire  [1:0]                   vo4iscd43mm129ts9g7;
  wire                          n5ajmphmp207ybl3ru6ee3p;
  wire                          r_te1f8papt089n46s6j2k;
  wire  [1:0]                   ao8xdzkmlvr9h6inuey9k;
  wire                          b6c9ysz1s8lqf83mno84; 
  wire                          gam1zdrkynr0puyhapwkq5fs; 
  wire                          w_bo91bpxaukiy9s3fyc9ib6; 
  wire                          yivyo1xc3okylkdzlkar; 
  wire                          acdtgtj2r5zy7qoh9ukv; 

  wire                          ejbq7zgkpgwgttfvvx5rp;
  wire                          agtve46c928tzy8367oy14bf;
  wire  [32-1:0]   pii5a6cmz40r9w30q_awu; 
  wire                          m6vmtqf14m_q0ahhpf9ys0t; 
  wire  [64-1:0]        hn4lhm3a_wcnqbxq84q;
  wire  [8-1:0]     pqhi5t7t91o9xtpy8r4_9o;
  wire  [2:0]                   zhc7g2_tfy2pqp2f8g5;
  wire  [1:0]                   edt_9_yofk03w8y7jt;
  wire                          zeqnplthuo3przg6v7sc;
  wire                          ia_e66cu_no6wwvfzv;
  wire  [1:0]                   ceg6dnmky0mxytf2e9bhe0;
  wire                          x934mbk53lq9pp23th7n5no0; 
  wire                          qw8c56hyyf3o9z35eb8m; 
  wire                          tpkr0onb62gbg0ddt7_pz4l; 
  wire                          j_e7kc3w9drko64cvqn5g; 
  wire                          fz8l_vym0or20pcgjct; 

  wire                          z9q40jbnm38zcodsjsd090z;
  wire                          i0znoodcvzhh4rexar7joqvk;
  wire                          g5a675dzhov32an3m  ;
  wire                          efz5oj5hqaeq_wptcenc10fq7;
  wire [64-1:0]         bhhfkcv51hmdpdenvztypn; 

  wire                          gcan4qd32d7splx9secvc8b;
  wire                          q2_zn_ozuoxddlj2se_t45w;
  wire                          ng9lxc1zr1snbj1p1b9  ;
  wire                          nykvnvl0i96asmogcmhlrpy;
  wire [64-1:0]         b_7_y71ywtomguvgnoq5; 

  
  wire                          zsp7u2uqvojc8zqnw0k6_p;
  wire                          mljh30sszwrhguqyc4f5e77l4;

  wire                          yp6atu2uzbb053onf7h7j_g3;
  wire                          vydbpbb7_kmw71ncfvuvj74;
  wire                          gl9dazcghkmei56i8tlb  ;
  wire                          k7x2rdsdsxkmoiyluje7bf2aa;
  wire [64-1:0]         j1utgrdwzlhqppb8rev5pbh55; 
 
  wire  [3-1:0]   pne0i0g6_hms5_ag22zyfpdmpf3; 
  wire  [3-1:0]   vk3aoj6halc2m4mdlurcg7joxd; 

















  localparam yvxy18k82q = 8;
  localparam q_x9wrwj4_y9o_9go_pa = (8-1);





  wire [8-1:0] kyu0c7rbs3tzasd;
  wire [8-1:0] m64tp4jpwoadr8w;
  wire [8-1:0] x5p4oi1vgjp37abo6;
  wire [8-1:0] iexhykoj1n453;
  wire [8-1:0] puxm_ue7jwuwh72gi;
  wire [8-1:0] g53evua7d3gpxw3;

  wire [8-1:0] welnckam1xqornvo_[8-1:0];
  wire [8-1:0] j23uvqn5e9vkkw0w2fht[8-1:0];
  wire [8-1:0] pnedptzdy93p4krxqb_p[8-1:0];
  wire [8-1:0] b700gcu8o4ko92g1i7kcc[8-1:0];
  wire [8-1:0] b2rl4ox_6rp8po4j2tz  [8-1:0];

  wire [8-1:0] f__yd2_rd0i7mgsj05bn;
  wire [8-1:0] buxvgnamnlcw3lpbel0;
  wire [8-1:0] d763qyon3q45pdbxztuo4;
  wire [8-1:0] asf2z47ldhqkwm15lbpzc;
  wire [8-1:0] kcgdolb8q4gs6fitbr3v_;

  wire [8-1:0] u5zzpdddo7nx53kgpobe;
  wire [8-1:0] ckambm7sahfb9bg1nm;
  wire [8-1:0] i801bchffjgm2eeav1c0;


  wire [8-1:0] ttgaf1h84fzp0d1oel7;
  wire [8-1:0] pup241nwugqoxaddw6o;
  wire [8-1:0] j6x4yktmu5u6_uil;
  wire [8-1:0] o8btl8op6tng90p0h;
  wire [8-1:0] n7nx9bfxwcqwv7;


  wire [8-1:0] mnch_edao2_c4_ni2;
  wire [8-1:0] ttgsuta_ewmr6;
  wire [8-1:0] ny0n30vi0dzifq_o;
  wire [8-1:0] cgst_q5rcj_eo2wfk;
  wire [8-1:0] n3k7lk4c5q;


  wire [8-1:0] mwvgay3ta4a2;
  wire [8-1:0] os4b0yseamo1t;
  wire [8-1:0] brv_ewhw27bxxr_;
  wire [8-1:0] rkx1mrv8yqxi8el;
  wire [8-1:0] a672uxn3mwn;

  
  wire [8-1:0] g7qqd7ejlmjzz7uab;
  wire [8-1:0] tg8y2zr5rfj4sw1xke8;
  wire [8-1:0] vkzm86ii21rro827o0;
  wire [8-1:0] oosv_ui3yrxrqb_nh89;
  wire [8-1:0] l_ldkrkpn59v4mhb_;

  wire [8-1:0] v84iwz704r1326150y;

  wire [8-1:0] ixtmkj78nheu_ghv7byt0w;
  wire [8-1:0] fa8x97zn7g9lhjdunyuqg;

  wire [8-1:0] w8u6pj2octqg9n0vi6;
  wire [8-1:0] ea8x6ufv3q0voque2u5o8;

  wire [8-1:0] e0umr420ntwlczrjba;
  wire [8-1:0] d7roxn5jsm8p278tf;

  wire [8-1:0] y206os9wqkqs1a7zyv;



  wire  [32-1:0] haaqh6wjlwi9jhnl     [8-1:0]; 
  wire                        xzc0imuvetgbn8    [8-1:0]; 
  wire                        halyb9c30hal    [8-1:0]; 
  wire                        pllepw4azlfujoh_i    [8-1:0];
  wire                        d1rzzdht0dlkdfjvs420q    [8-1:0];
  wire                        hwwn5fuw1ki6rpxis    [8-1:0];
  wire                        dmjcrnz0ai9_04   [8-1:0]; 
  wire                        t54w0z3ee_q       [8-1:0]; 
  wire                        a2oenic4uandesr_k9qocfw       [8-1:0]; 
  wire                        qp1mbsaizjipsj6     [8-1:0]; 
  wire                        rg7cda_918ahdww6p56mv81qg_     [8-1:0]; 
  wire                        v1bfb0aqght1_yfm5znt     [8-1:0]; 
  wire                        c3mjay1nkztzsfo3mf2     [8-1:0]; 
  wire                        cuslzq6_3njc_9dr     [8-1:0]; 
  wire  [64-1:0]    vsfpyprm4rivny0n4    [8-1:0];
  wire  [8-1:0]    zrhld0y35qav    [8-1:0];
  wire                        epo0qysbvw4gkmi     [8-1:0];     
  wire                        c274s6asp6_ptv     [8-1:0];     
  wire  [1:0]                 bx9szwl63ur     [8-1:0];
  wire                        knyt1bhi0tp16v3 [8-1:0];
  wire                        di2o65qovx5zvsf3rujmc [8-1:0];
  wire                        fizjb37qgnqc11y3usvo1jd8 [8-1:0];
  wire                        te3sgyqybgiz02r496eiram [8-1:0];
  wire                        hotgsfmzxnfg6u691gfcuem [8-1:0];
  wire                        dej8khi216rqhe3ebb4 [8-1:0];
  wire                        bk8m_k0vayvzu1ytxtuvky [8-1:0];

  wire  [64-1:0]    ypal30idlttlfu9s_qrvo    [8-1:0];

  wire                        xezq29zs58h59dv     [8-1:0];
  wire                        hmqlykdc12wo5_r73zg8 [8-1:0];

  wire  [64-1:0]    b9i1i44zz7lsiekhgww  [8-1:0];


  wire [3-1:0] gtbu9zcij35aw_0ph1j;


  wire [3-1:0] jgfckxgs0fo048;


  wire [3-1:0] s8ol0xfe2arkosb;


  wire [3-1:0] fnvtppgr2s0i78;


  wire [8-1:0] zlgnht9uo2fb7p;
  wire [8-1:0] yel5kfjrg5ib6;

  wire xnmbaecrrzbadq6w;

  wire yed5vav_1mz5nme_ = 1'b1;

  wire blwju8dk7oqctm5;
  wire tm4v0w70xpfbnl8980;

  wire c62fn41h9xt61kf = sej7ti3911672ok72k & z2s7c4x2upx2k94;
  wire cz_zhjm1li1y_udg = blwju8dk7oqctm5 & tm4v0w70xpfbnl8980;
  wire nt8ye4twu46q1ra9 = r57mgw9ntmg26lxok & cac59gne730vqiq;
  wire rl6bkzjo4zmfl3x = xnmbaecrrzbadq6w & yed5vav_1mz5nme_;

  wire wf8kpn_u83u2_gj9bsb = c62fn41h9xt61kf;
  wire p_hc6rswvpztv26i = rl6bkzjo4zmfl3x;

  wire huqvm9m1hvosa8sc4xjt;

  wire w3ss3ti2t0dj2tvx = cz_zhjm1li1y_udg;
  wire k23tmhod3m0plvdlp = nt8ye4twu46q1ra9 | huqvm9m1hvosa8sc4xjt;




  wire nynvaiovg4pie7ruixtjath;
  wire qri2yyksd_33u_zx9tmmo = ~nynvaiovg4pie7ruixtjath;
  wire iq0_stqcjlb0emx654f0dk = (gtbu9zcij35aw_0ph1j == q_x9wrwj4_y9o_9go_pa[3-1:0]) & wf8kpn_u83u2_gj9bsb;

  ux607_gnrl_dfflr #(1) lg_sd24qiy5gzxm32adh286j7 (iq0_stqcjlb0emx654f0dk, qri2yyksd_33u_zx9tmmo, nynvaiovg4pie7ruixtjath, gf33atgy, ru_wi);

  wire [3-1:0] uiml967ah3fw9vrc3; 

  assign uiml967ah3fw9vrc3 = iq0_stqcjlb0emx654f0dk ? 3'b0 : (gtbu9zcij35aw_0ph1j + {{3-1{1'b0}},1'b1});

  ux607_gnrl_dfflr #(3) kfpcc28arqmpkgegqy5f (wf8kpn_u83u2_gj9bsb, uiml967ah3fw9vrc3, gtbu9zcij35aw_0ph1j, gf33atgy, ru_wi);



  wire llbze9tcjwisi3ez26o;
  wire mlv5k08kf3rdk49ynxiyukcvr = ~llbze9tcjwisi3ez26o;
  wire l9zxwry2rkdqbd9t1stozgw9d = (jgfckxgs0fo048 == q_x9wrwj4_y9o_9go_pa[3-1:0]) & w3ss3ti2t0dj2tvx;

  ux607_gnrl_dfflr #(1) ku18ifaqt2n0vvgdvb6i0oz (l9zxwry2rkdqbd9t1stozgw9d, mlv5k08kf3rdk49ynxiyukcvr, llbze9tcjwisi3ez26o, gf33atgy, ru_wi);

  wire [3-1:0] z4_eazngbw1kzt4di; 

  assign z4_eazngbw1kzt4di = l9zxwry2rkdqbd9t1stozgw9d ? 3'b0 : (jgfckxgs0fo048 + {{3-1{1'b0}},1'b1});

  ux607_gnrl_dfflr #(3) n9khdda4c5ce7f0ez_s5v0 (w3ss3ti2t0dj2tvx, z4_eazngbw1kzt4di, jgfckxgs0fo048, gf33atgy, ru_wi);



  wire j4rv0c1p5ke7krinra;
  wire m5ryw3seisurjxzarj03_e = ~j4rv0c1p5ke7krinra;
  wire y6ch3w746a2o9xh6rgtesaap = (s8ol0xfe2arkosb == q_x9wrwj4_y9o_9go_pa[3-1:0]) & k23tmhod3m0plvdlp;

  ux607_gnrl_dfflr #(1) a8yrgavnklzhe9lh1nm81ncj (y6ch3w746a2o9xh6rgtesaap, m5ryw3seisurjxzarj03_e, j4rv0c1p5ke7krinra, gf33atgy, ru_wi);

  wire [3-1:0] vmas7nkwq48y8ugl2co0d; 

  assign vmas7nkwq48y8ugl2co0d = y6ch3w746a2o9xh6rgtesaap ? 3'b0 : (s8ol0xfe2arkosb + {{3-1{1'b0}},1'b1});

  ux607_gnrl_dfflr #(3) mjylwfiae8dfustolnvqz4 (k23tmhod3m0plvdlp, vmas7nkwq48y8ugl2co0d, s8ol0xfe2arkosb, gf33atgy, ru_wi);



  wire pn2h5gfpc4kw0y66t9;
  wire d5jrixpw82rcyxb77lqvpjt = ~pn2h5gfpc4kw0y66t9;
  wire hy_qezp81icfs3e8q66_zj = (fnvtppgr2s0i78 == q_x9wrwj4_y9o_9go_pa[3-1:0]) & p_hc6rswvpztv26i;

  ux607_gnrl_dfflr #(1) ewhzmr84uhd837_1ww13puh2w (hy_qezp81icfs3e8q66_zj, d5jrixpw82rcyxb77lqvpjt, pn2h5gfpc4kw0y66t9, gf33atgy, ru_wi);

  wire [3-1:0] ezrpbzwi3v7u6fhcl3; 

  assign ezrpbzwi3v7u6fhcl3 = hy_qezp81icfs3e8q66_zj ? 3'b0 : (fnvtppgr2s0i78 + {{3-1{1'b0}},1'b1});

  ux607_gnrl_dfflr #(3) uvdo2wx6icjwr698e11ob (p_hc6rswvpztv26i, ezrpbzwi3v7u6fhcl3, fnvtppgr2s0i78, gf33atgy, ru_wi);

  assign bda77mp8zde61a_ = (fnvtppgr2s0i78 == gtbu9zcij35aw_0ph1j) &   (pn2h5gfpc4kw0y66t9 == nynvaiovg4pie7ruixtjath);
  assign tlwo81ky1a6b8  = (fnvtppgr2s0i78 == gtbu9zcij35aw_0ph1j) & (~(pn2h5gfpc4kw0y66t9 == nynvaiovg4pie7ruixtjath));


  wire [3-1:0] jbuu2xdq0qw_wi19r = p_hc6rswvpztv26i ? ezrpbzwi3v7u6fhcl3 : fnvtppgr2s0i78;
  wire [3-1:0] ytx4fsx0_lffvqrj = wf8kpn_u83u2_gj9bsb ? uiml967ah3fw9vrc3 : gtbu9zcij35aw_0ph1j;
  wire r5bo9n9q6a8c5e5mv29k6wr = iq0_stqcjlb0emx654f0dk ? qri2yyksd_33u_zx9tmmo : nynvaiovg4pie7ruixtjath;
  wire ofznhzgl9ab2i_x2bpo1bvzos = hy_qezp81icfs3e8q66_zj ? d5jrixpw82rcyxb77lqvpjt : pn2h5gfpc4kw0y66t9;
  assign l9x1ubg9wznb6ixv1i  = (jbuu2xdq0qw_wi19r == ytx4fsx0_lffvqrj) & (~(ofznhzgl9ab2i_x2bpo1bvzos == r5bo9n9q6a8c5e5mv29k6wr));

  assign z2s7c4x2upx2k94 = ~tlwo81ky1a6b8;

  wire rwsuwy1bu82silyha06rggrf;
  wire rkpp17fj9tfksrejydcwru1;

  ux607_gnrl_fifo # (
   .CUT_READY(0),
   .DP(qrt6p0l7zsi7heuq),
   .DW(ynlkel_xoan9ow)
  ) oxeuy_ujjxzsn1i_ptt3rckm3frq (
   .i_vld(rwsuwy1bu82silyha06rggrf),
   .i_rdy(), 
   .i_dat(nc91g6pv91sa5ofkv6oqrzywy),
   .o_vld(), 
   .o_rdy(rkpp17fj9tfksrejydcwru1), 
   .o_dat(p738fnhowqrqokqjpa0a748b),

   .clk  (gf33atgy  ),
   .rst_n(ru_wi)  
  );

  wire ica3vfgm5bata1asuow;
  wire n_0k_24nqbeq5go0i17i;

  ux607_gnrl_fifo # (
   .CUT_READY(0),
   .DP(qrt6p0l7zsi7heuq),
   .DW(ynlkel_xoan9ow)
  ) zz64t3zdn7gcdp_b41b__5wfely (
   .i_vld(ica3vfgm5bata1asuow),
   .i_rdy(), 
   .i_dat(pwi4opocymgcqmwe_vq4sm0),
   .o_vld(), 
   .o_rdy(n_0k_24nqbeq5go0i17i), 
   .o_dat(tq4o19u3oc43c2v2sc9hsityj),

   .clk  (gf33atgy  ),
   .rst_n(ru_wi)  
  );

  wire mvud0s01b7n5fysigki_efg3zysp4bk1lts;
  wire p11an_iatsqmyhotqeai;
  wire fwlog0iiy2aq1zwy865vg9mu;

  ux607_gnrl_fifo # (
   .CUT_READY(0),
   .DP(qrt6p0l7zsi7heuq),
   .DW(ynlkel_xoan9ow)
  ) axemvggs77p4nuq3ztdby0lpni1t4 (
   .i_vld(mvud0s01b7n5fysigki_efg3zysp4bk1lts),
   .i_rdy(), 
   .i_dat(pne0i0g6_hms5_ag22zyfpdmpf3),
   .o_vld(), 
   .o_rdy(fwlog0iiy2aq1zwy865vg9mu), 
   .o_dat(vk3aoj6halc2m4mdlurcg7joxd),
 
   .clk  (gf33atgy  ),
   .rst_n(ru_wi)  
  );

        
  wire lidm0bbo5jcorhwlodeg2t = ((xpd4oma8mrw21r9b0mc8c | ytx0p13ahjuk751e8crl_0) & (~ghikvq604upn2v)) | ohprpkw231g_f2qqzmq;

  wire                          k6uqslf4yjz0;
  wire [3-1:0]   ibegorpv3fon9ktf; 

  genvar i;
  generate 
      for (i=0; i<yvxy18k82q; i=i+1) begin:filydm41n5gf3jyfic

        assign kyu0c7rbs3tzasd[i] = wf8kpn_u83u2_gj9bsb & (gtbu9zcij35aw_0ph1j == i[3-1:0]);
        assign m64tp4jpwoadr8w[i] = p_hc6rswvpztv26i & (fnvtppgr2s0i78 == i[3-1:0]);
        assign x5p4oi1vgjp37abo6[i] = kyu0c7rbs3tzasd[i] | m64tp4jpwoadr8w[i];
        assign iexhykoj1n453[i] = kyu0c7rbs3tzasd[i];

        ux607_gnrl_dfflr #(1) jo7q74300uyjp8gq3 (x5p4oi1vgjp37abo6[i], iexhykoj1n453[i], g53evua7d3gpxw3[i], gf33atgy, ru_wi);

          assign welnckam1xqornvo_[i][0] = kyu0c7rbs3tzasd[i] 
                                          & g53evua7d3gpxw3[0] & (~n7nx9bfxwcqwv7[0])
                                          & (


                                              (g2x5gi27ly4aw24 & dmjcrnz0ai9_04[0])
                                              | 
                                              ( 

                                                   (vx_fynrmojs7gx ^ qp1mbsaizjipsj6[0]) & 


                                                   (hdwldkfk3vetnqg3us[32-1:3] == haaqh6wjlwi9jhnl[0][32-1:3])
                                              )
                                            )
                                            & (~pup241nwugqoxaddw6o[0])
                                          ;
          assign j23uvqn5e9vkkw0w2fht[i][0] = b2rl4ox_6rp8po4j2tz[i][0] & pup241nwugqoxaddw6o[0];
          assign pnedptzdy93p4krxqb_p[i][0] = welnckam1xqornvo_[i][0] | j23uvqn5e9vkkw0w2fht[i][0];
          assign b700gcu8o4ko92g1i7kcc[i][0] = welnckam1xqornvo_[i][0];
        ux607_gnrl_dfflr #(1) eeyfqt3ks9t8f8f0_dfflr (pnedptzdy93p4krxqb_p[i][0], b700gcu8o4ko92g1i7kcc[i][0], b2rl4ox_6rp8po4j2tz[i][0], gf33atgy, ru_wi);
          assign welnckam1xqornvo_[i][1] = kyu0c7rbs3tzasd[i] 
                                          & g53evua7d3gpxw3[1] & (~n7nx9bfxwcqwv7[1])
                                          & (


                                              (g2x5gi27ly4aw24 & dmjcrnz0ai9_04[1])
                                              | 
                                              ( 

                                                   (vx_fynrmojs7gx ^ qp1mbsaizjipsj6[1]) & 


                                                   (hdwldkfk3vetnqg3us[32-1:3] == haaqh6wjlwi9jhnl[1][32-1:3])
                                              )
                                            )
                                            & (~pup241nwugqoxaddw6o[1])
                                          ;
          assign j23uvqn5e9vkkw0w2fht[i][1] = b2rl4ox_6rp8po4j2tz[i][1] & pup241nwugqoxaddw6o[1];
          assign pnedptzdy93p4krxqb_p[i][1] = welnckam1xqornvo_[i][1] | j23uvqn5e9vkkw0w2fht[i][1];
          assign b700gcu8o4ko92g1i7kcc[i][1] = welnckam1xqornvo_[i][1];
        ux607_gnrl_dfflr #(1) eeyfqt3ks9t8f8f1_dfflr (pnedptzdy93p4krxqb_p[i][1], b700gcu8o4ko92g1i7kcc[i][1], b2rl4ox_6rp8po4j2tz[i][1], gf33atgy, ru_wi);
          assign welnckam1xqornvo_[i][2] = kyu0c7rbs3tzasd[i] 
                                          & g53evua7d3gpxw3[2] & (~n7nx9bfxwcqwv7[2])
                                          & (


                                              (g2x5gi27ly4aw24 & dmjcrnz0ai9_04[2])
                                              | 
                                              ( 

                                                   (vx_fynrmojs7gx ^ qp1mbsaizjipsj6[2]) & 


                                                   (hdwldkfk3vetnqg3us[32-1:3] == haaqh6wjlwi9jhnl[2][32-1:3])
                                              )
                                            )
                                            & (~pup241nwugqoxaddw6o[2])
                                          ;
          assign j23uvqn5e9vkkw0w2fht[i][2] = b2rl4ox_6rp8po4j2tz[i][2] & pup241nwugqoxaddw6o[2];
          assign pnedptzdy93p4krxqb_p[i][2] = welnckam1xqornvo_[i][2] | j23uvqn5e9vkkw0w2fht[i][2];
          assign b700gcu8o4ko92g1i7kcc[i][2] = welnckam1xqornvo_[i][2];
        ux607_gnrl_dfflr #(1) eeyfqt3ks9t8f8f2_dfflr (pnedptzdy93p4krxqb_p[i][2], b700gcu8o4ko92g1i7kcc[i][2], b2rl4ox_6rp8po4j2tz[i][2], gf33atgy, ru_wi);
          assign welnckam1xqornvo_[i][3] = kyu0c7rbs3tzasd[i] 
                                          & g53evua7d3gpxw3[3] & (~n7nx9bfxwcqwv7[3])
                                          & (


                                              (g2x5gi27ly4aw24 & dmjcrnz0ai9_04[3])
                                              | 
                                              ( 

                                                   (vx_fynrmojs7gx ^ qp1mbsaizjipsj6[3]) & 


                                                   (hdwldkfk3vetnqg3us[32-1:3] == haaqh6wjlwi9jhnl[3][32-1:3])
                                              )
                                            )
                                            & (~pup241nwugqoxaddw6o[3])
                                          ;
          assign j23uvqn5e9vkkw0w2fht[i][3] = b2rl4ox_6rp8po4j2tz[i][3] & pup241nwugqoxaddw6o[3];
          assign pnedptzdy93p4krxqb_p[i][3] = welnckam1xqornvo_[i][3] | j23uvqn5e9vkkw0w2fht[i][3];
          assign b700gcu8o4ko92g1i7kcc[i][3] = welnckam1xqornvo_[i][3];
        ux607_gnrl_dfflr #(1) eeyfqt3ks9t8f8f3_dfflr (pnedptzdy93p4krxqb_p[i][3], b700gcu8o4ko92g1i7kcc[i][3], b2rl4ox_6rp8po4j2tz[i][3], gf33atgy, ru_wi);
          assign welnckam1xqornvo_[i][4] = kyu0c7rbs3tzasd[i] 
                                          & g53evua7d3gpxw3[4] & (~n7nx9bfxwcqwv7[4])
                                          & (


                                              (g2x5gi27ly4aw24 & dmjcrnz0ai9_04[4])
                                              | 
                                              ( 

                                                   (vx_fynrmojs7gx ^ qp1mbsaizjipsj6[4]) & 


                                                   (hdwldkfk3vetnqg3us[32-1:3] == haaqh6wjlwi9jhnl[4][32-1:3])
                                              )
                                            )
                                            & (~pup241nwugqoxaddw6o[4])
                                          ;
          assign j23uvqn5e9vkkw0w2fht[i][4] = b2rl4ox_6rp8po4j2tz[i][4] & pup241nwugqoxaddw6o[4];
          assign pnedptzdy93p4krxqb_p[i][4] = welnckam1xqornvo_[i][4] | j23uvqn5e9vkkw0w2fht[i][4];
          assign b700gcu8o4ko92g1i7kcc[i][4] = welnckam1xqornvo_[i][4];
        ux607_gnrl_dfflr #(1) eeyfqt3ks9t8f8f4_dfflr (pnedptzdy93p4krxqb_p[i][4], b700gcu8o4ko92g1i7kcc[i][4], b2rl4ox_6rp8po4j2tz[i][4], gf33atgy, ru_wi);
          assign welnckam1xqornvo_[i][5] = kyu0c7rbs3tzasd[i] 
                                          & g53evua7d3gpxw3[5] & (~n7nx9bfxwcqwv7[5])
                                          & (


                                              (g2x5gi27ly4aw24 & dmjcrnz0ai9_04[5])
                                              | 
                                              ( 

                                                   (vx_fynrmojs7gx ^ qp1mbsaizjipsj6[5]) & 


                                                   (hdwldkfk3vetnqg3us[32-1:3] == haaqh6wjlwi9jhnl[5][32-1:3])
                                              )
                                            )
                                            & (~pup241nwugqoxaddw6o[5])
                                          ;
          assign j23uvqn5e9vkkw0w2fht[i][5] = b2rl4ox_6rp8po4j2tz[i][5] & pup241nwugqoxaddw6o[5];
          assign pnedptzdy93p4krxqb_p[i][5] = welnckam1xqornvo_[i][5] | j23uvqn5e9vkkw0w2fht[i][5];
          assign b700gcu8o4ko92g1i7kcc[i][5] = welnckam1xqornvo_[i][5];
        ux607_gnrl_dfflr #(1) eeyfqt3ks9t8f8f5_dfflr (pnedptzdy93p4krxqb_p[i][5], b700gcu8o4ko92g1i7kcc[i][5], b2rl4ox_6rp8po4j2tz[i][5], gf33atgy, ru_wi);
          assign welnckam1xqornvo_[i][6] = kyu0c7rbs3tzasd[i] 
                                          & g53evua7d3gpxw3[6] & (~n7nx9bfxwcqwv7[6])
                                          & (


                                              (g2x5gi27ly4aw24 & dmjcrnz0ai9_04[6])
                                              | 
                                              ( 

                                                   (vx_fynrmojs7gx ^ qp1mbsaizjipsj6[6]) & 


                                                   (hdwldkfk3vetnqg3us[32-1:3] == haaqh6wjlwi9jhnl[6][32-1:3])
                                              )
                                            )
                                            & (~pup241nwugqoxaddw6o[6])
                                          ;
          assign j23uvqn5e9vkkw0w2fht[i][6] = b2rl4ox_6rp8po4j2tz[i][6] & pup241nwugqoxaddw6o[6];
          assign pnedptzdy93p4krxqb_p[i][6] = welnckam1xqornvo_[i][6] | j23uvqn5e9vkkw0w2fht[i][6];
          assign b700gcu8o4ko92g1i7kcc[i][6] = welnckam1xqornvo_[i][6];
        ux607_gnrl_dfflr #(1) eeyfqt3ks9t8f8f6_dfflr (pnedptzdy93p4krxqb_p[i][6], b700gcu8o4ko92g1i7kcc[i][6], b2rl4ox_6rp8po4j2tz[i][6], gf33atgy, ru_wi);
          assign welnckam1xqornvo_[i][7] = kyu0c7rbs3tzasd[i] 
                                          & g53evua7d3gpxw3[7] & (~n7nx9bfxwcqwv7[7])
                                          & (


                                              (g2x5gi27ly4aw24 & dmjcrnz0ai9_04[7])
                                              | 
                                              ( 

                                                   (vx_fynrmojs7gx ^ qp1mbsaizjipsj6[7]) & 


                                                   (hdwldkfk3vetnqg3us[32-1:3] == haaqh6wjlwi9jhnl[7][32-1:3])
                                              )
                                            )
                                            & (~pup241nwugqoxaddw6o[7])
                                          ;
          assign j23uvqn5e9vkkw0w2fht[i][7] = b2rl4ox_6rp8po4j2tz[i][7] & pup241nwugqoxaddw6o[7];
          assign pnedptzdy93p4krxqb_p[i][7] = welnckam1xqornvo_[i][7] | j23uvqn5e9vkkw0w2fht[i][7];
          assign b700gcu8o4ko92g1i7kcc[i][7] = welnckam1xqornvo_[i][7];
        ux607_gnrl_dfflr #(1) eeyfqt3ks9t8f8f7_dfflr (pnedptzdy93p4krxqb_p[i][7], b700gcu8o4ko92g1i7kcc[i][7], b2rl4ox_6rp8po4j2tz[i][7], gf33atgy, ru_wi);


        assign puxm_ue7jwuwh72gi[i] = x5p4oi1vgjp37abo6[i] ? iexhykoj1n453[i] : g53evua7d3gpxw3[i];


        assign mnch_edao2_c4_ni2[i] = kyu0c7rbs3tzasd[i];
        assign ttgsuta_ewmr6[i] = (w3ss3ti2t0dj2tvx & (jgfckxgs0fo048 == i[3-1:0])); 
        assign ny0n30vi0dzifq_o[i] = mnch_edao2_c4_ni2[i] | ttgsuta_ewmr6[i];
        assign cgst_q5rcj_eo2wfk[i] = mnch_edao2_c4_ni2[i];

        ux607_gnrl_dfflr #(1) ttzwehxbic556a_d7k (ny0n30vi0dzifq_o[i], cgst_q5rcj_eo2wfk[i], n3k7lk4c5q[i], gf33atgy, ru_wi);

        assign ttgaf1h84fzp0d1oel7[i] = (f__yd2_rd0i7mgsj05bn[i] | buxvgnamnlcw3lpbel0[i] 
                                                  | d763qyon3q45pdbxztuo4[i]  
                                                );
        assign pup241nwugqoxaddw6o[i] = m64tp4jpwoadr8w[i];
        assign j6x4yktmu5u6_uil[i] = ttgaf1h84fzp0d1oel7[i] | pup241nwugqoxaddw6o[i];
        assign o8btl8op6tng90p0h[i] = ttgaf1h84fzp0d1oel7[i];

        ux607_gnrl_dfflr #(1) hctuzh67uuch1pgax5 (j6x4yktmu5u6_uil[i], o8btl8op6tng90p0h[i], n7nx9bfxwcqwv7[i], gf33atgy, ru_wi);

        assign mwvgay3ta4a2[i] = k23tmhod3m0plvdlp & (s8ol0xfe2arkosb == i[3-1:0]);
        assign os4b0yseamo1t[i] = m64tp4jpwoadr8w[i];
        assign brv_ewhw27bxxr_[i] = mwvgay3ta4a2[i] | os4b0yseamo1t[i];
        assign rkx1mrv8yqxi8el[i] = (~os4b0yseamo1t[i]);

        ux607_gnrl_dfflr #(1) bliew68hvg4vlv (brv_ewhw27bxxr_[i], rkx1mrv8yqxi8el[i], a672uxn3mwn[i], gf33atgy, ru_wi);

        assign g7qqd7ejlmjzz7uab[i] = kyu0c7rbs3tzasd[i] & lidm0bbo5jcorhwlodeg2t; 
        assign tg8y2zr5rfj4sw1xke8[i] = (k6uqslf4yjz0 & (ibegorpv3fon9ktf == i[3-1:0]));
        assign vkzm86ii21rro827o0[i] = g7qqd7ejlmjzz7uab[i] | tg8y2zr5rfj4sw1xke8[i];
        assign oosv_ui3yrxrqb_nh89[i] = g7qqd7ejlmjzz7uab[i];
  
        ux607_gnrl_dfflr #(1) b23grdf9umzw5pvfrk (vkzm86ii21rro827o0[i], oosv_ui3yrxrqb_nh89[i], l_ldkrkpn59v4mhb_[i], gf33atgy, ru_wi); 





        assign rg7cda_918ahdww6p56mv81qg_[i] = v1bfb0aqght1_yfm5znt[i] & (~pllepw4azlfujoh_i[i]);

        assign a2oenic4uandesr_k9qocfw[i] = g53evua7d3gpxw3[i] & (~rg7cda_918ahdww6p56mv81qg_[i]) & (~knyt1bhi0tp16v3[i]);

        assign ixtmkj78nheu_ghv7byt0w[i] = g53evua7d3gpxw3[i] & (
                                      w8u6pj2octqg9n0vi6[i]
                                    );

        assign fa8x97zn7g9lhjdunyuqg[i] = puxm_ue7jwuwh72gi[i] & (
                                      ea8x6ufv3q0voque2u5o8[i]
                                    );


        assign e0umr420ntwlczrjba[i] = g53evua7d3gpxw3[i] & n3k7lk4c5q[i]
                                     & (~(|b2rl4ox_6rp8po4j2tz[i]))
                                     ;

        assign d7roxn5jsm8p278tf[i] = g53evua7d3gpxw3[i] & (~a672uxn3mwn[i]) & (a2oenic4uandesr_k9qocfw[i] ? n7nx9bfxwcqwv7[i] : 1'b1) & (~ixtmkj78nheu_ghv7byt0w[i]);

        assign y206os9wqkqs1a7zyv[i] = g53evua7d3gpxw3[i] & (~n3k7lk4c5q[i])  & (a672uxn3mwn[i] | mwvgay3ta4a2[i])  & (a2oenic4uandesr_k9qocfw[i] ? n7nx9bfxwcqwv7[i] : 1'b1 ) 
                                   & (~l_ldkrkpn59v4mhb_[i])  
                                   ;


        ux607_gnrl_dfflr #(32) mff371e7jrp6xy2kf        (kyu0c7rbs3tzasd[i], hdwldkfk3vetnqg3us    , haaqh6wjlwi9jhnl[i]    , gf33atgy, ru_wi);
        ux607_gnrl_dfflr #(              1) fpc3o8kyopchwataqd26m8y  (kyu0c7rbs3tzasd[i], kix9_o92mst68vescu79v, w8u6pj2octqg9n0vi6[i]   , gf33atgy, ru_wi);
        ux607_gnrl_dfflr #(              1) h5y3th04w9g6n6pfpk2w8tlycgx(kyu0c7rbs3tzasd[i], lidm0bbo5jcorhwlodeg2t, v84iwz704r1326150y[i]   , gf33atgy, ru_wi);
        ux607_gnrl_dfflr #(              1) xwc6j4xipx7zwusa9m       (kyu0c7rbs3tzasd[i], ihkz9tebg3jd5f47z   , xzc0imuvetgbn8[i]   , gf33atgy, ru_wi);
        ux607_gnrl_dfflr #(              1) osyiapt643wo2u9l83hq       (kyu0c7rbs3tzasd[i], tu1v8ryo2rv95crsvz   , halyb9c30hal[i]   , gf33atgy, ru_wi);
        ux607_gnrl_dfflr #(              1) ansd5452q3j9yoioodd3c       (kyu0c7rbs3tzasd[i], ghikvq604upn2v   , pllepw4azlfujoh_i[i]   , gf33atgy, ru_wi);
        ux607_gnrl_dfflr #(              1) ec2fhj42e0_595ilw8ph_yes  (kyu0c7rbs3tzasd[i], t4leke6w3uzo3gxu3yhk   , d1rzzdht0dlkdfjvs420q[i]   , gf33atgy, ru_wi);
        ux607_gnrl_dfflr #(              1) nbl_y00g5syozwfapc7s_  (kyu0c7rbs3tzasd[i], oodqv7hv99boddj3kk48j   , hwwn5fuw1ki6rpxis[i]   , gf33atgy, ru_wi);
        ux607_gnrl_dfflr #(              1) r2fn9h5s8ufgqk08tu      (kyu0c7rbs3tzasd[i], g2x5gi27ly4aw24  , dmjcrnz0ai9_04[i]  , gf33atgy, ru_wi);
        ux607_gnrl_dfflr #(              1) t8pozfv3tulwroc          (kyu0c7rbs3tzasd[i], g16len3w2wk22u      , t54w0z3ee_q[i]      , gf33atgy, ru_wi);
        ux607_gnrl_dfflr #(              1) ibf2pe731u9m4ypy4j        (kyu0c7rbs3tzasd[i], vx_fynrmojs7gx    , qp1mbsaizjipsj6[i]    , gf33atgy, ru_wi);
        ux607_gnrl_dfflr #(              1) z82u8p8s8s3a2x_k0nrsa53b  (kyu0c7rbs3tzasd[i], ytx0p13ahjuk751e8crl_0, v1bfb0aqght1_yfm5znt[i], gf33atgy, ru_wi);
        ux607_gnrl_dfflr #(              1) pq62u9k16z_6dgspya60eb_   (kyu0c7rbs3tzasd[i], xpd4oma8mrw21r9b0mc8c, cuslzq6_3njc_9dr[i], gf33atgy, ru_wi);
        ux607_gnrl_dfflr #(8   ) xazi9t8l7j3pcrhbkygr       (kyu0c7rbs3tzasd[i], v0uq3fcdfb8eatt3   , zrhld0y35qav[i]   , gf33atgy, ru_wi);
        ux607_gnrl_dfflr #(              1) c7n7gm06n57jim8r1d        (kyu0c7rbs3tzasd[i], c4otadutq6rav14ed2    , epo0qysbvw4gkmi[i]    , gf33atgy, ru_wi);
        ux607_gnrl_dfflr #(              1) zb1etj2bs_m7pgmcq1ky        (kyu0c7rbs3tzasd[i], mw8uaelv0i5zfav    , c274s6asp6_ptv[i]    , gf33atgy, ru_wi);
        ux607_gnrl_dfflr #(              2) m3ghcb2zi5xdumhrh        (kyu0c7rbs3tzasd[i], uq0oocqz_ys0no4o_t    , bx9szwl63ur[i]    , gf33atgy, ru_wi);
        ux607_gnrl_dfflr #(              1) w6ymwa79qgeczx2cyoz0zk9    (kyu0c7rbs3tzasd[i], ohprpkw231g_f2qqzmq, knyt1bhi0tp16v3[i], gf33atgy, ru_wi);
        ux607_gnrl_dfflr #(              1) ccj3a_yjcxh5930v3tmzx54hyan    (kyu0c7rbs3tzasd[i], e3l8n6__k56uw5o7jujwibr, fizjb37qgnqc11y3usvo1jd8[i], gf33atgy, ru_wi);
        ux607_gnrl_dfflr #(              1) klzm1myvh7p8_ru5qio_uu3_jp7    (kyu0c7rbs3tzasd[i], rwmac6nity_ikz7xbj_ta1nce, te3sgyqybgiz02r496eiram[i], gf33atgy, ru_wi);
        ux607_gnrl_dfflr #(              1) zhzi5ja7x0xy8b8enfgmd2yvz1    (kyu0c7rbs3tzasd[i], en9ogfq6nx_uirma3y2jiigbh, hotgsfmzxnfg6u691gfcuem[i], gf33atgy, ru_wi);
        ux607_gnrl_dfflr #(              1) gs27edv_5la14fjjtpla2hz7k3    (kyu0c7rbs3tzasd[i], t9otq6y33fc5qs21p9d2rc3zn, dej8khi216rqhe3ebb4[i], gf33atgy, ru_wi);
        ux607_gnrl_dfflr #(              1) baxbr0x6sx7c4_8aiiuspg    (kyu0c7rbs3tzasd[i], xpbzeko14yty79dehft9e2l, bk8m_k0vayvzu1ytxtuvky[i], gf33atgy, ru_wi);

        assign c3mjay1nkztzsfo3mf2[i]      = kyu0c7rbs3tzasd[i] ? ytx0p13ahjuk751e8crl_0      : v1bfb0aqght1_yfm5znt     [i];
        assign di2o65qovx5zvsf3rujmc[i]        = kyu0c7rbs3tzasd[i] ? ohprpkw231g_f2qqzmq        : knyt1bhi0tp16v3       [i];
        assign ea8x6ufv3q0voque2u5o8[i]      = kyu0c7rbs3tzasd[i] ? kix9_o92mst68vescu79v      : w8u6pj2octqg9n0vi6     [i];


        assign f__yd2_rd0i7mgsj05bn[i]  = rkpp17fj9tfksrejydcwru1 & (p738fnhowqrqokqjpa0a748b == i[3-1:0]); 
        assign buxvgnamnlcw3lpbel0[i]  = n_0k_24nqbeq5go0i17i & (tq4o19u3oc43c2v2sc9hsityj == i[3-1:0]); 
        assign d763qyon3q45pdbxztuo4[i] = fwlog0iiy2aq1zwy865vg9mu & (vk3aoj6halc2m4mdlurcg7joxd == i[3-1:0]); 

        assign {asf2z47ldhqkwm15lbpzc[i], kcgdolb8q4gs6fitbr3v_[i], ypal30idlttlfu9s_qrvo[i] }     = (
                               ({64+2{f__yd2_rd0i7mgsj05bn[i] }} & {ng9lxc1zr1snbj1p1b9 , nykvnvl0i96asmogcmhlrpy , b_7_y71ywtomguvgnoq5 }) 
                             | ({64+2{buxvgnamnlcw3lpbel0[i] }} & {g5a675dzhov32an3m , efz5oj5hqaeq_wptcenc10fq7 , bhhfkcv51hmdpdenvztypn })
                             | ({64+2{d763qyon3q45pdbxztuo4[i]}} & {gl9dazcghkmei56i8tlb, k7x2rdsdsxkmoiyluje7bf2aa, j1utgrdwzlhqppb8rev5pbh55})
                 );


        ux607_gnrl_dfflr #(1) br9k93zt31tzcac6bf23_     (ttgaf1h84fzp0d1oel7[i], asf2z47ldhqkwm15lbpzc[i]    , xezq29zs58h59dv[i]    , gf33atgy, ru_wi);
        ux607_gnrl_dfflr #(1) mpeybvah3z0_lm2b52c5ity (ttgaf1h84fzp0d1oel7[i], kcgdolb8q4gs6fitbr3v_[i], hmqlykdc12wo5_r73zg8[i], gf33atgy, ru_wi);

        assign u5zzpdddo7nx53kgpobe[i] = qp1mbsaizjipsj6[i] & ttgaf1h84fzp0d1oel7[i];
        assign ckambm7sahfb9bg1nm[i] = (kyu0c7rbs3tzasd[i] & (~vx_fynrmojs7gx)); 

        assign i801bchffjgm2eeav1c0[i] = ckambm7sahfb9bg1nm[i] 
                                     | u5zzpdddo7nx53kgpobe[i]; 

        assign b9i1i44zz7lsiekhgww[i] = u5zzpdddo7nx53kgpobe[i] ? ypal30idlttlfu9s_qrvo[i] : uacpumgrbwt0fmb;

        ux607_gnrl_dfflr #(64) ifckjvpl4sc3th1gfl (i801bchffjgm2eeav1c0[i], b9i1i44zz7lsiekhgww[i], vsfpyprm4rivny0n4[i], gf33atgy, ru_wi);

        assign zlgnht9uo2fb7p[i]  = (v1bfb0aqght1_yfm5znt[i] | cuslzq6_3njc_9dr[i]) & g53evua7d3gpxw3[i] & 
                       (z8alxhlwgz117[32-1:5] == haaqh6wjlwi9jhnl[i][32-1:5]);
        assign yel5kfjrg5ib6[i]  = (v1bfb0aqght1_yfm5znt[i] | cuslzq6_3njc_9dr[i]) & g53evua7d3gpxw3[i] & 
                       (q4j831gvqooep12[32-1:5] == haaqh6wjlwi9jhnl[i][32-1:5]);
      end
  endgenerate

  assign y5otpn351odm3mnpnfdshm = ~(| (g53evua7d3gpxw3 & (~ixtmkj78nheu_ghv7byt0w)));
  assign rnlnwebfnqcg8g5oq_2gv0 = ~(| (puxm_ue7jwuwh72gi & (~fa8x97zn7g9lhjdunyuqg)));

  wire nl2n_jy0ye9rq9j0hteu;
  wire bvwt0k4qftqv4to2lj6d46_;
  wire xerurm1znxab6ednf5rf;
  wire ocz7civlapwkb3oe78oqt2fw;

  assign yafkacaefbdmi3hm6rvuao = (| zlgnht9uo2fb7p) | nl2n_jy0ye9rq9j0hteu | bvwt0k4qftqv4to2lj6d46_;
  assign u4frf_hcy8c0dh_aqkgsrp = (| yel5kfjrg5ib6) | xerurm1znxab6ednf5rf | ocz7civlapwkb3oe78oqt2fw;

  assign pwi4opocymgcqmwe_vq4sm0  = jgfckxgs0fo048; 
  assign nc91g6pv91sa5ofkv6oqrzywy  = jgfckxgs0fo048; 
  assign pne0i0g6_hms5_ag22zyfpdmpf3 = jgfckxgs0fo048; 

  wire b2b_rqtoetzhmz2za = qp1mbsaizjipsj6[jgfckxgs0fo048];
  wire as6c9asy2pmyim1mpl6 = knyt1bhi0tp16v3[jgfckxgs0fo048];
  wire nhhkvz0vlgwkhroehttknd4 = fizjb37qgnqc11y3usvo1jd8[jgfckxgs0fo048];
  wire vvszajn57xalwihwqb10 = te3sgyqybgiz02r496eiram[jgfckxgs0fo048];
  wire fs6va8zhb7c7up7raca6re8y_4 = hotgsfmzxnfg6u691gfcuem[jgfckxgs0fo048];
  wire za44bo8vauicq1_d2xn8u9xau = dej8khi216rqhe3ebb4[jgfckxgs0fo048];
  wire ymqea1d98jlrnw9zubeo = bk8m_k0vayvzu1ytxtuvky[jgfckxgs0fo048];

  wire ot8jvy0c6kgqefqv = ~(v84iwz704r1326150y[jgfckxgs0fo048]);
  wire bfr5u4s_wl1y3qg = ot8jvy0c6kgqefqv & b2b_rqtoetzhmz2za;  
  wire dpkcph27_2sm8d0l = ot8jvy0c6kgqefqv & (~b2b_rqtoetzhmz2za);   
  wire aoooi7kgel8pjm = ~ot8jvy0c6kgqefqv;

  assign zfu2vonacwweg65jwl5h  = blwju8dk7oqctm5 & bfr5u4s_wl1y3qg;
  assign ejbq7zgkpgwgttfvvx5rp  = blwju8dk7oqctm5 & dpkcph27_2sm8d0l;
  assign zsp7u2uqvojc8zqnw0k6_p = blwju8dk7oqctm5 & aoooi7kgel8pjm;

  assign tm4v0w70xpfbnl8980 = (
                            (ecc0pa6dsujd5fk_ztk1odty  & bfr5u4s_wl1y3qg)
                          | (agtve46c928tzy8367oy14bf  & dpkcph27_2sm8d0l)
                          | (mljh30sszwrhguqyc4f5e77l4 & aoooi7kgel8pjm)
              );


  assign i0znoodcvzhh4rexar7joqvk = 1'b1;
  assign q2_zn_ozuoxddlj2se_t45w = 1'b1;
  assign vydbpbb7_kmw71ncfvuvj74 = 1'b1;

  assign ica3vfgm5bata1asuow = zfu2vonacwweg65jwl5h & ecc0pa6dsujd5fk_ztk1odty;
  assign rwsuwy1bu82silyha06rggrf = ejbq7zgkpgwgttfvvx5rp & agtve46c928tzy8367oy14bf;
  wire   fegv040vs2cbidgh74h_gtkeg;
  assign p11an_iatsqmyhotqeai = zsp7u2uqvojc8zqnw0k6_p & mljh30sszwrhguqyc4f5e77l4;
  assign mvud0s01b7n5fysigki_efg3zysp4bk1lts = p11an_iatsqmyhotqeai & fegv040vs2cbidgh74h_gtkeg;

  assign n_0k_24nqbeq5go0i17i = z9q40jbnm38zcodsjsd090z & i0znoodcvzhh4rexar7joqvk;
  assign rkpp17fj9tfksrejydcwru1 = gcan4qd32d7splx9secvc8b & q2_zn_ozuoxddlj2se_t45w;
  assign fwlog0iiy2aq1zwy865vg9mu = yp6atu2uzbb053onf7h7j_g3 & vydbpbb7_kmw71ncfvuvj74;

  assign p2m0mydv1zb_6iqetg5 = 1'b1; 
  assign m6vmtqf14m_q0ahhpf9ys0t = 1'b0; 

  assign a01toa5fu8pmct9z1qeb  = 64'b0;
  assign ex_5rp8vtq6iwx6hm_w  = 8'b0;

  assign hn4lhm3a_wcnqbxq84q  = vsfpyprm4rivny0n4 [jgfckxgs0fo048];
  assign pqhi5t7t91o9xtpy8r4_9o  = zrhld0y35qav [jgfckxgs0fo048];

  assign t60xfh0jvayj7nnp_3swk1v   = haaqh6wjlwi9jhnl  [jgfckxgs0fo048]; 
  assign m_zge7ydxw1me0bp66_b  = 3'b0;
  assign vo4iscd43mm129ts9g7   = 2'b0;
  assign n5ajmphmp207ybl3ru6ee3p   = epo0qysbvw4gkmi  [jgfckxgs0fo048];
  assign r_te1f8papt089n46s6j2k   = c274s6asp6_ptv  [jgfckxgs0fo048];
  assign ao8xdzkmlvr9h6inuey9k   = bx9szwl63ur  [jgfckxgs0fo048];
  assign b6c9ysz1s8lqf83mno84  = xzc0imuvetgbn8 [jgfckxgs0fo048]; 
  assign gam1zdrkynr0puyhapwkq5fs  = halyb9c30hal [jgfckxgs0fo048]; 
  assign w_bo91bpxaukiy9s3fyc9ib6  = pllepw4azlfujoh_i [jgfckxgs0fo048]; 
  assign yivyo1xc3okylkdzlkar = dmjcrnz0ai9_04[jgfckxgs0fo048]; 
  assign acdtgtj2r5zy7qoh9ukv     = t54w0z3ee_q    [jgfckxgs0fo048]; 
  assign fegv040vs2cbidgh74h_gtkeg     = a2oenic4uandesr_k9qocfw[jgfckxgs0fo048]; 

  assign pii5a6cmz40r9w30q_awu   = t60xfh0jvayj7nnp_3swk1v  ; 
  assign zhc7g2_tfy2pqp2f8g5  = m_zge7ydxw1me0bp66_b ;
  assign edt_9_yofk03w8y7jt   = vo4iscd43mm129ts9g7  ;
  assign zeqnplthuo3przg6v7sc   = n5ajmphmp207ybl3ru6ee3p  ;
  assign ia_e66cu_no6wwvfzv   = r_te1f8papt089n46s6j2k  ;
  assign ceg6dnmky0mxytf2e9bhe0   = ao8xdzkmlvr9h6inuey9k  ;
  assign x934mbk53lq9pp23th7n5no0  = b6c9ysz1s8lqf83mno84 ; 
  assign qw8c56hyyf3o9z35eb8m  = gam1zdrkynr0puyhapwkq5fs ; 
  assign tpkr0onb62gbg0ddt7_pz4l  = w_bo91bpxaukiy9s3fyc9ib6 ; 
  assign j_e7kc3w9drko64cvqn5g = yivyo1xc3okylkdzlkar; 
  assign fz8l_vym0or20pcgjct     = acdtgtj2r5zy7qoh9ukv    ; 


  assign huqvm9m1hvosa8sc4xjt  = ixtmkj78nheu_ghv7byt0w[s8ol0xfe2arkosb] & (~a672uxn3mwn[s8ol0xfe2arkosb]);
  wire   kxncstfuoj9lu6kva4j = a2oenic4uandesr_k9qocfw[s8ol0xfe2arkosb];

  assign blwju8dk7oqctm5 = e0umr420ntwlczrjba[jgfckxgs0fo048];
  assign r57mgw9ntmg26lxok = d7roxn5jsm8p278tf[s8ol0xfe2arkosb];

  assign ypuolenm4dvdg     = kxncstfuoj9lu6kva4j ? xezq29zs58h59dv    [s8ol0xfe2arkosb] : 1'b0;
  assign yu5m552dobcb8gbsq = kxncstfuoj9lu6kva4j ? hmqlykdc12wo5_r73zg8[s8ol0xfe2arkosb] : 1'b0;
  assign bo_q_t246zgg3q   = kxncstfuoj9lu6kva4j ? vsfpyprm4rivny0n4      [s8ol0xfe2arkosb] : 64'b0;
  assign d4k4iwwrjuzjqt    = haaqh6wjlwi9jhnl[s8ol0xfe2arkosb];

  assign xnmbaecrrzbadq6w = y206os9wqkqs1a7zyv[fnvtppgr2s0i78];

  localparam uw3hbdikblihw1_r3o = (32+1+64+8+3+2+1+1+2+5);
  localparam szbi56su117rxsuhhun = (1+1+64);

  wire [uw3hbdikblihw1_r3o-1:0] a23lzk9_jpf1wt6gpoa3t;
  wire [uw3hbdikblihw1_r3o-1:0] nzcpulhcv_r50wph3pz9;
  wire [szbi56su117rxsuhhun-1:0] kti_aenofx1syww4og3;
  wire [szbi56su117rxsuhhun-1:0] cmvo1gt96vee3wmg9e;

  assign 
       a23lzk9_jpf1wt6gpoa3t = { 
       t60xfh0jvayj7nnp_3swk1v, 
       p2m0mydv1zb_6iqetg5, 
       a01toa5fu8pmct9z1qeb,
       ex_5rp8vtq6iwx6hm_w,
       m_zge7ydxw1me0bp66_b,
       vo4iscd43mm129ts9g7,
       n5ajmphmp207ybl3ru6ee3p,
       r_te1f8papt089n46s6j2k,
       ao8xdzkmlvr9h6inuey9k,
       b6c9ysz1s8lqf83mno84, 
       gam1zdrkynr0puyhapwkq5fs, 
       w_bo91bpxaukiy9s3fyc9ib6, 
       yivyo1xc3okylkdzlkar, 
       acdtgtj2r5zy7qoh9ukv};

  assign 
       nzcpulhcv_r50wph3pz9 = { 
       pii5a6cmz40r9w30q_awu, 
       m6vmtqf14m_q0ahhpf9ys0t, 
       hn4lhm3a_wcnqbxq84q,
       pqhi5t7t91o9xtpy8r4_9o,
       zhc7g2_tfy2pqp2f8g5,
       edt_9_yofk03w8y7jt,
       zeqnplthuo3przg6v7sc,
       ia_e66cu_no6wwvfzv,
       ceg6dnmky0mxytf2e9bhe0,
       x934mbk53lq9pp23th7n5no0, 
       qw8c56hyyf3o9z35eb8m, 
       tpkr0onb62gbg0ddt7_pz4l, 
       j_e7kc3w9drko64cvqn5g, 
       fz8l_vym0or20pcgjct};

  assign {
                                    g5a675dzhov32an3m  ,
                                    efz5oj5hqaeq_wptcenc10fq7,
                                    bhhfkcv51hmdpdenvztypn} = kti_aenofx1syww4og3; 

  assign {
                                    ng9lxc1zr1snbj1p1b9  ,
                                    nykvnvl0i96asmogcmhlrpy,
                                    b_7_y71ywtomguvgnoq5} = cmvo1gt96vee3wmg9e; 


  
  
  
  
  
  
  
  
  
  
  
  
  
  wire                          bidjco9v6uwp91tvsqnp72df_u0q;
  wire                          m83gf40i8n5qmmo860pq3w7n5n5f;
  wire  [32-1:0]   q064m0tgrtkrz7vn_qf2bjb; 
  wire                          xxrb4v2suklf9djaeyf0rkmedjz3; 
  wire  [64-1:0]        hrn1giqg1k6gbt6q7lrxzxaqztx;
  wire  [8-1:0]     xw04i4vzqgn2m2ihbdv55m4bvtr;
  wire  [2:0]                   h_9b0wqhlkmvxkfizht97cqp;
  wire  [1:0]                   ycmo1kcbjq1scw4gwg4uiwd_;
  wire                          ocdu63ksnvvgacaermakucm0f4g;
  wire                          oxlxxz2rxp0amufq1s9jqrry3y;
  wire  [1:0]                   rcpyv929ixr6xhyeyg2p0cgtj;
  wire                          n169ohp8pq9l7goaugowzjfa; 
  wire                          psec5ihpqk4slg2u90eq4yzyy; 
  wire                          cv6960ns7f2dyrvj6ij_phb0; 
  wire                          kxqipwn8s_54dje1dpjvcgaye6t; 
  wire                          gc_aq81uy3hbdq8ns7y1_ckg; 

  wire                          vkjwr2hxue8911qmv5ro35cg;
  wire                          xronfobw50555i02avvye82b;
  wire  [32-1:0]   kbbc76s46hvu_3te0ihj3hb2nl; 
  wire                          g33u_ys44gmrebks2nd9y8o; 
  wire  [64-1:0]      y5gfh4gmog9i5iq47qq3nmc95_fnd;
  wire  [8-1:0]      bafx6nbdipfv60zavyhkpt5ulfqp;
  wire  [2:0]                   wfq3yog1gp3v5k8ew8aazeio5q9qm;
  wire  [1:0]                   bkec53bqczw0o6vx2ouxlbp;
  wire                          o347ncxtm6aeg09kb47k1oggzcw;
  wire                          pfkm_ekt4p23xk05wj0f5ei8wut2;
  wire  [1:0]                   rx7d01wkjl49umakx8rnira0bvj;
  wire                          bpetbkuwyy1k6fa142bfw3rz7sjpi; 
  wire                          vsn6zt6npfa5qvbab0qrm7ya; 
  wire                          c_saxxol2d2vxelssdxtjul5uxmn; 
  wire                          yueav99q0b7x3rcm9_x625j6yd; 
  wire                          c7y5emtdpd3rk_dus5ixb7r44; 

  wire                          xnvidl2ouve1vln7ywwu6a5v;
  wire                          k0ue65kc80maq9qkm04zau8h4bz;
  wire                          we3r29j8uhskq7kyw558l15b7  ;
  wire                          vsf0g6h63ew3evcsozmlfhinvhq;
  wire[64-1:0]        yzi326ahunke54273wsh5pgc7kka; 
  
  wire                          qp6hat5pdku7yc9bq1vsm6hb_w9;
  wire                          n0pfd6t_58aep4y4wg7wl9vo7ejyz;
  wire                          f1t_hrt88trjzo1oeoj3ui9lhcu  ;
  wire                          qah4iiv5ntbmab46ir87_rkxcqzih4;
  wire[64-1:0]        nud3tr5ire99qpl6xy6s2vj0; 

  wire                          flb64u531jaudptz5l9y7ju5;
  wire                          so7wnp3pfxe74elogsol7qrvj_5;
  wire  [32-1:0]   z6x6vtfm5ozsb8e1g3ek9mxcaavx; 
  wire                          nsvtf_9m6sep1hb1kltgl2hlnqn; 
  wire  [64-1:0]        odd4wynvno2o6hjyvi65l10zi;
  wire  [8-1:0]     zbpyr_m9c2hqfkc019qkpou4krbxw;
  wire  [2:0]                   l0tlr34v20v3hk8a6gie4uk91yp1w;
  wire  [1:0]                   riimr6qwir1dx_guosj51l91;
  wire                          szfy9s6lzimlb2j3cs5_vlwl;
  wire                          vqq0vkkbq8gqc1tz1k_ud7rm42za;
  wire  [1:0]                   frs0vh2vwgovicyibkf_d3sr6_;
  wire                          x7bhi63pp_k_4diubx18eq_x6c; 
  wire                          vmucahlss7dpuvf0zo7r14es8mw4e; 
  wire                          j46f_ypuqx8_ubhj2dqsl2nvo3xl2; 
  wire                          s5m9cu2ee3zjqralllxvdcnv_nr; 
  wire                          hycfweaqoatse84iuu9rp; 

  wire                          lxdia3j_hv2zwfjcp0_5bnsv3xu;
  wire                          kf17agt2l21y8meszqlaks6n;
  wire  [32-1:0]   w2rebtphwb45_nf6qw5dy26z; 
  wire                          ypdw34_kup0gaiwjzl4bcthak; 
  wire  [64-1:0]      yg5d3o1ke2l9iz9fexcwz4ndh;
  wire  [8-1:0]      t43psmvm15g070eibanybptz7;
  wire  [2:0]                   wz17_6fsan5b1vvg2gbkburw2;
  wire  [1:0]                   wbp0e817xt2uj0bm5047co29g9jr;
  wire                          kzneydeew74np7qbndwhvw_;
  wire                          rywjhkc2m319gtnl68n6yia0h;
  wire  [1:0]                   xqr6qbo6fxrb8hni14at1bkd1o;
  wire                          rr_kd00n0nzd08jhv6de62tu5w2e; 
  wire                          ci_vdf2vqsfb45ipjbbj2kf0g; 
  wire                          cm2iw9jkt_zvly6ri5f7s0sz3q; 
  wire                          r048om6_elh04xzuybqp1x5ynfs4um; 
  wire                          zjg4nl981npxovpev0e_yqz4; 

  wire                          duzcgyd7bbw3jp7bax5m_im68gt;
  wire                          w0414mghkbrhfheu2cmwalfj9g0;
  wire                          ibfxlpjz4f428kdyrvz2l243b__  ;
  wire                          zdq146b5sl9b_zsw84kq0l8u51ph;
  wire[64-1:0]        b49a3gf23ov9g7xpe88_11si96vh; 
  
  wire                          rwfis2p5oqcxun3vrabpu4ehd;
  wire                          ssgsllp8a48t220i6zawign01kjs;
  wire                          pb5hz9n6i21hdl1f9ktx2pf4s  ;
  wire                          gqcennvw7i4s9ra6nufl5auv9n2;
  wire[64-1:0]        zie7s8nvi9nxy9tbeenymedx2ch; 


  wire                          rinamilgle00i5xmx_vt;
  wire                          j8wlfupbw25hdmohz5q0;
  wire  [32-1:0]   z64bwdr23steb7s9y9j; 
  wire                          bg1spy6_v2kbo75pz1d6; 
  wire  [64-1:0]        xyeq7c6icdac80_y0jup;
  wire  [8-1:0]     za5ms2soyuucfxo_jbn;
  wire  [2:0]                   b7aet1zp_fcfxn8h7rw0u1;
  wire  [1:0]                   t3szwnvfo2nj3wk6r5kvt;
  wire                          m4x1_gvw8v_sc8h7c8_6;
  wire                          hpeqnhpztp9l_d3yx16l;
  wire  [1:0]                   bngbyv57e7juc0vkk2y8i;
  wire                          cneu8a119tg3vmie6zr2h_; 
  wire                          jw2dzv9gi7gygudyqql6fz; 
  wire                          o_7kpry6inkqpqi1bf1nd; 
  wire                          f97tgz_qybmvln6nz5dqt458; 
  wire                          znotwr53pu47f5m1agm; 

  wire                          zf_v02okbs8_euhd64;
  wire                          wq4r8m45isqp8_o4pdtitz;
  wire  [32-1:0]   qpzo6lin6brrytho7; 
  wire                          k7j6g0757jovg8xstgrvwf; 
  wire  [64-1:0]      nwx86gohbrn08nvh60789;
  wire  [8-1:0]      bebhplbk2k43sfoehvt66w;
  wire  [2:0]                   ljk3q52m5tirt6shbcwbf;
  wire  [1:0]                   ucj9poqgl683ej1pihkh;
  wire                          u9hi0xtx8u0mn0l_7p;
  wire                          rm04yhu6ondli9u0g6din;
  wire  [1:0]                   o5fmtstd7kef7z4m7jefm;
  wire                          vvadj6ew1h5wq9z5askkzr9; 
  wire                          lop06h0_z_4tt1s04up; 
  wire                          ivllgcn1kiix2iamzwf0u; 
  wire                          rnmvpk356vfgxd_045g; 
  wire                          a46c4xo4texvc9o; 

  wire                          ze2bfnigu62i9937pcxnjc;
  wire                          c86b14qr2qo45_qw2ns;
  
  wire                          mm70cenjp_1wmcs135nh4wl;
  wire                          p4dpiqc4w_g42ni5jsaj;


  wire [uw3hbdikblihw1_r3o-1:0] hgzu6a1jtp0nlbtwfmavcuox3sbr;
  wire [uw3hbdikblihw1_r3o-1:0] mu65khgqx0z95knlzx6iei9q0;
  wire [uw3hbdikblihw1_r3o-1:0] xvd66h85myby1si3gcpihi2q;
  wire [uw3hbdikblihw1_r3o-1:0] ahdyrung86cgxxtsd2oudlh;
  wire [uw3hbdikblihw1_r3o-1:0] yhwduf8bvuhcs65ehz;
  wire [uw3hbdikblihw1_r3o-1:0] w7k_388auwycpor_bf4;

  wire [uw3hbdikblihw1_r3o-1:0] of253wss1uu2rupz6abzptzor3a;
  wire [uw3hbdikblihw1_r3o-1:0] cioxj8lmdlu0ysr1dt0ogp6gjf;

  assign 
       hgzu6a1jtp0nlbtwfmavcuox3sbr = { 
       q064m0tgrtkrz7vn_qf2bjb, 
       xxrb4v2suklf9djaeyf0rkmedjz3, 
       hrn1giqg1k6gbt6q7lrxzxaqztx,
       xw04i4vzqgn2m2ihbdv55m4bvtr,
       h_9b0wqhlkmvxkfizht97cqp,
       ycmo1kcbjq1scw4gwg4uiwd_,
       ocdu63ksnvvgacaermakucm0f4g,
       oxlxxz2rxp0amufq1s9jqrry3y,
       rcpyv929ixr6xhyeyg2p0cgtj,
       n169ohp8pq9l7goaugowzjfa, 
       psec5ihpqk4slg2u90eq4yzyy, 
       cv6960ns7f2dyrvj6ij_phb0, 
       kxqipwn8s_54dje1dpjvcgaye6t, 
       gc_aq81uy3hbdq8ns7y1_ckg};

  assign 
       mu65khgqx0z95knlzx6iei9q0 = { 
       kbbc76s46hvu_3te0ihj3hb2nl, 
       g33u_ys44gmrebks2nd9y8o, 
       y5gfh4gmog9i5iq47qq3nmc95_fnd,
       bafx6nbdipfv60zavyhkpt5ulfqp,
       wfq3yog1gp3v5k8ew8aazeio5q9qm,
       bkec53bqczw0o6vx2ouxlbp,
       o347ncxtm6aeg09kb47k1oggzcw,
       pfkm_ekt4p23xk05wj0f5ei8wut2,
       rx7d01wkjl49umakx8rnira0bvj,
       bpetbkuwyy1k6fa142bfw3rz7sjpi, 
       vsn6zt6npfa5qvbab0qrm7ya, 
       c_saxxol2d2vxelssdxtjul5uxmn, 
       yueav99q0b7x3rcm9_x625j6yd, 
       c7y5emtdpd3rk_dus5ixb7r44};

  assign 
       xvd66h85myby1si3gcpihi2q = { 
       z6x6vtfm5ozsb8e1g3ek9mxcaavx, 
       nsvtf_9m6sep1hb1kltgl2hlnqn, 
       odd4wynvno2o6hjyvi65l10zi,
       zbpyr_m9c2hqfkc019qkpou4krbxw,
       l0tlr34v20v3hk8a6gie4uk91yp1w,
       riimr6qwir1dx_guosj51l91,
       szfy9s6lzimlb2j3cs5_vlwl,
       vqq0vkkbq8gqc1tz1k_ud7rm42za,
       frs0vh2vwgovicyibkf_d3sr6_,
       x7bhi63pp_k_4diubx18eq_x6c, 
       vmucahlss7dpuvf0zo7r14es8mw4e, 
       j46f_ypuqx8_ubhj2dqsl2nvo3xl2, 
       s5m9cu2ee3zjqralllxvdcnv_nr, 
       hycfweaqoatse84iuu9rp};

  assign  
       ahdyrung86cgxxtsd2oudlh = { 
       w2rebtphwb45_nf6qw5dy26z, 
       ypdw34_kup0gaiwjzl4bcthak, 
       yg5d3o1ke2l9iz9fexcwz4ndh,
       t43psmvm15g070eibanybptz7,
       wz17_6fsan5b1vvg2gbkburw2,
       wbp0e817xt2uj0bm5047co29g9jr,
       kzneydeew74np7qbndwhvw_,
       rywjhkc2m319gtnl68n6yia0h,
       xqr6qbo6fxrb8hni14at1bkd1o,
       rr_kd00n0nzd08jhv6de62tu5w2e, 
       ci_vdf2vqsfb45ipjbbj2kf0g, 
       cm2iw9jkt_zvly6ri5f7s0sz3q, 
       r048om6_elh04xzuybqp1x5ynfs4um, 
       zjg4nl981npxovpev0e_yqz4};

  assign 
       { 
       z64bwdr23steb7s9y9j, 
       bg1spy6_v2kbo75pz1d6, 
       xyeq7c6icdac80_y0jup,
       za5ms2soyuucfxo_jbn,
       b7aet1zp_fcfxn8h7rw0u1,
       t3szwnvfo2nj3wk6r5kvt,
       m4x1_gvw8v_sc8h7c8_6,
       hpeqnhpztp9l_d3yx16l,
       bngbyv57e7juc0vkk2y8i,
       cneu8a119tg3vmie6zr2h_, 
       jw2dzv9gi7gygudyqql6fz, 
       o_7kpry6inkqpqi1bf1nd, 
       f97tgz_qybmvln6nz5dqt458, 
       znotwr53pu47f5m1agm} =
       yhwduf8bvuhcs65ehz;

  assign  
       {
       qpzo6lin6brrytho7, 
       k7j6g0757jovg8xstgrvwf, 
       nwx86gohbrn08nvh60789,
       bebhplbk2k43sfoehvt66w,
       ljk3q52m5tirt6shbcwbf,
       ucj9poqgl683ej1pihkh,
       u9hi0xtx8u0mn0l_7p,
       rm04yhu6ondli9u0g6din,
       o5fmtstd7kef7z4m7jefm,
       vvadj6ew1h5wq9z5askkzr9, 
       lop06h0_z_4tt1s04up, 
       ivllgcn1kiix2iamzwf0u, 
       rnmvpk356vfgxd_045g, 
       a46c4xo4texvc9o} = 
       w7k_388auwycpor_bf4;

  assign 
       { 
       a45qubts5uovcopirpl9jxs7uia, 
       kwbu6olmnnt53fot6kfntm2q7t, 
       kq9lkjt85jst7fa5smg1nud,
       mekhipn8vmxn5adno3jrpek8nkm,
       wbwviedmyjzfiwi2t1yh0ibf7wv3,
       h99v8xeu9gkycpsn1wl3lrow7,
       jvloelo3plm6zwbisesi7fwa,
       ecz8u30wtuyonhyfwfrfrc30g,
       vxwea8jbxv6m5tu7nkqtf6,
       jsswxoezxjsdw154f5xt1omqrup, 
       e5cyxxxkg4061gq3_ksqdax_7op, 
       m3pduyvpfh4ximuy0dl6k_wjuc, 
       xhts19tgn12c186fduss6cfjyz, 
       zt7xddfgq3m2nsc8s_3a48r8} =
       of253wss1uu2rupz6abzptzor3a;

  assign 
       { 
       gi8g2jgc5r69ozgg2517f4, 
       nqq4y60r7eh5lbir_nzlqf2q7k, 
       rf_rtoowzj9m6zi6taqyqn6ku,
       kqa4ro7t84z342uqr2plzmi1,
       d50l6nnxdfj7iuhnqe9gjobewaj4,
       ziqf65e93q9kc_6bj_n4gd2op,
       lkflakila483fdjdz1hrtobjiz,
       zg0qkr8fhe1v0eku3at17q,
       gu2ufdscjjb3hvpwrwu6c8h,
       pn9rf9nl21n4t8clpsygzbo72n, 
       u6t2h_hm580phvwuvdedyagaqg, 
       h1p8zhyrvirdo9c78wx8cmal83, 
       d11v3v5k967aul6l7_up53azs, 
       tnfd_mhtdr0hw58lveup8w8} =
       cioxj8lmdlu0ysr1dt0ogp6gjf;

  wire [szbi56su117rxsuhhun-1:0] v4756d8xk0jqi9j0qedfnm2;
  wire [szbi56su117rxsuhhun-1:0] v7pt_kohuazs2hduan3ewo5r7j;
  wire [szbi56su117rxsuhhun-1:0] xmygo7hdickwkqu1107gh0ofld;
  wire [szbi56su117rxsuhhun-1:0] c9hib9fb61pjgp772_89fllik;
  wire [szbi56su117rxsuhhun-1:0] mavn74e1rxaempydhr;
  wire [szbi56su117rxsuhhun-1:0] yda8t9dlz43knw4vi;

  wire [szbi56su117rxsuhhun-1:0] ot_thh6tdm6pci9nju5b6t;
  wire [szbi56su117rxsuhhun-1:0] o0oddj2hd8ur16vx2shbs8_;

  assign {
                                    we3r29j8uhskq7kyw558l15b7  ,
                                    vsf0g6h63ew3evcsozmlfhinvhq,
                                    yzi326ahunke54273wsh5pgc7kka} = v4756d8xk0jqi9j0qedfnm2; 

  assign {
                                    ibfxlpjz4f428kdyrvz2l243b__  ,
                                    zdq146b5sl9b_zsw84kq0l8u51ph,
                                    b49a3gf23ov9g7xpe88_11si96vh} = v7pt_kohuazs2hduan3ewo5r7j; 


  assign {
                                    f1t_hrt88trjzo1oeoj3ui9lhcu  ,
                                    qah4iiv5ntbmab46ir87_rkxcqzih4,
                                    nud3tr5ire99qpl6xy6s2vj0} = xmygo7hdickwkqu1107gh0ofld; 

  assign {
                                    pb5hz9n6i21hdl1f9ktx2pf4s  ,
                                    gqcennvw7i4s9ra6nufl5auv9n2,
                                    zie7s8nvi9nxy9tbeenymedx2ch} = c9hib9fb61pjgp772_89fllik; 


  assign ot_thh6tdm6pci9nju5b6t = {
                                    gz2qngl9towiwc_nk48gu38p9  ,
                                    saolr4xnpfm570snrsqk7hazshkz,
                                    b85cqul2sjbg0c5ta0bcpgpluvma};

  assign o0oddj2hd8ur16vx2shbs8_ = {
                                    byn2o0bi_9ggzegrnvskn  ,
                                    m12x1nn4kvsdeqofo9rqi8aawa,
                                    e0xiuuzhk1qbwdjlub9o_cca5};

  wire no360dfthc_r812ltoqdhrz;
  wire piosx1_uvpor01vn8ll66_yhit;
  wire j9o_ty1uw4uvham3ak;
  
  
  
  wire  xzz_39w6q2zpq6egp9ojdui_ = 
        (bidjco9v6uwp91tvsqnp72df_u0q & (~flb64u531jaudptz5l9y7ju5)) 
      | (bidjco9v6uwp91tvsqnp72df_u0q & flb64u531jaudptz5l9y7ju5 & (j9o_ty1uw4uvham3ak == 1'b0));

  wire  s8ld7ymugb8dqx60x5okhsd3 = 
        (flb64u531jaudptz5l9y7ju5 & (~bidjco9v6uwp91tvsqnp72df_u0q)) 
      | (flb64u531jaudptz5l9y7ju5 & bidjco9v6uwp91tvsqnp72df_u0q & (j9o_ty1uw4uvham3ak == 1'b1));

  wire  ef5131xxhh6i_flah2f1mpt = 
        (vkjwr2hxue8911qmv5ro35cg & (~lxdia3j_hv2zwfjcp0_5bnsv3xu)) 
      | (vkjwr2hxue8911qmv5ro35cg & lxdia3j_hv2zwfjcp0_5bnsv3xu & (j9o_ty1uw4uvham3ak == 1'b0));

  wire  dvtbmm8px0fy141v1gn67d = 
        (lxdia3j_hv2zwfjcp0_5bnsv3xu & (~vkjwr2hxue8911qmv5ro35cg)) 
      | (lxdia3j_hv2zwfjcp0_5bnsv3xu & vkjwr2hxue8911qmv5ro35cg & (j9o_ty1uw4uvham3ak == 1'b1));

  wire  opa_i9g_7se8iof9su_mxicjyu = 
        (no360dfthc_r812ltoqdhrz & (~piosx1_uvpor01vn8ll66_yhit)) 
      | (no360dfthc_r812ltoqdhrz & piosx1_uvpor01vn8ll66_yhit & (j9o_ty1uw4uvham3ak == 1'b0));

  wire  n1bimos0aw0citrgtz3yco = 
        (piosx1_uvpor01vn8ll66_yhit & (~no360dfthc_r812ltoqdhrz)) 
      | (piosx1_uvpor01vn8ll66_yhit & no360dfthc_r812ltoqdhrz & (j9o_ty1uw4uvham3ak == 1'b1));


  wire rj0pmrnp69j8jdw7m77j;

  f2w7478x4kvdp7gsxub2tls31 #(
    .f16zrowg1s1f5   (uw3hbdikblihw1_r3o),
    .mp26klefy4v2f   (szbi56su117rxsuhhun),
    .cu7ihzi5k8   (nsy582liduihtlix7j5),
    .cqf2oxizzealhe   (1) 
  ) bvan0yb0t_khtcy6f2vix4fp(
  
    .ffckqqivts0p     (xzz_39w6q2zpq6egp9ojdui_),
    .yseo05ez9cr0r     (s8ld7ymugb8dqx60x5okhsd3),
    .g5ptjmebcoo5nwcg (bidjco9v6uwp91tvsqnp72df_u0q),
    .pjmu7ih6ul43bacz (m83gf40i8n5qmmo860pq3w7n5n5f),
    .s6tktwbreyy7r  (hgzu6a1jtp0nlbtwfmavcuox3sbr ),
    .h014w4n6dlj78fr3 (ycmo1kcbjq1scw4gwg4uiwd_[0]),
    .jf6zw884wuj   (ycmo1kcbjq1scw4gwg4uiwd_[1]),
  
    .l1mjv4a3o1i7qxeru (xnvidl2ouve1vln7ywwu6a5v),
    .vmc_730ubm6z6mit (k0ue65kc80maq9qkm04zau8h4bz),
    .ok1b1b_3nv0  (v4756d8xk0jqi9j0qedfnm2 ),
  
    .sgk1y63o9l50k3 (flb64u531jaudptz5l9y7ju5),
    .gqhewm9l9lvfgkbf7 (so7wnp3pfxe74elogsol7qrvj_5),
    .mchi632scfby1t0n  (xvd66h85myby1si3gcpihi2q ),
    .ofjszjvfai0r49q (riimr6qwir1dx_guosj51l91[0]),
    .mlewhkn_ph   (riimr6qwir1dx_guosj51l91[1]),
  
    .eapg2epq1a388t4 (duzcgyd7bbw3jp7bax5m_im68gt),
    .osuxnyc17r3xf (w0414mghkbrhfheu2cmwalfj9g0),
    .sy8hpqbz5umprdog  (v7pt_kohuazs2hduan3ewo5r7j ),
  
    .nk9dw9ied4zd2h  (rinamilgle00i5xmx_vt),
    .czec2uuagggq  (j8wlfupbw25hdmohz5q0),
    .d5xonxqryf7   (yhwduf8bvuhcs65ehz),
  
    .qegs8svpsb6wzol  (ze2bfnigu62i9937pcxnjc),
    .k0csx0ynvoz54fjx  (c86b14qr2qo45_qw2ns),
    .c20li_6i3x   (mavn74e1rxaempydhr),
  
    .f5lbzfpsc02anbqy (rj0pmrnp69j8jdw7m77j),

    .gf33atgy         (gf33atgy),
    .ru_wi       (ru_wi)
  );

  wire d4ky0qxli8vpovkpsv1;

  f2w7478x4kvdp7gsxub2tls31 #(
    .f16zrowg1s1f5   (uw3hbdikblihw1_r3o),
    .mp26klefy4v2f   (szbi56su117rxsuhhun),
    .cu7ihzi5k8   (nsy582liduihtlix7j5),
    .cqf2oxizzealhe   (1) 
  ) bx03gkfg2cg7g92__pvji45cje(

    .ffckqqivts0p     (ef5131xxhh6i_flah2f1mpt),
    .yseo05ez9cr0r     (dvtbmm8px0fy141v1gn67d),
  
    .g5ptjmebcoo5nwcg (vkjwr2hxue8911qmv5ro35cg),
    .pjmu7ih6ul43bacz (xronfobw50555i02avvye82b),
    .s6tktwbreyy7r  (mu65khgqx0z95knlzx6iei9q0 ),
    .h014w4n6dlj78fr3 (bkec53bqczw0o6vx2ouxlbp[0]),
    .jf6zw884wuj   (bkec53bqczw0o6vx2ouxlbp[1]),
  
    .l1mjv4a3o1i7qxeru (qp6hat5pdku7yc9bq1vsm6hb_w9),
    .vmc_730ubm6z6mit (n0pfd6t_58aep4y4wg7wl9vo7ejyz),
    .ok1b1b_3nv0  (xmygo7hdickwkqu1107gh0ofld ),
  
    .sgk1y63o9l50k3 (lxdia3j_hv2zwfjcp0_5bnsv3xu),
    .gqhewm9l9lvfgkbf7 (kf17agt2l21y8meszqlaks6n),
    .mchi632scfby1t0n  (ahdyrung86cgxxtsd2oudlh ),
    .ofjszjvfai0r49q (wbp0e817xt2uj0bm5047co29g9jr[0]),
    .mlewhkn_ph   (wbp0e817xt2uj0bm5047co29g9jr[1]),
  
    .eapg2epq1a388t4 (rwfis2p5oqcxun3vrabpu4ehd),
    .osuxnyc17r3xf (ssgsllp8a48t220i6zawign01kjs),
    .sy8hpqbz5umprdog  (c9hib9fb61pjgp772_89fllik ),
  
    .nk9dw9ied4zd2h  (zf_v02okbs8_euhd64),
    .czec2uuagggq  (wq4r8m45isqp8_o4pdtitz),
    .d5xonxqryf7   (w7k_388auwycpor_bf4),
  
    .qegs8svpsb6wzol  (mm70cenjp_1wmcs135nh4wl),
    .k0csx0ynvoz54fjx  (p4dpiqc4w_g42ni5jsaj),
    .c20li_6i3x   (yda8t9dlz43knw4vi),

    .f5lbzfpsc02anbqy (d4ky0qxli8vpovkpsv1 ),
  
    .gf33atgy         (gf33atgy),
    .ru_wi       (ru_wi)
  );

  wire vi4wgos18sjty012c =  rinamilgle00i5xmx_vt;
  wire i3d14osds0zjqeii = ~rinamilgle00i5xmx_vt;


  f2w7478x4kvdp7gsxub2tls31 #(
    .f16zrowg1s1f5   (uw3hbdikblihw1_r3o),
    .mp26klefy4v2f   (szbi56su117rxsuhhun),
    .cu7ihzi5k8   (nsy582liduihtlix7j5),
    .cqf2oxizzealhe   (1) 
  ) vfp2x5uo14ndbi3ii8i3giuu(

    .ffckqqivts0p     (vi4wgos18sjty012c),
    .yseo05ez9cr0r     (i3d14osds0zjqeii),
  
    .g5ptjmebcoo5nwcg (rinamilgle00i5xmx_vt),
    .pjmu7ih6ul43bacz (j8wlfupbw25hdmohz5q0),
    .s6tktwbreyy7r  (yhwduf8bvuhcs65ehz ),
    .h014w4n6dlj78fr3 (t3szwnvfo2nj3wk6r5kvt[0]),
    .jf6zw884wuj   (t3szwnvfo2nj3wk6r5kvt[1]),
  
    .l1mjv4a3o1i7qxeru (ze2bfnigu62i9937pcxnjc),
    .vmc_730ubm6z6mit (c86b14qr2qo45_qw2ns),
    .ok1b1b_3nv0  (mavn74e1rxaempydhr ),
  
    .sgk1y63o9l50k3 (zfu2vonacwweg65jwl5h),
    .gqhewm9l9lvfgkbf7 (ecc0pa6dsujd5fk_ztk1odty),
    .mchi632scfby1t0n  (a23lzk9_jpf1wt6gpoa3t ),
    .ofjszjvfai0r49q (vo4iscd43mm129ts9g7[0]),
    .mlewhkn_ph   (vo4iscd43mm129ts9g7[1]),
  
    .eapg2epq1a388t4 (z9q40jbnm38zcodsjsd090z),
    .osuxnyc17r3xf (i0znoodcvzhh4rexar7joqvk),
    .sy8hpqbz5umprdog  (kti_aenofx1syww4og3 ),
  
    .nk9dw9ied4zd2h  (rjy1ysvx9590bpklijsn0ucgaga),
    .czec2uuagggq  (d_933icutbtk8nknxip5t1ds),
    .d5xonxqryf7   (of253wss1uu2rupz6abzptzor3a),
  
    .qegs8svpsb6wzol  (fp_qm6eq7380_uydc6pb2sw7),
    .k0csx0ynvoz54fjx  (z9eviza6dmjc6u7jbuzirzh8z1ce),
    .c20li_6i3x   (ot_thh6tdm6pci9nju5b6t),
  
    .f5lbzfpsc02anbqy (),

    .gf33atgy         (gf33atgy),
    .ru_wi       (ru_wi)
  );

  wire amyj2vwd59trjfwu3  =  zf_v02okbs8_euhd64;
  wire vm5sjyldzo48q7w = ~zf_v02okbs8_euhd64;


  f2w7478x4kvdp7gsxub2tls31 #(
    .f16zrowg1s1f5   (uw3hbdikblihw1_r3o),
    .mp26klefy4v2f   (szbi56su117rxsuhhun),
    .cu7ihzi5k8   (nsy582liduihtlix7j5),
    .cqf2oxizzealhe   (1) 
  ) x9yzda0b_kj2ulywb3g9jf(
    .ffckqqivts0p     (amyj2vwd59trjfwu3),
    .yseo05ez9cr0r     (vm5sjyldzo48q7w),
  
    .g5ptjmebcoo5nwcg (zf_v02okbs8_euhd64),
    .pjmu7ih6ul43bacz (wq4r8m45isqp8_o4pdtitz),
    .s6tktwbreyy7r  (w7k_388auwycpor_bf4 ),
    .h014w4n6dlj78fr3 (ucj9poqgl683ej1pihkh[0]),
    .jf6zw884wuj   (ucj9poqgl683ej1pihkh[1]),
  
    .l1mjv4a3o1i7qxeru (mm70cenjp_1wmcs135nh4wl),
    .vmc_730ubm6z6mit (p4dpiqc4w_g42ni5jsaj),
    .ok1b1b_3nv0  (yda8t9dlz43knw4vi ),
  
    .sgk1y63o9l50k3 (ejbq7zgkpgwgttfvvx5rp),
    .gqhewm9l9lvfgkbf7 (agtve46c928tzy8367oy14bf),
    .mchi632scfby1t0n  (nzcpulhcv_r50wph3pz9 ),
    .ofjszjvfai0r49q (edt_9_yofk03w8y7jt[0]),
    .mlewhkn_ph   (edt_9_yofk03w8y7jt[1]),
  
    .eapg2epq1a388t4 (gcan4qd32d7splx9secvc8b),
    .osuxnyc17r3xf (q2_zn_ozuoxddlj2se_t45w),
    .sy8hpqbz5umprdog  (cmvo1gt96vee3wmg9e ),
  
    .nk9dw9ied4zd2h  (pkm6vgcr8iz_el5103gzwdew0hki),
    .czec2uuagggq  (vdbkch1krpijvuukam8k5_9g6h4d),
    .d5xonxqryf7   (cioxj8lmdlu0ysr1dt0ogp6gjf),
  
    .qegs8svpsb6wzol  (me8sa0hl_2m6xmtdm4r_1tn7cer4),
    .k0csx0ynvoz54fjx  (gv_wy8qy9rm50mn4yg66yvagb60l),
    .c20li_6i3x   (o0oddj2hd8ur16vx2shbs8_),
  
    .f5lbzfpsc02anbqy (),

    .gf33atgy         (gf33atgy),
    .ru_wi       (ru_wi)
  );

  wire                       khbwxlyuzlnl1c8t8_3og_5mq; 
  wire [64-1:0] qnthfit20wgbpxec8thtex71gzm7;  
  wire                       ddrezcee7228fcb3xe5ptlosy;  

  wire                       kn4nyomkyc9nib4jk3q9v9u; 
  wire [64-1:0] ms19_yn0emkdebo5xds5no7own3k;  
  wire                       koyy03uze4eek43dncxyfucn2;  
  
  wire                       hystveyc5mdp2fsv1prg; 
  wire [64-1:0] cqnseh0h9l57x_6_lagpk2_zv;  
  wire                       zi8qhl5upl3l4fr_x69d9;  

  wire                       xirk22lqyoyt4_ojp1k3vkzye; 
  wire [64-1:0] bo3wo9aretoipldnjadceyp2kgl;  
  wire                       li46sayiwuz6fbzu8n2xux;  
  
  wire                       tzuvc0ejdqdp8s;
  wire [64-1:0] yf9xpz2g2m0w8qlt13b21y2;  
  wire                       loifq6epc1ba16z5f;  

  wire                       ozyjhnq394jxng;
  wire [64-1:0] b0r1ara7cbtyek7a_1z;  
  wire                       n0qoqq4p_4wb45uxep7;  


  assign tzuvc0ejdqdp8s      = d4ky0qxli8vpovkpsv1 ? kn4nyomkyc9nib4jk3q9v9u      :  khbwxlyuzlnl1c8t8_3og_5mq     ;
  assign yf9xpz2g2m0w8qlt13b21y2 = d4ky0qxli8vpovkpsv1 ? ms19_yn0emkdebo5xds5no7own3k :  qnthfit20wgbpxec8thtex71gzm7;
  assign loifq6epc1ba16z5f     = d4ky0qxli8vpovkpsv1 ? koyy03uze4eek43dncxyfucn2     :  ddrezcee7228fcb3xe5ptlosy    ;
  
  assign ozyjhnq394jxng      = rj0pmrnp69j8jdw7m77j ? xirk22lqyoyt4_ojp1k3vkzye      :  hystveyc5mdp2fsv1prg     ;
  assign b0r1ara7cbtyek7a_1z = rj0pmrnp69j8jdw7m77j ? bo3wo9aretoipldnjadceyp2kgl :  cqnseh0h9l57x_6_lagpk2_zv;
  assign n0qoqq4p_4wb45uxep7     = rj0pmrnp69j8jdw7m77j ? li46sayiwuz6fbzu8n2xux     :  zi8qhl5upl3l4fr_x69d9    ;
  
  wire                          lr0ugrb30q4zc;
  wire [64-1:0]    uq8tdw3q3f22qrubbs;  
  wire                          n7_nwy7dhha;  

  assign lr0ugrb30q4zc      = ozyjhnq394jxng ? ozyjhnq394jxng      :  tzuvc0ejdqdp8s     ;
  assign uq8tdw3q3f22qrubbs = ozyjhnq394jxng ? b0r1ara7cbtyek7a_1z :  yf9xpz2g2m0w8qlt13b21y2;
  assign n7_nwy7dhha     = ozyjhnq394jxng ? n0qoqq4p_4wb45uxep7     :  loifq6epc1ba16z5f    ;
  
  ux607_gnrl_dffr #(1)                bvdctt0qoczifysk       (            lr0ugrb30q4zc,      tjzl_75hfxv6m,      gf33atgy, ru_wi);

  ux607_gnrl_dfflr #(64) ypcw7brxx3f57v4hkekd_62 (lr0ugrb30q4zc, uq8tdw3q3f22qrubbs, ay20xnz1tx3gv1k, gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1)               yuqi8sfyk58ynnr     (lr0ugrb30q4zc, n7_nwy7dhha    , fyo0ut7e82c,     gf33atgy, ru_wi);


  wire                        ye2fnsl_jl2n9kk6; 
  wire                        ctqj_dyrttnfzu9lcud3g_3; 

  wire                        i2hiwgez7xp0bc_3mg35a4rb;
  wire                        lwl5fn5x_gxnq3f3a1tt0qyrd;

  wire [32-1:0]  gwy4w6j_23g_d3t; 
  wire                        xknh2ut7lctvrugsz5wb; 
  wire                        g3itms8el25jimpco2t_yu4; 
  wire [64-1:0]       w_fuqyygyv_7yus0ow9k;
  wire [8-1:0]    ld964zre2gsugp9blpo;
  wire                        h5986karddzxifsa9t; 
  wire                        ya7g9x7j5jke20pxxk; 
  wire                        hyiwh018ufcuat94ohr4; 
  wire                        mdw031z1stmwv1atvh9pla6; 
  wire                        kqe4mxh6t85yt1es15h_kv3y_; 
  wire                        eidxuo2trad883370opeq; 
  wire                        yz4xms1_6ldn__afmhfdxic; 
  wire                        k6aoxxoxugbmismespiv2pfhf; 
  wire                        g6zc5qflpket_8b_30jviei4n; 
  wire                        ff8kz54m27i8p1qxp4c_n1y; 
  wire                        lm8vcj797bp12bltgigc6lk76ei1; 
  wire                        cnh34kai5koa_4iw5boo0p; 

  wire                        lszyvs15rstcbyhj96v090d;
  wire                        iqj11baw8n07djxz1m45yxd  ;
  wire                        wx_fs2ijrykfgpoqldrgukw  ;
  wire[64-1:0]        tfwuip_0npwfy19ek9gpoc; 
 



  wire                          on12sjnlw0b975rtxnj;
  wire                          m91uirvkay9adfjui930dyv4;
  wire                          a_i3c4odzkmjpufk2pffcu;

  wire                          i691bnr_y8gmwnd0nsaw;
  wire                          isqt1ng7lccfet8bj5hym5c;
  wire [24-1:0]  ije4h78_umvknjj6az4_5qf92e3iydh;
  wire [24-1:0]  sro97_d1rgt1fmqi2b_fitscvexczye2;
  wire [32-1:0]  v2tse065uysfbl8f4z8hlpkg5o68;
  wire [32-1:0]  kwczwxezdeidftn2_p2fpzik3gt;
  wire [32-1:0]  o58xzacx8hg_9zcqk21v9m0rqqsap22_;
  wire [32-1:0]  q0xni3yf49f2fj7ymo_nvdurqx1okyv;

  wire                          rbkhb89tyu_ucjpo;  
  wire [6-1:0]  sqvgnqdrkexeg2lziofadt;
  wire                          bwtzw5pqhc62g9v9w ;
  wire [24-1:0]  nwbvll63g8yq6vbpxok;          
  
  wire                          e4ui35hoxqcwkgfaol;  
  wire [6-1:0]  f1uy000fu6355gukzxt9r4y; 
  wire                          avudrqvyzx1dringrt4rs ;
  wire [24-1:0]  hz5leo9sklh2v25_50;          


  wire                          ofg0te04_oeiba586;  
  wire [8-1:0] dm0uaanzcp_7hojw2_h; 
  wire [4-1:0] yddyulfbyf7p2wvl6dyk;
  wire [32-1:0] j233e_ya9xhnxg7flb9d3;          
  
  wire                          mq3a_g7zrfyfdil1;  
  wire [8-1:0] f9ekxi98w3bnnfm3t1vyt1; 
  wire [4-1:0] k1vhaduoq3xy5cx6jr0;
  wire [32-1:0] hwo9njh5b4299teslcl;          
 
  wire                          shxdziymfk57c49e0;  
  wire [8-1:0] s_fatq1jfpqkf7q9d40n; 
  wire [4-1:0] ruix76vs69a8gynr7yydnp;
  wire [32-1:0] y0s6zoimyz170437bgkne;          

  wire                          nsyif4pw3tzuggdakg2;  
  wire [8-1:0] e4zsuzpz_sgcgql5k19iv; 
  wire [4-1:0] fvzgpoei5_ffhtrv6r;
  wire [32-1:0] cnqt629_5e9xaypczfdt;         

  wire                        mvkoyonaqzuf3ip; 
  wire                        eca4wu5z1eltuvtu76r7ti6; 

  wire                        aq3hy9uuv5rnvzphrnaa3;
  wire                        rho1guu79090z97aekm9s16pn;

  wire [32-1:0]  xnmq3kuajinzxdfiu6q; 
  wire                        xdheobtph1wq8f9ui3h; 
  wire                        nni92t4rn44yvbfgt5yor94mh; 
  wire [64-1:0]       rft88ds492cdh634i;
  wire [8-1:0]    u87rvzwj0xs9vt8uwuot;
  wire                        wawfribsksiyhybl3m1fc; 
  wire                        zfmqdobuh7r4t0fza5uv; 
  wire                        jhiyy3sgiaizu4l4milff; 
  wire                        snm9n0s_9re1n13_p9tec; 
  wire                        ccf5m6bnqnibseotadeyu86cd0; 
  wire                        irncno4zcb4x06mlfiba16bh; 
  wire                        yc59czg2u_bbaxbn1ejpjm8w; 
  wire                        n3r6ftigei07xsagxiifpct; 
  wire                        j8lpsrktt_qs_wo43c_rre4; 
  wire                        ryz4vgf7dpx5dcq733ch1f5gm; 
  wire                        ulggxuvjbou5t00s_czahip80ud3; 
  wire                        kbt5xarx9to2rj956ik1zwwq; 

  wire                        qpzxk_hrtmppd7i7eplel;
  wire                        z85m6lb5ii_p8z196b1r  ;
  wire                        zg97ncjhsfhaqpc60t6wfdr  ;
  wire[64-1:0]        h987z8usv7pyyl5zqvzw4; 
 


  wire [2-1:0] merfg1jkbwck;
  wire [2-1:0] x974z3fncltxj;
  wire [2-1:0] hh2n5p_74cpa;
  wire [2-1:0] yo_tvqeum32rvou;
  wire [2-1:0] trycoh_sgdgtcdg;

  wire [2-1:0] iv9dhbb1gs4h19y;
  wire [2-1:0] k8b8v2d_8bexygcseus;
  wire [2-1:0] cj_amdiu4_4kyqh;
  wire [2-1:0] bcohnzslp6bf6pqn1;
  wire [2-1:0] xlnalzy_jsdbs;

  wire m2s492eolz_a4lrc;

  wire [3-1:0] nyrioysq5ovac5r8 [2-1:0] ;
  

  wire                          a5s2gi2_h7rplzkx1;
  wire                          gn916lc8_fzkp3rcqpob;
  wire                          nepu6mf61h2b2uewptpauek6v;

  wire                          xu6a8p2dk2fy9r7lnn_kd1l;
  wire                          pn1rzse3t9e6g_et37gv;
  wire [24-1:0]  lwmr8fyosc4w78ftaznb17d0wep6;
  wire [24-1:0]  g_lbo1t8r4bx4olr034dfi8fhfw1m6i;
  wire [32-1:0]  xmf6kblqlhyjpa44uj3tn_7hs9g;
  wire [32-1:0]  td_dxcgpaod7g2fvddly_mg4rjh2vgbk;
  wire [32-1:0]  l1mayxu6go0ni6a1uu2tn40qyps5l_;
  wire [32-1:0]  qdf9k5s3p4c0d8jxgmxlyi478ade;

  wire                          idcribpugamfq_39t;  
  wire [6-1:0]  nfuf_njr73sjp5jr12d7gc;
  wire                          hgm8yvqudk9e2ne6 ;
  wire [24-1:0]  ivt9rgs2qqjzyrq5zt4isy;          
  
  wire                          u6di3j5ypwgwjvnmcbsqh;  
  wire [6-1:0]  i7vlo92n37lvcod6oj; 
  wire                          ulp1cmdd07o0vc3p_65wi ;
  wire [24-1:0]  f9_zg3c33q9sbq6d82u;          


  wire                          mgc5k45s6iun0h64mg94n;  
  wire [8-1:0] kuhd9_39ag_1mza9vf7x; 
  wire [4-1:0] dbp3mo7p_zh0242q9;
  wire [32-1:0] enbd230u3ab6jrd2gt;          
  
  wire                          nwvjy589molbkspazci;  
  wire [8-1:0] hkv3jt_7_o_8sk0aait_0kp; 
  wire [4-1:0] dzca_d1t69gei8viv2q;
  wire [32-1:0] w7paq1qa9rrtadyr3v3cx;          
 
  wire                          ky3t5ldjtr_g__hnxr58s;  
  wire [8-1:0] l20gjym8j9s2t31_nhs8iuh; 
  wire [4-1:0] r3kh4eweep0kg7fak6rx6f;
  wire [32-1:0] vwj6zdjeua22z66vj;          

  wire                          tbykhfjbcc3ure59;  
  wire [8-1:0] v0oz07osad44us4h0pyd; 
  wire [4-1:0] xtiqejiid_qbh90nn_jv;
  wire [32-1:0] dzoe86_fm7z7_c7_4_zn;       


  
  wire o0nkaxltg92zc7_vvacwa = p11an_iatsqmyhotqeai;


  wire hy9lwz17ce;
  wire vvzs4gmapk7c ;

  
  wire m4kup76s12og17 = xlnalzy_jsdbs[j9o_ty1uw4uvham3ak];
  wire uy_5bn9r03ydi88m7 = 1'b1;
  wire aliwneheqa6be8dgn = m4kup76s12og17 & uy_5bn9r03ydi88m7;
  wire oyc0vwbyun6num5qh = aliwneheqa6be8dgn;



  wire d1rivbcy3w5oji6yoo = m91uirvkay9adfjui930dyv4 | on12sjnlw0b975rtxnj;
  wire y2f6a9k_hg3xfq93vb = gn916lc8_fzkp3rcqpob | a5s2gi2_h7rplzkx1;



  wire  bd3d3vhhigx1vbq1611n = 
        (d1rivbcy3w5oji6yoo & (~y2f6a9k_hg3xfq93vb)) 
      | (d1rivbcy3w5oji6yoo &   y2f6a9k_hg3xfq93vb & (j9o_ty1uw4uvham3ak == 1'b0));

  wire  rq6h3zj1i90esxh193v = 
        (y2f6a9k_hg3xfq93vb & (~d1rivbcy3w5oji6yoo)) 
      | (y2f6a9k_hg3xfq93vb &   d1rivbcy3w5oji6yoo & (j9o_ty1uw4uvham3ak == 1'b1));

  
  wire zs3i7m0dyc2b141ctfd;
  wire ee0lpnrpb0r5ezcvewy2 = ~zs3i7m0dyc2b141ctfd;
  wire q1t052cryjx59v5egpcc = (m2s492eolz_a4lrc == yjbrpsqyidt47leh_[1-1:0]) & o0nkaxltg92zc7_vvacwa;
  
  ux607_gnrl_dfflr #(1) gnezozmg7lduup3e_4m7un (q1t052cryjx59v5egpcc, ee0lpnrpb0r5ezcvewy2, zs3i7m0dyc2b141ctfd, gf33atgy, ru_wi);
  
  wire [1-1:0] gf0dpof_3vhwojox7c; 
  
  assign gf0dpof_3vhwojox7c = q1t052cryjx59v5egpcc ? 1'b0 : (m2s492eolz_a4lrc + {{1-1{1'b0}},1'b1});
  
  ux607_gnrl_dfflr #(1) uy4yu6hr_sw1839o33a2o7 (o0nkaxltg92zc7_vvacwa, gf0dpof_3vhwojox7c, m2s492eolz_a4lrc, gf33atgy, ru_wi);
      

  
  wire ovtnp77z94fvwwlmanp3m;
  wire ag1q8n1v0zdb0gd3mwnw = ~ovtnp77z94fvwwlmanp3m;
  wire aiadz_ucvzjlnyxt9c89_n = (j9o_ty1uw4uvham3ak == yjbrpsqyidt47leh_[1-1:0]) & oyc0vwbyun6num5qh;
  
  ux607_gnrl_dfflr #(1) jq3l62vfp3gv2vt48iaybpkho (aiadz_ucvzjlnyxt9c89_n, ag1q8n1v0zdb0gd3mwnw, ovtnp77z94fvwwlmanp3m, gf33atgy, ru_wi);
  
  wire [1-1:0] qda6sxg6ahx9dx7i5aio; 
  
  assign qda6sxg6ahx9dx7i5aio = aiadz_ucvzjlnyxt9c89_n ? 1'b0 : (j9o_ty1uw4uvham3ak + {{1-1{1'b0}},1'b1});

  ux607_gnrl_dfflr #(1) usdl9tgo_xp88gt90i85 (oyc0vwbyun6num5qh, qda6sxg6ahx9dx7i5aio, j9o_ty1uw4uvham3ak, gf33atgy, ru_wi);

  assign hy9lwz17ce = (j9o_ty1uw4uvham3ak == m2s492eolz_a4lrc) &   (ovtnp77z94fvwwlmanp3m == zs3i7m0dyc2b141ctfd);
  assign vvzs4gmapk7c  = (j9o_ty1uw4uvham3ak == m2s492eolz_a4lrc) & (~(ovtnp77z94fvwwlmanp3m == zs3i7m0dyc2b141ctfd));

  wire [1:0] jm4__y98e00ukvb4hiw_f = {eca4wu5z1eltuvtu76r7ti6, ctqj_dyrttnfzu9lcud3g_3};

  generate 
      for (i=0; i<yy567yahzg; i=i+1) begin:z8ha13bq2e55zoce36tle
  
        assign merfg1jkbwck[i] = o0nkaxltg92zc7_vvacwa & (m2s492eolz_a4lrc == i[1-1:0]);
        assign x974z3fncltxj[i] = oyc0vwbyun6num5qh & (j9o_ty1uw4uvham3ak == i[1-1:0]);
        assign hh2n5p_74cpa[i] = merfg1jkbwck[i] |   x974z3fncltxj[i];
        assign yo_tvqeum32rvou[i] = merfg1jkbwck[i];
  
        ux607_gnrl_dfflr #(1) c8n9altpe31o39ukpce (hh2n5p_74cpa[i], yo_tvqeum32rvou[i], trycoh_sgdgtcdg[i], gf33atgy, ru_wi);

        
        ux607_gnrl_dfflr #(3) m1ll7trcvgevi0m7oz8s (merfg1jkbwck[i], jgfckxgs0fo048, nyrioysq5ovac5r8[i], gf33atgy, ru_wi);

        assign iv9dhbb1gs4h19y[i] = jm4__y98e00ukvb4hiw_f[i];
        assign k8b8v2d_8bexygcseus[i] = x974z3fncltxj[i];
        assign cj_amdiu4_4kyqh[i] = iv9dhbb1gs4h19y[i] | k8b8v2d_8bexygcseus[i];
        assign bcohnzslp6bf6pqn1[i] = iv9dhbb1gs4h19y[i];
  
        ux607_gnrl_dfflr #(1) i0y9y21w9l9y4kflfhvjkp (cj_amdiu4_4kyqh[i], bcohnzslp6bf6pqn1[i], xlnalzy_jsdbs[i], gf33atgy, ru_wi);


      end
  endgenerate

  wire [3-1:0] n7fwy8f483ujgu2d = nyrioysq5ovac5r8[0];
  wire [3-1:0] qs3f0sj6kmhi5nn = nyrioysq5ovac5r8[1];


  assign k6uqslf4yjz0 = oyc0vwbyun6num5qh;
  assign ibegorpv3fon9ktf = j9o_ty1uw4uvham3ak ? qs3f0sj6kmhi5nn : n7fwy8f483ujgu2d; 

  assign i2hiwgez7xp0bc_3mg35a4rb = zsp7u2uqvojc8zqnw0k6_p & (~m2s492eolz_a4lrc);
  assign aq3hy9uuv5rnvzphrnaa3 = zsp7u2uqvojc8zqnw0k6_p &   m2s492eolz_a4lrc ;
  assign mljh30sszwrhguqyc4f5e77l4  = m2s492eolz_a4lrc ? rho1guu79090z97aekm9s16pn : lwl5fn5x_gxnq3f3a1tt0qyrd;

  
  assign yp6atu2uzbb053onf7h7j_g3 = lszyvs15rstcbyhj96v090d | qpzxk_hrtmppd7i7eplel;
  assign gl9dazcghkmei56i8tlb     = lszyvs15rstcbyhj96v090d ? iqj11baw8n07djxz1m45yxd     : z85m6lb5ii_p8z196b1r    ;
  assign k7x2rdsdsxkmoiyluje7bf2aa = lszyvs15rstcbyhj96v090d ? wx_fs2ijrykfgpoqldrgukw : zg97ncjhsfhaqpc60t6wfdr;
  assign j1utgrdwzlhqppb8rev5pbh55   = lszyvs15rstcbyhj96v090d ? tfwuip_0npwfy19ek9gpoc   : h987z8usv7pyyl5zqvzw4  ;

  assign gwy4w6j_23g_d3t     = haaqh6wjlwi9jhnl    [n7fwy8f483ujgu2d];
  assign xknh2ut7lctvrugsz5wb     = qp1mbsaizjipsj6    [n7fwy8f483ujgu2d];
  assign g3itms8el25jimpco2t_yu4     = a2oenic4uandesr_k9qocfw    [n7fwy8f483ujgu2d];
  assign w_fuqyygyv_7yus0ow9k    = vsfpyprm4rivny0n4   [n7fwy8f483ujgu2d];
  assign ld964zre2gsugp9blpo    = zrhld0y35qav   [n7fwy8f483ujgu2d];
  assign h5986karddzxifsa9t    = xzc0imuvetgbn8   [n7fwy8f483ujgu2d];
  assign ya7g9x7j5jke20pxxk    = halyb9c30hal   [n7fwy8f483ujgu2d];
  assign hyiwh018ufcuat94ohr4    = pllepw4azlfujoh_i   [n7fwy8f483ujgu2d];
  assign mdw031z1stmwv1atvh9pla6    = d1rzzdht0dlkdfjvs420q   [n7fwy8f483ujgu2d];
  assign kqe4mxh6t85yt1es15h_kv3y_    = hwwn5fuw1ki6rpxis   [n7fwy8f483ujgu2d];
  assign eidxuo2trad883370opeq    = v1bfb0aqght1_yfm5znt   [n7fwy8f483ujgu2d];
  assign yz4xms1_6ldn__afmhfdxic = knyt1bhi0tp16v3[n7fwy8f483ujgu2d];
  assign k6aoxxoxugbmismespiv2pfhf = fizjb37qgnqc11y3usvo1jd8[n7fwy8f483ujgu2d];
  assign g6zc5qflpket_8b_30jviei4n = te3sgyqybgiz02r496eiram[n7fwy8f483ujgu2d];
  assign ff8kz54m27i8p1qxp4c_n1y = hotgsfmzxnfg6u691gfcuem[n7fwy8f483ujgu2d];
  assign lm8vcj797bp12bltgigc6lk76ei1 = dej8khi216rqhe3ebb4[n7fwy8f483ujgu2d];
  assign cnh34kai5koa_4iw5boo0p = bk8m_k0vayvzu1ytxtuvky[n7fwy8f483ujgu2d];

  assign xnmq3kuajinzxdfiu6q     = haaqh6wjlwi9jhnl    [qs3f0sj6kmhi5nn];
  assign xdheobtph1wq8f9ui3h     = qp1mbsaizjipsj6    [qs3f0sj6kmhi5nn];
  assign nni92t4rn44yvbfgt5yor94mh     = a2oenic4uandesr_k9qocfw    [qs3f0sj6kmhi5nn];
  assign rft88ds492cdh634i    = vsfpyprm4rivny0n4   [qs3f0sj6kmhi5nn];
  assign u87rvzwj0xs9vt8uwuot    = zrhld0y35qav   [qs3f0sj6kmhi5nn];
  assign wawfribsksiyhybl3m1fc    = xzc0imuvetgbn8   [qs3f0sj6kmhi5nn];
  assign zfmqdobuh7r4t0fza5uv    = halyb9c30hal   [qs3f0sj6kmhi5nn];
  assign jhiyy3sgiaizu4l4milff    = pllepw4azlfujoh_i   [qs3f0sj6kmhi5nn];
  assign snm9n0s_9re1n13_p9tec    = d1rzzdht0dlkdfjvs420q   [qs3f0sj6kmhi5nn];
  assign ccf5m6bnqnibseotadeyu86cd0    = hwwn5fuw1ki6rpxis   [qs3f0sj6kmhi5nn];
  assign irncno4zcb4x06mlfiba16bh    = v1bfb0aqght1_yfm5znt   [qs3f0sj6kmhi5nn];
  assign yc59czg2u_bbaxbn1ejpjm8w = knyt1bhi0tp16v3[qs3f0sj6kmhi5nn];
  assign n3r6ftigei07xsagxiifpct = fizjb37qgnqc11y3usvo1jd8[qs3f0sj6kmhi5nn];
  assign j8lpsrktt_qs_wo43c_rre4 = te3sgyqybgiz02r496eiram[qs3f0sj6kmhi5nn];
  assign ryz4vgf7dpx5dcq733ch1f5gm = hotgsfmzxnfg6u691gfcuem[qs3f0sj6kmhi5nn];
  assign ulggxuvjbou5t00s_czahip80ud3 = dej8khi216rqhe3ebb4[qs3f0sj6kmhi5nn];
  assign kbt5xarx9to2rj956ik1zwwq = bk8m_k0vayvzu1ytxtuvky[qs3f0sj6kmhi5nn];

  wire                            agnsw48g8fdikd;
  wire                            x25ltyb13sb2td2;

  wire lt23vkvcmjwt0_0j           ;
  wire jrxv7dijvw894k_vlv2lhga    ;
  wire t7kciau00u9xy6cb157ewa429m       ;
  wire cw53t17pm78oskoyt49oivc7qh3ab8;

  wire                               o3ydhguk119jyhp47x106ib;
  wire[32-1:0]          enqm3v278hn097pt6_04p9n;
  wire                               hs3xn0evnbpy575ea7p5p3qto53;
  wire                               sycglehz7v8eijxjqe7ufoxp4j1y;
  wire                               pihkjnbghw4bk8y2477x7k82o93ug;
  wire                               crriagr_kegsjfrtly_v8yw9;
  wire                               p5u44x4jrltstcsbmk8kg5hnq0;
  wire                               ve1mua6_hp7e4a8tf03lfitualb;
  wire                               m7fr__lszd5b56qf13pbarusep;

  wire                               gg0tr7jpfos4ct46rnx8kikun5t6ee;
  wire                               vfxj481iib57qmfew_ggqin2rqaa;
  wire                               tl82sx3puyxv5f6eoxlnfunqhe8;

  k7eqwfmolitp9my9g4 vypajg4xg8j7p72(

    .hv39pppvbmeqy8b6        (no360dfthc_r812ltoqdhrz       ),
    .dukd0zozp1ektzmt7f        (o3ydhguk119jyhp47x106ib       ),
    .t6l88yqbe4wokkhiso9t       (enqm3v278hn097pt6_04p9n      ),
    .hyec__ebnw8lbcssd81       (hs3xn0evnbpy575ea7p5p3qto53      ),
    .vs2610q9_on1r996p      (sycglehz7v8eijxjqe7ufoxp4j1y     ),
    .coy3buxdw6yq3duh21azuwflk (pihkjnbghw4bk8y2477x7k82o93ug),
    .r_8h5lxb39ug57zli04e_o      (crriagr_kegsjfrtly_v8yw9     ),
    .pv7q0ikpayogkay57rgyr      (p5u44x4jrltstcsbmk8kg5hnq0     ),
    .dsq8f3rhmb7yc876v8     (ve1mua6_hp7e4a8tf03lfitualb    ),
    .enu_vumk17eoj1fma5ilz0    (m7fr__lszd5b56qf13pbarusep),
                             
    .ou74jmm5p6th0y0kcdwpqv2ey (gg0tr7jpfos4ct46rnx8kikun5t6ee),
    .adwzzx09c_s_x1seh      (vfxj481iib57qmfew_ggqin2rqaa     ),
    .zp0aylmm0k4yw4w561bgzh    (tl82sx3puyxv5f6eoxlnfunqhe8   ),

    .kd96ha16hcj4wyo0          (tq5w2fd0flcywep677l  ),
    .j9kszxa35hle0cl9         (k6_e3_saw0oup16pudov ),
    .myqlprv648_pqf92vvj        (zpq6nysk8b654ynyt4zj9k),

    .zpdvh58o0evhzt           (lt23vkvcmjwt0_0j           ),
    .q0duv6epk3ccff620vhhx2    (jrxv7dijvw894k_vlv2lhga    ),
    .rpkosm9pbcpggwup90_ge9       (t7kciau00u9xy6cb157ewa429m       ),
    .xwmkl_9n7oehwe7hh_a6aompojzukuik(cw53t17pm78oskoyt49oivc7qh3ab8),

    .z8alxhlwgz117             (z8alxhlwgz117), 
    .q4j831gvqooep12             (q4j831gvqooep12), 
    .tyg8z9t16af4e8xtdiw       (nl2n_jy0ye9rq9j0hteu),
    .qkl9_olndwlohzaurunzkg       (xerurm1znxab6ednf5rf),

    .fpihselr34pn79               (ye2fnsl_jl2n9kk6               ),
    .jm4__y98e00ukvb4hiw_f        (ctqj_dyrttnfzu9lcud3g_3        ),
                                                         
    .w4sit6hoc28giqb51t3n6       (i2hiwgez7xp0bc_3mg35a4rb       ),
    .tbli88os0gfvjlfl6ttv1       (lwl5fn5x_gxnq3f3a1tt0qyrd       ),
                                    
    .hxvldlso5zpp81            (gwy4w6j_23g_d3t            ),
    .ahhi0t6w86wbz891shq            (xknh2ut7lctvrugsz5wb            ),
    .zkqavy8j9jzdikz_29v7am     (g3itms8el25jimpco2t_yu4            ),
    .bl79n71wkynirgcs3           (w_fuqyygyv_7yus0ow9k           ),
    .o8smcfmzt25hxpwcn           (ld964zre2gsugp9blpo           ),
    .y4tsxz4rprpynubw3rvm           (h5986karddzxifsa9t           ),
    .n7jh1zclcr_s0l4bgd           (ya7g9x7j5jke20pxxk           ),
    .wunjscg6om1d0yu8o           (hyiwh018ufcuat94ohr4           ),
    .f24hbj6y6nq5sy45lqzm5s           (mdw031z1stmwv1atvh9pla6           ),
    .od57enqth4m5g9lpdduxdx           (kqe4mxh6t85yt1es15h_kv3y_           ),
    .ibt51xz_a6yo4yknr5mx1      (eidxuo2trad883370opeq        ),
    .vqfoysp81h8x_kvfv1sg56        (yz4xms1_6ldn__afmhfdxic        ),
    .l03z9wtep77xkwohwq0e_1lm     (k6aoxxoxugbmismespiv2pfhf        ),
    .e4wqef4o71wrrp_crj0dw8     (g6zc5qflpket_8b_30jviei4n        ),
    .eymxkl1knoowfwizivwrzpsi     (ff8kz54m27i8p1qxp4c_n1y        ),
    .rbrj5qqhjrxh023fhy4v2ce     (lm8vcj797bp12bltgigc6lk76ei1        ),
    .xdyys2soinatq_bm7r2g35ie     (cnh34kai5koa_4iw5boo0p        ),

                                   
    .yp6atu2uzbb053onf7h7j_g3      (lszyvs15rstcbyhj96v090d      ),
    .gl9dazcghkmei56i8tlb        (iqj11baw8n07djxz1m45yxd        ),
    .k7x2rdsdsxkmoiyluje7bf2aa    (wx_fs2ijrykfgpoqldrgukw    ),
    .j1utgrdwzlhqppb8rev5pbh55      (tfwuip_0npwfy19ek9gpoc      ),
                                                          
    .rinamilgle00i5xmx_vt        (bidjco9v6uwp91tvsqnp72df_u0q        ),
    .j8wlfupbw25hdmohz5q0        (m83gf40i8n5qmmo860pq3w7n5n5f        ),
    .z64bwdr23steb7s9y9j         (q064m0tgrtkrz7vn_qf2bjb         ),
    .bg1spy6_v2kbo75pz1d6         (xxrb4v2suklf9djaeyf0rkmedjz3         ),
    .xyeq7c6icdac80_y0jup        (hrn1giqg1k6gbt6q7lrxzxaqztx        ),
    .za5ms2soyuucfxo_jbn        (xw04i4vzqgn2m2ihbdv55m4bvtr        ),
    .b7aet1zp_fcfxn8h7rw0u1        (h_9b0wqhlkmvxkfizht97cqp        ),
    .t3szwnvfo2nj3wk6r5kvt         (ycmo1kcbjq1scw4gwg4uiwd_         ),
    .m4x1_gvw8v_sc8h7c8_6         (ocdu63ksnvvgacaermakucm0f4g         ),
    .hpeqnhpztp9l_d3yx16l         (oxlxxz2rxp0amufq1s9jqrry3y         ),
    .bngbyv57e7juc0vkk2y8i         (rcpyv929ixr6xhyeyg2p0cgtj         ),
    .cneu8a119tg3vmie6zr2h_        (n169ohp8pq9l7goaugowzjfa        ),
    .jw2dzv9gi7gygudyqql6fz        (psec5ihpqk4slg2u90eq4yzyy        ),
    .o_7kpry6inkqpqi1bf1nd        (cv6960ns7f2dyrvj6ij_phb0        ),
    .f97tgz_qybmvln6nz5dqt458       (kxqipwn8s_54dje1dpjvcgaye6t       ),
    .znotwr53pu47f5m1agm           (gc_aq81uy3hbdq8ns7y1_ckg           ),
                  
    .zf_v02okbs8_euhd64        (vkjwr2hxue8911qmv5ro35cg        ),
    .wq4r8m45isqp8_o4pdtitz        (xronfobw50555i02avvye82b        ),
    .qpzo6lin6brrytho7         (kbbc76s46hvu_3te0ihj3hb2nl         ),
    .k7j6g0757jovg8xstgrvwf         (g33u_ys44gmrebks2nd9y8o         ),
    .nwx86gohbrn08nvh60789        (y5gfh4gmog9i5iq47qq3nmc95_fnd        ),
    .bebhplbk2k43sfoehvt66w        (bafx6nbdipfv60zavyhkpt5ulfqp        ),
    .ljk3q52m5tirt6shbcwbf        (wfq3yog1gp3v5k8ew8aazeio5q9qm        ),
    .ucj9poqgl683ej1pihkh         (bkec53bqczw0o6vx2ouxlbp         ),
    .u9hi0xtx8u0mn0l_7p         (o347ncxtm6aeg09kb47k1oggzcw         ),
    .rm04yhu6ondli9u0g6din         (pfkm_ekt4p23xk05wj0f5ei8wut2         ),
    .o5fmtstd7kef7z4m7jefm         (rx7d01wkjl49umakx8rnira0bvj         ),
    .vvadj6ew1h5wq9z5askkzr9        (bpetbkuwyy1k6fa142bfw3rz7sjpi        ),
    .lop06h0_z_4tt1s04up        (vsn6zt6npfa5qvbab0qrm7ya        ),
    .ivllgcn1kiix2iamzwf0u        (c_saxxol2d2vxelssdxtjul5uxmn        ),
    .rnmvpk356vfgxd_045g       (yueav99q0b7x3rcm9_x625j6yd       ),
    .a46c4xo4texvc9o           (c7y5emtdpd3rk_dus5ixb7r44           ),
                 
    .ze2bfnigu62i9937pcxnjc        (xnvidl2ouve1vln7ywwu6a5v        ),
    .c86b14qr2qo45_qw2ns        (k0ue65kc80maq9qkm04zau8h4bz        ),
    .dm5b92mx0redfbuhs1u3d          (we3r29j8uhskq7kyw558l15b7          ),
    .c4cb28s8l8rdx2e53vww      (vsf0g6h63ew3evcsozmlfhinvhq      ),
    .c3vtv1izxu7rm5646jsmmke        (yzi326ahunke54273wsh5pgc7kka        ),
                
    .mm70cenjp_1wmcs135nh4wl        (qp6hat5pdku7yc9bq1vsm6hb_w9        ),
    .p4dpiqc4w_g42ni5jsaj        (n0pfd6t_58aep4y4wg7wl9vo7ejyz        ),
    .ezntrtg3q1must0tfcgn          (f1t_hrt88trjzo1oeoj3ui9lhcu          ),
    .h99vs7dtnw2w96vts56dhc2      (qah4iiv5ntbmab46ir87_rkxcqzih4      ),
    .glqyhrpm6zzwddhsd6mcd1u        (nud3tr5ire99qpl6xy6s2vj0        ),
               
    .c9oejgc5s6_v8ooyy8c0x1          (khbwxlyuzlnl1c8t8_3og_5mq          ),
    .sktjnm1h7yu59cy6lnbf0gx40e_     (qnthfit20wgbpxec8thtex71gzm7     ),
    .izozgg91hphikoatw0xsa         (ddrezcee7228fcb3xe5ptlosy         ),
              
    .m7rpuph0hm25ukmyralijiy          (hystveyc5mdp2fsv1prg          ),
    .r_13gm13ck84al5d7ty5lf_m     (cqnseh0h9l57x_6_lagpk2_zv     ),
    .ck7dirv94s9jkefjfed0h0mp         (zi8qhl5upl3l4fr_x69d9         ),
              
             
    .jkq984ky8fozrzq               (on12sjnlw0b975rtxnj),
    .g3_8p4g7w5grnl62xy            (m91uirvkay9adfjui930dyv4            ),
    .vqwqaofc8sz_yjccd            (a_i3c4odzkmjpufk2pffcu            ),
                               
    .tyxs3jzhr2i2gq9dt7            (i691bnr_y8gmwnd0nsaw            ),
    .zti98n829owa2p            (isqt1ng7lccfet8bj5hym5c            ),
    .ye256knohacnaakiw2nqck6     (ije4h78_umvknjj6az4_5qf92e3iydh),
    .hyxeikuobvxjumz2hibay     (sro97_d1rgt1fmqi2b_fitscvexczye2),
    .zkojor8433oflab2kpvtzi1z9     (v2tse065uysfbl8f4z8hlpkg5o68     ),
    .nx6i4o0_cbqmlan1ylpodj9y     (kwczwxezdeidftn2_p2fpzik3gt     ),
    .tgfv2w2s7qhwkl0pdpf_79v4e     (o58xzacx8hg_9zcqk21v9m0rqqsap22_     ),
    .qfjl6250hpfb57pxl0t53q6fd     (q0xni3yf49f2fj7ymo_nvdurqx1okyv     ),
            
    .j2kcz1faqhvh1ler6j           (rbkhb89tyu_ucjpo           ),
    .a6gdkt5h77dh0mcj8t4gq         (sqvgnqdrkexeg2lziofadt         ),
    .wixbtbeqlhzelg4t           (bwtzw5pqhc62g9v9w           ),
    .uh_ekyw7cw8c3d3xj1          (nwbvll63g8yq6vbpxok          ),
           
    .uf44audysjgtvdnua67           (e4ui35hoxqcwkgfaol           ),
    .qtcasxm90cy0bwaqaxz         (f1uy000fu6355gukzxt9r4y         ),
    .y38seii6ja77q2jy08           (avudrqvyzx1dringrt4rs           ),
    .f42g8ulc2y43ntmai5          (hz5leo9sklh2v25_50          ),
          
    .cgnsvvj7srbljqst             (agnsw48g8fdikd             ),
        
    .rgf8pa4kn20jusruz           (ofg0te04_oeiba586           ),
    .wjwjffxr_4lulivwz         (dm0uaanzcp_7hojw2_h         ),
    .z6udkjbx164gh9yo1o          (yddyulfbyf7p2wvl6dyk          ),
    .frkunk72hlttw0ar0np          (j233e_ya9xhnxg7flb9d3          ),
       
    .r2tvaf8px0p9vlw4we           (mq3a_g7zrfyfdil1           ),
    .srfn4smswwo6hbyaa         (f9ekxi98w3bnnfm3t1vyt1         ),
    .a_u2kfmgv2ho357c          (k1vhaduoq3xy5cx6jr0          ),
    .svj88sv2u56fepzmg          (hwo9njh5b4299teslcl          ),
      
    .rzf167thmprvps0tm62i           (shxdziymfk57c49e0           ),
    .lv7fu0hif2n2zhmgtcc         (s_fatq1jfpqkf7q9d40n         ),
    .oj5t3f0lq1n9ae82x          (ruix76vs69a8gynr7yydnp          ),
    .hat38salswlktk821          (y0s6zoimyz170437bgkne          ),
     
    .caxkrdjq0tjnnne9           (nsyif4pw3tzuggdakg2           ),
    .qpuk8ry0w9_r7ur4gcnx         (e4zsuzpz_sgcgql5k19iv         ),
    .v8jl1eh8o0n5g765          (fvzgpoei5_ffhtrv6r          ),
    .c0xnu9p8he2hw10h          (cnqt629_5e9xaypczfdt          ),
   .gf33atgy  (gf33atgy  ),
   .ru_wi(ru_wi)  
 
  );


  wire d0vr59qnksmk5qmvaie           ;
  wire v2hd81fxe604639r8kl8oye90    ;
  wire e94jesry36znm45r1soyhic0hk       ;
  wire zgp64zvc52r2j6zasb74b8wzx6nm68icc6;

  wire                               b4687t39adr64eo0i4lf5md;
  wire[32-1:0]          fsgnhdgr565rvtm7jewinuufhjm;
  wire                               ilmemra32cftf81jy7tb1tn;
  wire                               p8rx6454dkq9mcu0knbdrp4;
  wire                               oy5tnom44u2vm3zpklpy9_xsje_dh;
  wire                               enjo_thzs5fjl2yaorgzrh85sivo;
  wire                               eg3xuv8r03e6j0msnfyr8i2b;
  wire                               kc_oc1b1x6hj408h8pkuuwr09qnr;
  wire                               zjp7e4i7qt_0abds5ihh_dnqk;

  wire                               ydi3gh_3ks81b74d8g9vgn081jicdv8;
  wire                               ce_6thxzv8n4n8xdhg9y9ftl;
  wire                               xg81tsg3z29z7lie1domdmt86crlg;

  k7eqwfmolitp9my9g4 mifteg5b2oci7z4zj(

    .hv39pppvbmeqy8b6        (piosx1_uvpor01vn8ll66_yhit       ),
    .dukd0zozp1ektzmt7f        (b4687t39adr64eo0i4lf5md       ),
    .t6l88yqbe4wokkhiso9t       (fsgnhdgr565rvtm7jewinuufhjm      ),
    .hyec__ebnw8lbcssd81       (ilmemra32cftf81jy7tb1tn      ),
    .vs2610q9_on1r996p      (p8rx6454dkq9mcu0knbdrp4     ),
    .coy3buxdw6yq3duh21azuwflk (oy5tnom44u2vm3zpklpy9_xsje_dh),
    .r_8h5lxb39ug57zli04e_o      (enjo_thzs5fjl2yaorgzrh85sivo     ),
    .pv7q0ikpayogkay57rgyr      (eg3xuv8r03e6j0msnfyr8i2b     ),
    .dsq8f3rhmb7yc876v8     (kc_oc1b1x6hj408h8pkuuwr09qnr    ),
    .enu_vumk17eoj1fma5ilz0    (zjp7e4i7qt_0abds5ihh_dnqk),
                             
    .ou74jmm5p6th0y0kcdwpqv2ey (ydi3gh_3ks81b74d8g9vgn081jicdv8),
    .adwzzx09c_s_x1seh      (ce_6thxzv8n4n8xdhg9y9ftl     ),
    .zp0aylmm0k4yw4w561bgzh    (xg81tsg3z29z7lie1domdmt86crlg   ),

    .zpdvh58o0evhzt           (d0vr59qnksmk5qmvaie           ),
    .q0duv6epk3ccff620vhhx2    (v2hd81fxe604639r8kl8oye90    ),
    .rpkosm9pbcpggwup90_ge9       (e94jesry36znm45r1soyhic0hk       ),
    .xwmkl_9n7oehwe7hh_a6aompojzukuik(zgp64zvc52r2j6zasb74b8wzx6nm68icc6),

    .kd96ha16hcj4wyo0          (juwj_oo3r8yt2a4hg  ),
    .j9kszxa35hle0cl9         (pzfb_24lrjd770iigjx4sm ),
    .myqlprv648_pqf92vvj        (d2lstp52x9w9900ioarrtfk),

    .z8alxhlwgz117             (z8alxhlwgz117), 
    .q4j831gvqooep12             (q4j831gvqooep12), 
    .tyg8z9t16af4e8xtdiw       (bvwt0k4qftqv4to2lj6d46_),
    .qkl9_olndwlohzaurunzkg       (ocz7civlapwkb3oe78oqt2fw),
    .fpihselr34pn79               (mvkoyonaqzuf3ip               ),
    .jm4__y98e00ukvb4hiw_f        (eca4wu5z1eltuvtu76r7ti6        ),
                                                         
    .w4sit6hoc28giqb51t3n6       (aq3hy9uuv5rnvzphrnaa3       ),
    .tbli88os0gfvjlfl6ttv1       (rho1guu79090z97aekm9s16pn       ),
                                    
    .hxvldlso5zpp81            (xnmq3kuajinzxdfiu6q            ),
    .ahhi0t6w86wbz891shq            (xdheobtph1wq8f9ui3h            ),
    .zkqavy8j9jzdikz_29v7am     (nni92t4rn44yvbfgt5yor94mh            ),
    .bl79n71wkynirgcs3           (rft88ds492cdh634i           ),
    .o8smcfmzt25hxpwcn           (u87rvzwj0xs9vt8uwuot           ),
    .y4tsxz4rprpynubw3rvm           (wawfribsksiyhybl3m1fc           ),
    .n7jh1zclcr_s0l4bgd           (zfmqdobuh7r4t0fza5uv           ),
    .wunjscg6om1d0yu8o           (jhiyy3sgiaizu4l4milff           ),
    .f24hbj6y6nq5sy45lqzm5s           (snm9n0s_9re1n13_p9tec           ),
    .od57enqth4m5g9lpdduxdx           (ccf5m6bnqnibseotadeyu86cd0           ),
    .ibt51xz_a6yo4yknr5mx1      (irncno4zcb4x06mlfiba16bh      ),
    .vqfoysp81h8x_kvfv1sg56        (yc59czg2u_bbaxbn1ejpjm8w        ),
    .l03z9wtep77xkwohwq0e_1lm     (n3r6ftigei07xsagxiifpct     ),
    .e4wqef4o71wrrp_crj0dw8     (j8lpsrktt_qs_wo43c_rre4     ),
    .eymxkl1knoowfwizivwrzpsi     (ryz4vgf7dpx5dcq733ch1f5gm     ),
    .rbrj5qqhjrxh023fhy4v2ce     (ulggxuvjbou5t00s_czahip80ud3     ),
    .xdyys2soinatq_bm7r2g35ie     (kbt5xarx9to2rj956ik1zwwq     ),
                                   
    .yp6atu2uzbb053onf7h7j_g3      (qpzxk_hrtmppd7i7eplel      ),
    .gl9dazcghkmei56i8tlb        (z85m6lb5ii_p8z196b1r        ),
    .k7x2rdsdsxkmoiyluje7bf2aa    (zg97ncjhsfhaqpc60t6wfdr    ),
    .j1utgrdwzlhqppb8rev5pbh55      (h987z8usv7pyyl5zqvzw4      ),
                                                          
    .rinamilgle00i5xmx_vt        (flb64u531jaudptz5l9y7ju5        ),
    .j8wlfupbw25hdmohz5q0        (so7wnp3pfxe74elogsol7qrvj_5        ),
    .z64bwdr23steb7s9y9j         (z6x6vtfm5ozsb8e1g3ek9mxcaavx         ),
    .bg1spy6_v2kbo75pz1d6         (nsvtf_9m6sep1hb1kltgl2hlnqn         ),
    .xyeq7c6icdac80_y0jup        (odd4wynvno2o6hjyvi65l10zi        ),
    .za5ms2soyuucfxo_jbn        (zbpyr_m9c2hqfkc019qkpou4krbxw        ),
    .b7aet1zp_fcfxn8h7rw0u1        (l0tlr34v20v3hk8a6gie4uk91yp1w        ),
    .t3szwnvfo2nj3wk6r5kvt         (riimr6qwir1dx_guosj51l91         ),
    .m4x1_gvw8v_sc8h7c8_6         (szfy9s6lzimlb2j3cs5_vlwl         ),
    .hpeqnhpztp9l_d3yx16l         (vqq0vkkbq8gqc1tz1k_ud7rm42za         ),
    .bngbyv57e7juc0vkk2y8i         (frs0vh2vwgovicyibkf_d3sr6_         ),
    .cneu8a119tg3vmie6zr2h_        (x7bhi63pp_k_4diubx18eq_x6c        ),
    .jw2dzv9gi7gygudyqql6fz        (vmucahlss7dpuvf0zo7r14es8mw4e        ),
    .o_7kpry6inkqpqi1bf1nd        (j46f_ypuqx8_ubhj2dqsl2nvo3xl2        ),
    .f97tgz_qybmvln6nz5dqt458       (s5m9cu2ee3zjqralllxvdcnv_nr       ),
    .znotwr53pu47f5m1agm           (hycfweaqoatse84iuu9rp           ),
                  
    .zf_v02okbs8_euhd64        (lxdia3j_hv2zwfjcp0_5bnsv3xu        ),
    .wq4r8m45isqp8_o4pdtitz        (kf17agt2l21y8meszqlaks6n        ),
    .qpzo6lin6brrytho7         (w2rebtphwb45_nf6qw5dy26z         ),
    .k7j6g0757jovg8xstgrvwf         (ypdw34_kup0gaiwjzl4bcthak         ),
    .nwx86gohbrn08nvh60789        (yg5d3o1ke2l9iz9fexcwz4ndh        ),
    .bebhplbk2k43sfoehvt66w        (t43psmvm15g070eibanybptz7        ),
    .ljk3q52m5tirt6shbcwbf        (wz17_6fsan5b1vvg2gbkburw2        ),
    .ucj9poqgl683ej1pihkh         (wbp0e817xt2uj0bm5047co29g9jr         ),
    .u9hi0xtx8u0mn0l_7p         (kzneydeew74np7qbndwhvw_         ),
    .rm04yhu6ondli9u0g6din         (rywjhkc2m319gtnl68n6yia0h         ),
    .o5fmtstd7kef7z4m7jefm         (xqr6qbo6fxrb8hni14at1bkd1o         ),
    .vvadj6ew1h5wq9z5askkzr9        (rr_kd00n0nzd08jhv6de62tu5w2e        ),
    .lop06h0_z_4tt1s04up        (ci_vdf2vqsfb45ipjbbj2kf0g        ),
    .ivllgcn1kiix2iamzwf0u        (cm2iw9jkt_zvly6ri5f7s0sz3q        ),
    .rnmvpk356vfgxd_045g       (r048om6_elh04xzuybqp1x5ynfs4um       ),
    .a46c4xo4texvc9o           (zjg4nl981npxovpev0e_yqz4           ),
                 
    .ze2bfnigu62i9937pcxnjc        (duzcgyd7bbw3jp7bax5m_im68gt        ),
    .c86b14qr2qo45_qw2ns        (w0414mghkbrhfheu2cmwalfj9g0        ),
    .dm5b92mx0redfbuhs1u3d          (ibfxlpjz4f428kdyrvz2l243b__          ),
    .c4cb28s8l8rdx2e53vww      (zdq146b5sl9b_zsw84kq0l8u51ph      ),
    .c3vtv1izxu7rm5646jsmmke        (b49a3gf23ov9g7xpe88_11si96vh        ),
                
    .mm70cenjp_1wmcs135nh4wl        (rwfis2p5oqcxun3vrabpu4ehd        ),
    .p4dpiqc4w_g42ni5jsaj        (ssgsllp8a48t220i6zawign01kjs        ),
    .ezntrtg3q1must0tfcgn          (pb5hz9n6i21hdl1f9ktx2pf4s          ),
    .h99vs7dtnw2w96vts56dhc2      (gqcennvw7i4s9ra6nufl5auv9n2      ),
    .glqyhrpm6zzwddhsd6mcd1u        (zie7s8nvi9nxy9tbeenymedx2ch        ),
               
    .c9oejgc5s6_v8ooyy8c0x1          (kn4nyomkyc9nib4jk3q9v9u          ),
    .sktjnm1h7yu59cy6lnbf0gx40e_     (ms19_yn0emkdebo5xds5no7own3k     ),
    .izozgg91hphikoatw0xsa         (koyy03uze4eek43dncxyfucn2         ),
              
    .m7rpuph0hm25ukmyralijiy          (xirk22lqyoyt4_ojp1k3vkzye          ),
    .r_13gm13ck84al5d7ty5lf_m     (bo3wo9aretoipldnjadceyp2kgl     ),
    .ck7dirv94s9jkefjfed0h0mp         (li46sayiwuz6fbzu8n2xux         ),
              
             
    .jkq984ky8fozrzq               (a5s2gi2_h7rplzkx1),
    .g3_8p4g7w5grnl62xy            (gn916lc8_fzkp3rcqpob            ),
    .vqwqaofc8sz_yjccd            (nepu6mf61h2b2uewptpauek6v            ),
                               
    .tyxs3jzhr2i2gq9dt7            (xu6a8p2dk2fy9r7lnn_kd1l            ),
    .zti98n829owa2p            (pn1rzse3t9e6g_et37gv            ),
    .ye256knohacnaakiw2nqck6     (lwmr8fyosc4w78ftaznb17d0wep6),
    .hyxeikuobvxjumz2hibay     (g_lbo1t8r4bx4olr034dfi8fhfw1m6i),
    .zkojor8433oflab2kpvtzi1z9     (xmf6kblqlhyjpa44uj3tn_7hs9g     ),
    .nx6i4o0_cbqmlan1ylpodj9y     (td_dxcgpaod7g2fvddly_mg4rjh2vgbk     ),
    .tgfv2w2s7qhwkl0pdpf_79v4e     (l1mayxu6go0ni6a1uu2tn40qyps5l_     ),
    .qfjl6250hpfb57pxl0t53q6fd     (qdf9k5s3p4c0d8jxgmxlyi478ade     ),
            
    .j2kcz1faqhvh1ler6j           (idcribpugamfq_39t           ),
    .a6gdkt5h77dh0mcj8t4gq         (nfuf_njr73sjp5jr12d7gc         ),
    .wixbtbeqlhzelg4t           (hgm8yvqudk9e2ne6           ),
    .uh_ekyw7cw8c3d3xj1          (ivt9rgs2qqjzyrq5zt4isy          ),
           
    .uf44audysjgtvdnua67           (u6di3j5ypwgwjvnmcbsqh           ),
    .qtcasxm90cy0bwaqaxz         (i7vlo92n37lvcod6oj         ),
    .y38seii6ja77q2jy08           (ulp1cmdd07o0vc3p_65wi           ),
    .f42g8ulc2y43ntmai5          (f9_zg3c33q9sbq6d82u          ),
          

    .cgnsvvj7srbljqst             (x25ltyb13sb2td2             ),
        
    .rgf8pa4kn20jusruz           (mgc5k45s6iun0h64mg94n           ),
    .wjwjffxr_4lulivwz         (kuhd9_39ag_1mza9vf7x         ),
    .z6udkjbx164gh9yo1o          (dbp3mo7p_zh0242q9          ),
    .frkunk72hlttw0ar0np          (enbd230u3ab6jrd2gt          ),
       
    .r2tvaf8px0p9vlw4we           (nwvjy589molbkspazci           ),
    .srfn4smswwo6hbyaa         (hkv3jt_7_o_8sk0aait_0kp         ),
    .a_u2kfmgv2ho357c          (dzca_d1t69gei8viv2q          ),
    .svj88sv2u56fepzmg          (w7paq1qa9rrtadyr3v3cx          ),
      
    .rzf167thmprvps0tm62i           (ky3t5ldjtr_g__hnxr58s           ),
    .lv7fu0hif2n2zhmgtcc         (l20gjym8j9s2t31_nhs8iuh         ),
    .oj5t3f0lq1n9ae82x          (r3kh4eweep0kg7fak6rx6f          ),
    .hat38salswlktk821          (vwj6zdjeua22z66vj          ),
     
    .caxkrdjq0tjnnne9           (tbykhfjbcc3ure59           ),
    .qpuk8ry0w9_r7ur4gcnx         (v0oz07osad44us4h0pyd         ),
    .v8jl1eh8o0n5g765          (xtiqejiid_qbh90nn_jv          ),
    .c0xnu9p8he2hw10h          (dzoe86_fm7z7_c7_4_zn          ),

    .gf33atgy  (gf33atgy  ),
    .ru_wi(ru_wi)  
  );


  
  assign a03er8qo6p0zpb            = lt23vkvcmjwt0_0j     | d0vr59qnksmk5qmvaie    ;
  assign z8uuyp_3l6aqut86nkd__vvwgs     = (lt23vkvcmjwt0_0j & jrxv7dijvw894k_vlv2lhga) | (d0vr59qnksmk5qmvaie & v2hd81fxe604639r8kl8oye90);

  assign bzsjo5unerpy5i0e_q_6eqn        = t7kciau00u9xy6cb157ewa429m | e94jesry36znm45r1soyhic0hk;
  assign ctfhepdgvm53k59kbbe0s0924he0ijd = (t7kciau00u9xy6cb157ewa429m & cw53t17pm78oskoyt49oivc7qh3ab8) | (e94jesry36znm45r1soyhic0hk & zgp64zvc52r2j6zasb74b8wzx6nm68icc6);

  wire imzw3o6xtgdmikumc =  g3_8p4g7w5grnl62xy & vqwqaofc8sz_yjccd;
  wire yhwk19tompbv5zx = (tyxs3jzhr2i2gq9dt7 & zti98n829owa2p);

  wire bekul5xbo28zkmc90zy = (rq6h3zj1i90esxh193v & 1'b1) | (bd3d3vhhigx1vbq1611n & 1'b0);
  wire ap0oygari76txu48a;

  ux607_gnrl_fifo # (
   .CUT_READY(0),
   .DP(d8ba36mdzefszkfe3pwmzqxhwx),
   .DW(fumremxmy8mtkpij650zgfe79i)
  ) rdn_5jx1mqh6wucg6pbl0 (
   .i_vld(imzw3o6xtgdmikumc),
   .i_rdy(), 
   .i_dat(bekul5xbo28zkmc90zy),
   .o_vld(), 
   .o_rdy(yhwk19tompbv5zx), 
   .o_dat(ap0oygari76txu48a),
 
   .clk  (gf33atgy  ),
   .rst_n(ru_wi)  
  );


  assign i691bnr_y8gmwnd0nsaw = tyxs3jzhr2i2gq9dt7 & (~ap0oygari76txu48a);
  assign xu6a8p2dk2fy9r7lnn_kd1l = tyxs3jzhr2i2gq9dt7 & ap0oygari76txu48a;

  assign zti98n829owa2p = ap0oygari76txu48a ? pn1rzse3t9e6g_et37gv : isqt1ng7lccfet8bj5hym5c;

  assign v2tse065uysfbl8f4z8hlpkg5o68 = zkojor8433oflab2kpvtzi1z9;
  assign kwczwxezdeidftn2_p2fpzik3gt = nx6i4o0_cbqmlan1ylpodj9y;
  assign o58xzacx8hg_9zcqk21v9m0rqqsap22_ = tgfv2w2s7qhwkl0pdpf_79v4e;
  assign q0xni3yf49f2fj7ymo_nvdurqx1okyv = qfjl6250hpfb57pxl0t53q6fd;

  assign xmf6kblqlhyjpa44uj3tn_7hs9g = zkojor8433oflab2kpvtzi1z9;
  assign td_dxcgpaod7g2fvddly_mg4rjh2vgbk = nx6i4o0_cbqmlan1ylpodj9y;
  assign l1mayxu6go0ni6a1uu2tn40qyps5l_ = tgfv2w2s7qhwkl0pdpf_79v4e;
  assign qdf9k5s3p4c0d8jxgmxlyi478ade = qfjl6250hpfb57pxl0t53q6fd;

  assign ije4h78_umvknjj6az4_5qf92e3iydh = ye256knohacnaakiw2nqck6;
  assign sro97_d1rgt1fmqi2b_fitscvexczye2 = hyxeikuobvxjumz2hibay;
  assign lwmr8fyosc4w78ftaznb17d0wep6 = ye256knohacnaakiw2nqck6;
  assign g_lbo1t8r4bx4olr034dfi8fhfw1m6i = hyxeikuobvxjumz2hibay;
  
   



  assign jkq984ky8fozrzq = a5s2gi2_h7rplzkx1 | on12sjnlw0b975rtxnj;
  assign g3_8p4g7w5grnl62xy = bekul5xbo28zkmc90zy ? gn916lc8_fzkp3rcqpob : m91uirvkay9adfjui930dyv4;
  assign a_i3c4odzkmjpufk2pffcu = vqwqaofc8sz_yjccd & (~bekul5xbo28zkmc90zy);
  assign nepu6mf61h2b2uewptpauek6v = vqwqaofc8sz_yjccd & bekul5xbo28zkmc90zy;


  assign agnsw48g8fdikd     = cgnsvvj7srbljqst;
  assign x25ltyb13sb2td2     = cgnsvvj7srbljqst;
 
  assign j2kcz1faqhvh1ler6j   = bekul5xbo28zkmc90zy ? idcribpugamfq_39t   : rbkhb89tyu_ucjpo    ;   
  assign a6gdkt5h77dh0mcj8t4gq = bekul5xbo28zkmc90zy ? nfuf_njr73sjp5jr12d7gc : sqvgnqdrkexeg2lziofadt  ;
  assign wixbtbeqlhzelg4t   = bekul5xbo28zkmc90zy ? hgm8yvqudk9e2ne6   : bwtzw5pqhc62g9v9w    ;
  assign uh_ekyw7cw8c3d3xj1  = bekul5xbo28zkmc90zy ? ivt9rgs2qqjzyrq5zt4isy  : nwbvll63g8yq6vbpxok   ;        
                          
  assign uf44audysjgtvdnua67   = bekul5xbo28zkmc90zy ? u6di3j5ypwgwjvnmcbsqh   : e4ui35hoxqcwkgfaol    ;
  assign qtcasxm90cy0bwaqaxz = bekul5xbo28zkmc90zy ? i7vlo92n37lvcod6oj : f1uy000fu6355gukzxt9r4y  ;
  assign y38seii6ja77q2jy08   = bekul5xbo28zkmc90zy ? ulp1cmdd07o0vc3p_65wi   : avudrqvyzx1dringrt4rs    ;
  assign f42g8ulc2y43ntmai5  = bekul5xbo28zkmc90zy ? f9_zg3c33q9sbq6d82u  : hz5leo9sklh2v25_50   ;        
                           
                        
  assign rgf8pa4kn20jusruz   = bekul5xbo28zkmc90zy ? mgc5k45s6iun0h64mg94n   : ofg0te04_oeiba586    ;
  assign wjwjffxr_4lulivwz = bekul5xbo28zkmc90zy ? kuhd9_39ag_1mza9vf7x : dm0uaanzcp_7hojw2_h  ;
  assign z6udkjbx164gh9yo1o  = bekul5xbo28zkmc90zy ? dbp3mo7p_zh0242q9  : yddyulfbyf7p2wvl6dyk   ;
  assign frkunk72hlttw0ar0np  = bekul5xbo28zkmc90zy ? enbd230u3ab6jrd2gt  : j233e_ya9xhnxg7flb9d3   ;        
                       
  assign r2tvaf8px0p9vlw4we   = bekul5xbo28zkmc90zy ? nwvjy589molbkspazci   : mq3a_g7zrfyfdil1    ;
  assign srfn4smswwo6hbyaa = bekul5xbo28zkmc90zy ? hkv3jt_7_o_8sk0aait_0kp : f9ekxi98w3bnnfm3t1vyt1  ;
  assign a_u2kfmgv2ho357c  = bekul5xbo28zkmc90zy ? dzca_d1t69gei8viv2q  : k1vhaduoq3xy5cx6jr0   ;
  assign svj88sv2u56fepzmg  = bekul5xbo28zkmc90zy ? w7paq1qa9rrtadyr3v3cx  : hwo9njh5b4299teslcl   ;        
                         
  assign rzf167thmprvps0tm62i   = bekul5xbo28zkmc90zy ? ky3t5ldjtr_g__hnxr58s   : shxdziymfk57c49e0    ;
  assign lv7fu0hif2n2zhmgtcc = bekul5xbo28zkmc90zy ? l20gjym8j9s2t31_nhs8iuh : s_fatq1jfpqkf7q9d40n  ;
  assign oj5t3f0lq1n9ae82x  = bekul5xbo28zkmc90zy ? r3kh4eweep0kg7fak6rx6f  : ruix76vs69a8gynr7yydnp   ;
  assign hat38salswlktk821  = bekul5xbo28zkmc90zy ? vwj6zdjeua22z66vj  : y0s6zoimyz170437bgkne   ;        
                        
  assign caxkrdjq0tjnnne9   = bekul5xbo28zkmc90zy ? tbykhfjbcc3ure59   : nsyif4pw3tzuggdakg2    ;
  assign qpuk8ry0w9_r7ur4gcnx = bekul5xbo28zkmc90zy ? v0oz07osad44us4h0pyd : e4zsuzpz_sgcgql5k19iv  ;
  assign v8jl1eh8o0n5g765  = bekul5xbo28zkmc90zy ? xtiqejiid_qbh90nn_jv  : fvzgpoei5_ffhtrv6r   ;
  assign c0xnu9p8he2hw10h  = bekul5xbo28zkmc90zy ? dzoe86_fm7z7_c7_4_zn  : cnqt629_5e9xaypczfdt   ;  



  assign ktkt_7t0wo1gkg8gormhm = rjy1ysvx9590bpklijsn0ucgaga;
  assign s9lcmqjp282zoimy_nw6kv2u = pkm6vgcr8iz_el5103gzwdew0hki;

  assign o3ydhguk119jyhp47x106ib = opa_i9g_7se8iof9su_mxicjyu;
  assign b4687t39adr64eo0i4lf5md = n1bimos0aw0citrgtz3yco;

  assign hv39pppvbmeqy8b6        = opa_i9g_7se8iof9su_mxicjyu ? no360dfthc_r812ltoqdhrz        : piosx1_uvpor01vn8ll66_yhit        ;
  assign t6l88yqbe4wokkhiso9t       = opa_i9g_7se8iof9su_mxicjyu ? enqm3v278hn097pt6_04p9n       : fsgnhdgr565rvtm7jewinuufhjm       ;
  assign hyec__ebnw8lbcssd81       = opa_i9g_7se8iof9su_mxicjyu ? hs3xn0evnbpy575ea7p5p3qto53       : ilmemra32cftf81jy7tb1tn       ;
  assign vs2610q9_on1r996p      = opa_i9g_7se8iof9su_mxicjyu ? sycglehz7v8eijxjqe7ufoxp4j1y      : p8rx6454dkq9mcu0knbdrp4      ;
  assign coy3buxdw6yq3duh21azuwflk = opa_i9g_7se8iof9su_mxicjyu ? pihkjnbghw4bk8y2477x7k82o93ug : oy5tnom44u2vm3zpklpy9_xsje_dh ;
  assign r_8h5lxb39ug57zli04e_o      = opa_i9g_7se8iof9su_mxicjyu ? crriagr_kegsjfrtly_v8yw9      : enjo_thzs5fjl2yaorgzrh85sivo      ;
  assign pv7q0ikpayogkay57rgyr      = opa_i9g_7se8iof9su_mxicjyu ? p5u44x4jrltstcsbmk8kg5hnq0      : eg3xuv8r03e6j0msnfyr8i2b      ;
  assign ou74jmm5p6th0y0kcdwpqv2ey = opa_i9g_7se8iof9su_mxicjyu ? gg0tr7jpfos4ct46rnx8kikun5t6ee : ydi3gh_3ks81b74d8g9vgn081jicdv8 ;
  assign adwzzx09c_s_x1seh      = opa_i9g_7se8iof9su_mxicjyu ? vfxj481iib57qmfew_ggqin2rqaa      : ce_6thxzv8n4n8xdhg9y9ftl      ;

  assign ve1mua6_hp7e4a8tf03lfitualb     = dsq8f3rhmb7yc876v8  ;
  assign tl82sx3puyxv5f6eoxlnfunqhe8    = zp0aylmm0k4yw4w561bgzh ;
  assign m7fr__lszd5b56qf13pbarusep    = enu_vumk17eoj1fma5ilz0 ;
  assign kc_oc1b1x6hj408h8pkuuwr09qnr     = dsq8f3rhmb7yc876v8  ;
  assign xg81tsg3z29z7lie1domdmt86crlg    = zp0aylmm0k4yw4w561bgzh ;
  assign zjp7e4i7qt_0abds5ihh_dnqk    = enu_vumk17eoj1fma5ilz0 ;

endmodule






















module ktpcxlh_26k125r(

  input  rm1dxjejhq7dh3q5m,
  input sxvvsxtbhyvt,

  input [8*32-1:0] pcr4upio7_tx37, 
  input [8*1-1:0] uzklqlncpqqm1rav,
  input [8*1-1:0] ortueunvnkx_l5m_j,
  input [8*1-1:0] hwuhtb7ucto_utk56,
  input [8*2-1:0] i1env2kmns7qvvuuc,
  input [8*1-1:0] g3s3vpafvy3i,


  input  c4ughu0qm5sfai,

  input  tia1md5dyh6kj4,

  input  indfp6mwqdqamez0mex,
  
  output                          p7ah58va5_2njbtv, 
  output [64-1:0]         u981qrwkgi5h0e72b__gg19w,  
  output                          p0i2i3v3j1tclelx51,  


  input  j8cjhcuf0m6xjvemdaz,
  output s_eowfyzlvx7gjv542upo,
  input  q7ru87fmzxczveihcxcwh,
  input  umc_2tn6um_9xaiy7_ksg0w,
  input  uiyh4da4134sjv7gnmc,

  output r5hpbriny8m67sv9e_ylgo1,
  output dyl5g2vgrvy4mb3,

  
  
  
  input                                    ysnexkrvlg2s55ajc5g69tm,           
  input  [74-1:0]       p7832rg37bbm7_ssxunhcj7,          
  output                                   t1xtkdoie_8djygqlt1br56pwt,         
  output                                   w33zvryieg8hhgy58581ny437h9,           
  output                                   lv96t6re1w44borcb7do83ndua3vjy,      






  input                           th06du2c8e2_b7k,
  output                          irjoi8wvo25u209f_5,

  input  [32-1:0]    zvk11dhgg2s67mkq, 
  input                           fbzs0o4ysyuzeg_qdj, 
  input                           me1n4pvwxa7n3u8l05, 
  input                           qaidts35dk5jcji0n, 
  input                           uo0ftugxv_yuoh, 
  input                           dcj485cah5, 
  input                           zxe59xihintdqfy9d, 
  input  [64-1:0]       u4r4b_6kp09q767q,
  input  [8-1:0]       lhibcc3xwm6cy,
  input                           hc2ava5u3xa_bw0,     
  input                           erz5xg5fnrald,     
  input  [1:0]                    r19ik0uppwcr,


  output                          klkflmsyyf5w7ar,
  input                           wy36iirxspfw56864,
  output                          lkjqs6kiuyj,
  output                          u245it8jnyhc3eqcy0,
  output [64-1:0]         h7f6k_ims_9p3, 



  output                          cv0k9k_ijjnnylw1s7b_0d,

  output                          swpk4h0gei3t_34xogbqncbo4,
  input                           u9qmfl3rwx0dhr92z875vx7q,
  output  [32-1:0]   unu_x_i6jmr33nz0yitzk, 
  output                          bei3qhdtd0euq2emblogsu_x, 
  output  [64-1:0]        bf0_ynb648lqi7s93eieo0ln,
  output  [8-1:0]     wf8o7p9_qfthhoxs747wyeuwkky,
  output  [2:0]                   ygro7xue7x7rtdafkj3o4q4,
  output  [1:0]                   drrly3q0ocg8d4pwh3m9o77,
  output                          g654a6a9cesbee7xs6_uu9lu5,
  output                          x7fex0jf9da6a5v1c28upl72t,
  output  [1:0]                   ege0_1ufqm8i68zo4il6cwe46d,
  output                          ngyxf4n1cpcgks_s2zmgfb260, 
  output                          c7m50uaw8lmp_iv4ci38q2, 
  output                          m04a1mtbabwezldp1crh4rg6z, 
  output                          hwjq1ubtaei44lpk609fm2hb8, 
  output                          e28p_fu1k484ncul0p85ko, 

  output                          a0_d_zdz9h9fgk46e8arf,

  output                          twr9y24wxhs3qj2z9f2hzpaig6,
  input                           w8b46r9cof57xvd5zo1u4zh8,
  output  [32-1:0]   wn1l4cmih7rwce1rb7wk3f9wy, 
  output                          cgnzbuo_1yz6v42seb25duv, 
  output  [64-1:0]        zopev7f487spn9mwvuowqo,
  output  [8-1:0]     p32jk0lb8g31kqlpvmllo75qim,
  output  [2:0]                   g973rcaou05i456suvk_89dm,
  output  [1:0]                   wflv6rhfdwyxttak111v1l,
  output                          ggsmt4nzx8pwlowehinqvk60f,
  output                          xu8494ii8ectqb91224uuer,
  output  [1:0]                   r6rk128ijo839ougen9stbe,
  output                          xo6ciibewn8p8xey97jcsqi5, 
  output                          evz1w_girwszyfnlcg4mwvtjo, 
  output                          ju5f9fb1erjep_bv8gpfn6, 
  output                          hadi1_f3quoaotjv5758x8kksot2, 
  output                          bdi4gjlb0po4ejcztowoqil7, 



  input                           bvg_3t_ujbpur7b_h7f63jse,
  output                          m5l6wu3uz_jfqasz8e3tsvrm,
  input                           g9so28ythfl0q7xnk66p1  ,
  input                           e66wluxk71p2ldu3a1qk994bq,
  input [64-1:0]          ig2roj0y08x8_ntp3knz9rd, 

  input                           m7tq_t57mr5bovbb9ghffl4k,
  output                          gpcgdcri3e6_fxrw8wwtysoqqr,
  input                           a6s4kxg1ibr6mntc85jik  ,
  input                           hizzalmpwr8cqkxqi80wvbt65x,

  
  
  output                          mum8f1rtatle7p_55y84,  
  output [6-1:0]  pn5bpwlp5ijfako9m5ao,
  output                          g3s0qe2adsxsx8e6z ,
  output [24-1:0]  a1rl4lmhqp8ydyk07kqkn,          
  input  [24-1:0]  apnns9jlj7y3y5bg8ynz,
   
  output                          pmz7e4mgvbnmimqp0nghk,  
  output [6-1:0]  j61algpxjoycxbswhgsuf, 
  output                          omq1ehm8hp4q9jgp5n5vn ,
  output [24-1:0]  fbv1q6sraswzp91zcn,          
  input  [24-1:0]  jv8kv41vzuir6an4iod,


  
  
  output                          qgl4363n31jx6xjyo05zkn,  
  output [8-1:0] zec78nyllxlfwmpsgncluudf, 
  output [4-1:0] dwvnjl0vxqkgd8t6dtvg5z,
  output [32-1:0] gngmcj5c1jd85csel9ntru,          
  input  [32-1:0] tkt93y5lfluzkia5plvksp,
                                                
  output                          km7co8hqm563od8ga_03_g,  
  output [8-1:0] j4mas6g26o63wvnsdquh8c4p, 
  output [4-1:0] nniah5mh0cunkhyln9,
  output [32-1:0] rcy_v3911lf33nza5j,          
  input  [32-1:0] g4nfgu53_rgc0632w8z97,
                                                
  output                          xzgkclcxsgfuseg87,  
  output [8-1:0] djwlah5bo0r6myit6cal0t, 
  output [4-1:0] qu_ju3lv6nvkdbo8h11uf,
  output [32-1:0] dydwz9i6k80alqfarffop,          
  input  [32-1:0] ql1c7hzoj9kf__7r97krm,
                                                
  output                          kp2j8kv1p1cjcg0lerwm,  
  output [8-1:0] v4a7g1wh3ivw0esp7dye0oiz, 
  output [4-1:0] x9zuk21gpaj58uszvm5,
  output [32-1:0] n_h5oz0c5bo5rpevwjcu8,          
  input  [32-1:0] ryid4_99ns1jc83at_88x,

  input  gf33atgy,
  input  ru_wi
  );


  wire                               hv39pppvbmeqy8b6;
  wire [32-1:0]           t6l88yqbe4wokkhiso9t;
  wire                               hyec__ebnw8lbcssd81;
  wire                               vs2610q9_on1r996p;
  wire                               coy3buxdw6yq3duh21azuwflk;
  wire                               r_8h5lxb39ug57zli04e_o;
  wire                               pv7q0ikpayogkay57rgyr;
  wire                               dsq8f3rhmb7yc876v8;
  wire                               enu_vumk17eoj1fma5ilz0;

  wire                               ou74jmm5p6th0y0kcdwpqv2ey;
  wire                               adwzzx09c_s_x1seh;
  wire                               zp0aylmm0k4yw4w561bgzh;


  localparam r4bbs1l72_cd3t_ = (6 + 1);

  wire yb5ru177dkq2qb; 
  wire c_0qdn252ww1o9nhj4m; 
  wire x0pxzzrure0tp8zh3; 
  wire nvlcc2cq4xv0339t;
  wire j55vt_3172gxi8el;
  wire t8yi927p43l4;
  wire bda77mp8zde61a_;
  wire re8ax_cpd2o8l;


  wire nmqf8r7zm2wfw8pz;
  wire o9jixjnak_33vfbl;


  assign r5hpbriny8m67sv9e_ylgo1 = 
                       | j55vt_3172gxi8el   
                       | (~bda77mp8zde61a_)
                       ;


  wire s_fxmgzl8pdoycnrftl7z7wz = 
                         yb5ru177dkq2qb 
                       | c_0qdn252ww1o9nhj4m 
                       | x0pxzzrure0tp8zh3 
                       | nvlcc2cq4xv0339t
                       | j55vt_3172gxi8el
                       | o9jixjnak_33vfbl
                       | (~bda77mp8zde61a_)
                       ;

  wire b9b7j_s1j6pzebjxovfv6t = 
                         s_fxmgzl8pdoycnrftl7z7wz 
                       | t8yi927p43l4
                       | th06du2c8e2_b7k
                       ;

  assign dyl5g2vgrvy4mb3 = b9b7j_s1j6pzebjxovfv6t | j8cjhcuf0m6xjvemdaz
                       | re8ax_cpd2o8l
                       | nmqf8r7zm2wfw8pz
                       ;



  wire                        qe0x130i0z960a1ld7jru7ma         = p7832rg37bbm7_ssxunhcj7[0    ];
  wire                        z2w73ziehrytb1m0t4jo_jr0ici        = p7832rg37bbm7_ssxunhcj7[1   ];
  wire                        qmpmjqpq_d69kzu6u9bxjr74w1y        = p7832rg37bbm7_ssxunhcj7[2  ];
  wire                        e09r0m8969cj0sl6_iwpy513ad9kih       = p7832rg37bbm7_ssxunhcj7[3];
  wire                        oithmqsqi28np858lo1dztmf         = p7832rg37bbm7_ssxunhcj7[4    ];
  wire                        axgfwdkn0nyose7m3bwgcx92jc5gl61      = p7832rg37bbm7_ssxunhcj7[5 ];
  wire                        dyw1ymrkp8_lbpgb36w25d8fef1      = p7832rg37bbm7_ssxunhcj7[6 ];
  wire                        gq9tfy8ozjrgv8isn05omqqolwzip      = p7832rg37bbm7_ssxunhcj7[7 ];
  wire                        pvt527iyu2jjdtrzg1dhd0zi084q0nmww = p7832rg37bbm7_ssxunhcj7[8 ];
  wire                        n3vgs5xww30vllhavnnqse8w0t8mrph = p7832rg37bbm7_ssxunhcj7[9 ];
  wire  [64-1:0] jkptde77bwbsv8niyj78xrgj8vz6mus1  = p7832rg37bbm7_ssxunhcj7[74-1:10  ];
  wire  [32-1:0] erg8nrhaecoc2m5idim8fol1zo25m         = jkptde77bwbsv8niyj78xrgj8vz6mus1[32-1:0];

  assign re8ax_cpd2o8l = ysnexkrvlg2s55ajc5g69tm;



  
  
  
  
  
  

  wire niejxpmibm8_c3z9;
  wire d8fgkbjcpmd8_4r;

  wire jo2m0mwneyhm = (t8yi927p43l4 & niejxpmibm8_c3z9);
  wire u3gm9gusc9log5m42rc = (nvlcc2cq4xv0339t & d8fgkbjcpmd8_4r);


  wire [32-1:0]    a7h_7269eov; 
  wire                          z7yrukhpu2yv7; 
  wire                          haj3ixozrokecb; 
  wire                          b1ojpuh8kzteazg; 
  wire                          al2dpsmo5cx28; 
  wire                          ulo4ekmq8z3kurrev0okj; 
  wire                          kqbdvrqc2ega5n0a; 
  wire                          go95at_xv3zz734; 
  wire                          w1uq15jgugrn3; 
  wire                          n15yjlq97s5vf9; 
  wire [64-1:0]       yqy4lcoychj91n;
  wire [8-1:0]       qnwoumw9i3v36;
  wire                          a5atqg2vaqg92ov;     
  wire                          ahxhj9pllg;     
  wire [1:0]                    y9f19nzrdlvvh;
  wire                          wzpsauw3j_6xyp0;     


  wire [32-1:0]    dm_t8xh6s80cssm; 
  wire                          lwq70xytakc30w; 
  wire                          d2lwzgwj549p; 
  wire                          vuqz2ck550pkhan; 
  wire                          gcio7gsqtef4lbth; 
  wire                          rrgpiz3c94ildst7z_; 
  wire                          v6m8pnzviydxj77_a_f6h; 
  wire                          dqpjx6e7kt6x2csta; 
  wire                          a7hxr7wh300y3; 
  wire                          io1dzzuksv6fh6w; 
  wire [64-1:0]       ctciq9lwt094amf;
  wire [8-1:0]       c04en6bt2lvr5;
  wire                          q8aypq1prdr34cq;     
  wire                          csirbohj0gm_cfs;     
  wire [1:0]                    gstkdmb4wbsp8xhi;
  wire                          rnj3s81yxus08gthgj;     

  wire [32-1:0]    pq05yc_ea9cb; 
  wire                          bqbd1vx7u6p; 
  wire                          io1o8wz_hhx_efhn; 
  wire                          ar75eg689jsahd; 
  wire                          lv2obxi3r4ob; 
  wire                          l3i_yp_t5k_ghmdbmvrk4; 
  wire                          ntwmchaa8jnutooi3_; 
  wire                          y2yeehopezll49cmf; 
  wire                          g5dm3flv9; 
  wire                          jxbtey15c3kkb7; 
  wire [64-1:0]       rxps0kbgar3hf;
  wire [8-1:0]       kogy6rrqymszp;
  wire                          hqchs835s6qbo2wr;     
  wire                          kfjijv_31s3;     
  wire [1:0]                    g6qm6ye0l65m;
  wire                          yqc55f6txw_pmexi;     

  
  wire [32-1:0]    fwgc_k58kjyp_va; 
  wire                          etwu6izome4p5cwa0gn; 
  wire                          xa3kdso6mkaf3rs_51f; 
  wire                          w8oyx6w2m20wkhtzop; 
  wire                          jab9p1mpwm16j6wmz3hs; 
  wire                          u3fovt7dw2e5zglu0b_3uen0m; 
  wire                          f4c6lj0xc31c5ibnegpv6ymsi_; 
  wire                          epi1zu1tfkun1al0l9; 
  wire                          n29ai3bkicr4tgyzgk; 
  wire                          hh6d0ibqo915gqaoole; 
  wire [64-1:0]       herh0nxfburswr1cgvh;
  wire [8-1:0]       l1ic10plktexvczv;
  wire                          g7m6bw52bw7jvu414;     
  wire                          gaqzi18ded72q1bbz4p;     
  wire [1:0]                    xkopv4_km4ey9cihevo2;
  wire                          v_9kfy4x1fk3adyoz6x2;     

  wire [32-1:0]    pte_y5zn1kqfnzxo5izs; 
  wire                          ne3qv25fuqotk2dk5; 
  wire                          ycqmiyj7jekquq0pxuy1uk; 
  wire                          dryvl0kbql72b720rm; 
  wire                          fsqkwjz0sanwked5rfthn; 
  wire                          m5uxjf11e0v1munmybb1n3fv; 
  wire                          eschp5gtzyhx77wg6jhl4z9ny; 
  wire                          wo477hsguadhf4cwa9bbl; 
  wire                          fsfq1s74k43eb5l; 
  wire                          yajgwlnlp6hvh354akt3lm; 
  wire [64-1:0]       gec3f9o0vmsnfdwup7xem;
  wire [8-1:0]       fy5zq5a7ou_6sownckex;
  wire                          xopz5es01zuocuhfzv;     
  wire                          j9ngo4gtwitbihmi5djct;     
  wire [1:0]                    hmaam0gy6lvgx07vlp6yo7;
  wire                          foma9juy1lv_7626wum__ceu;     

  localparam f16zrowg1s1f5 = (32+9+64+8+5); 

  wire [f16zrowg1s1f5-1:0] ez0jkdg20o7_ib;
  wire [f16zrowg1s1f5-1:0] se0zyj4n4upz;
  wire [f16zrowg1s1f5-1:0] cdqzid8vpi25lg6fx;
  wire [f16zrowg1s1f5-1:0] k8qtf1i196m8bfpmqi;

  assign ez0jkdg20o7_ib = {
                                           zvk11dhgg2s67mkq  
                                         , 1'b0
                                         , fbzs0o4ysyuzeg_qdj  
                                         , me1n4pvwxa7n3u8l05  
                                         , qaidts35dk5jcji0n 
                                         , 1'b0
                                         , 1'b0
                                         , uo0ftugxv_yuoh  
                                         , (dcj485cah5 | (~tia1md5dyh6kj4)) 
                                         , zxe59xihintdqfy9d  
                                         , u4r4b_6kp09q767q 
                                         , lhibcc3xwm6cy 
                                         , hc2ava5u3xa_bw0      
                                         , erz5xg5fnrald      
                                         , r19ik0uppwcr
                                         , 1'b0
                     };


  assign {
                                           a7h_7269eov  
                                         , z7yrukhpu2yv7
                                         , haj3ixozrokecb  
                                         , b1ojpuh8kzteazg  
                                         , al2dpsmo5cx28  
                                         , ulo4ekmq8z3kurrev0okj  
                                         , kqbdvrqc2ega5n0a  
                                         , go95at_xv3zz734  
                                         , w1uq15jgugrn3  
                                         , n15yjlq97s5vf9  
                                         , yqy4lcoychj91n 
                                         , qnwoumw9i3v36 
                                         , a5atqg2vaqg92ov      
                                         , ahxhj9pllg      
                                         , y9f19nzrdlvvh
                                         , wzpsauw3j_6xyp0
                                                             } = se0zyj4n4upz;



  wire [f16zrowg1s1f5-1:0] tv1vy00negaq6kq;
  assign {
                                           dm_t8xh6s80cssm  
                                         , lwq70xytakc30w  
                                         , d2lwzgwj549p  
                                         , vuqz2ck550pkhan  
                                         , gcio7gsqtef4lbth  
                                         , rrgpiz3c94ildst7z_  
                                         , v6m8pnzviydxj77_a_f6h  
                                         , dqpjx6e7kt6x2csta  
                                         , a7hxr7wh300y3  
                                         , io1dzzuksv6fh6w  
                                         , ctciq9lwt094amf 
                                         , c04en6bt2lvr5 
                                         , q8aypq1prdr34cq      
                                         , csirbohj0gm_cfs      
                                         , gstkdmb4wbsp8xhi 
                                         , rnj3s81yxus08gthgj 
                                         } = tv1vy00negaq6kq;

  wire [f16zrowg1s1f5-1:0] gs05ko46ogh5;
  wire [f16zrowg1s1f5-1:0] ts27sjuboaf8qsmg;

  assign {
                                           pq05yc_ea9cb  
                                         , bqbd1vx7u6p  
                                         , io1o8wz_hhx_efhn  
                                         , ar75eg689jsahd  
                                         , lv2obxi3r4ob  
                                         , l3i_yp_t5k_ghmdbmvrk4  
                                         , ntwmchaa8jnutooi3_  
                                         , y2yeehopezll49cmf  
                                         , g5dm3flv9  
                                         , jxbtey15c3kkb7  
                                         , rxps0kbgar3hf 
                                         , kogy6rrqymszp 
                                         , hqchs835s6qbo2wr      
                                         , kfjijv_31s3      
                                         , g6qm6ye0l65m 
                                         , yqc55f6txw_pmexi 
                                         } = gs05ko46ogh5;

  wire [32-1:0] fzebl49irts00yi4k6c; 

  assign ts27sjuboaf8qsmg = {
                                           fzebl49irts00yi4k6c  
                                         , lwq70xytakc30w  
                                         , d2lwzgwj549p  
                                         , vuqz2ck550pkhan  
                                         , gcio7gsqtef4lbth  
                                         , rrgpiz3c94ildst7z_  
                                         , v6m8pnzviydxj77_a_f6h  
                                         , dqpjx6e7kt6x2csta  
                                         , a7hxr7wh300y3  
                                         , io1dzzuksv6fh6w  
                                         , ctciq9lwt094amf 
                                         , c04en6bt2lvr5 
                                         , q8aypq1prdr34cq      
                                         , csirbohj0gm_cfs      
                                         , gstkdmb4wbsp8xhi 
                                         , rnj3s81yxus08gthgj 
                                         };


  wire [f16zrowg1s1f5-1:0] tvypfoh27qvczot = {f16zrowg1s1f5{1'b0}};
  wire [f16zrowg1s1f5-1:0] ky8zw277b8fa1dq1zk;

  assign {
                                           fwgc_k58kjyp_va  
                                         , etwu6izome4p5cwa0gn  
                                         , xa3kdso6mkaf3rs_51f  
                                         , w8oyx6w2m20wkhtzop  
                                         , jab9p1mpwm16j6wmz3hs  
                                         , u3fovt7dw2e5zglu0b_3uen0m  
                                         , f4c6lj0xc31c5ibnegpv6ymsi_  
                                         , epi1zu1tfkun1al0l9  
                                         , n29ai3bkicr4tgyzgk  
                                         , hh6d0ibqo915gqaoole  
                                         , herh0nxfburswr1cgvh 
                                         , l1ic10plktexvczv 
                                         , g7m6bw52bw7jvu414      
                                         , gaqzi18ded72q1bbz4p      
                                         , xkopv4_km4ey9cihevo2
                                         , v_9kfy4x1fk3adyoz6x2
                                         } = ky8zw277b8fa1dq1zk;


  assign cdqzid8vpi25lg6fx = {
                                           pte_y5zn1kqfnzxo5izs  
                                         , ne3qv25fuqotk2dk5  
                                         , ycqmiyj7jekquq0pxuy1uk  
                                         , dryvl0kbql72b720rm  
                                         , fsqkwjz0sanwked5rfthn  
                                         , m5uxjf11e0v1munmybb1n3fv  
                                         , eschp5gtzyhx77wg6jhl4z9ny  
                                         , wo477hsguadhf4cwa9bbl  
                                         , fsfq1s74k43eb5l  
                                         , yajgwlnlp6hvh354akt3lm  
                                         , gec3f9o0vmsnfdwup7xem 
                                         , fy5zq5a7ou_6sownckex 
                                         , xopz5es01zuocuhfzv      
                                         , j9ngo4gtwitbihmi5djct      
                                         , hmaam0gy6lvgx07vlp6yo7
                                         , foma9juy1lv_7626wum__ceu
                     };



  ux607_gnrl_bypbuf # (
   .DP(1),
   .DW(f16zrowg1s1f5)
  ) jesp83ag2itrtu0u991z (
   .i_vld(th06du2c8e2_b7k),
   .i_rdy(irjoi8wvo25u209f_5), 
   .i_dat(ez0jkdg20o7_ib ),
   .o_vld(t8yi927p43l4), 
   .o_rdy(niejxpmibm8_c3z9), 
   .o_dat(se0zyj4n4upz ),
 
   .clk  (gf33atgy  ),
   .rst_n(ru_wi)  
  );







  
  
  
  
  wire  bpmlbcph7uz4fmydd;
  wire brfek3hm0m1h_0qdx;
  wire t1cqzavxcqpcddy3yhtk;
  wire pn0blb6qozvruaiaccluecd;

  wire  dsrz57a4u1pediag;
  wire c5luf4ekdp8uxjd6phdb;
  wire cik9g8nrdjspswqucoa9;
  wire w3o65s8zjg4wgjw69l7iz58u;

  wire q6dwr6kors49;

  wire vc0fhfx87dxbgty02yd;
  wire stdkgs3cetkrgnprgzkr;
  wire ytaw26fvd4q2bkrmzdzc20exc7nofso;

  wire [2-1:0] qb0k_89eoa;
  
    
  wire jgd_t54t3z41vhe = jo2m0mwneyhm | stdkgs3cetkrgnprgzkr;
  
    
  wire ypahzv06s1rdg2 = (q6dwr6kors49 & (~vc0fhfx87dxbgty02yd)) | ytaw26fvd4q2bkrmzdzc20exc7nofso;

  wire jflxgnf39_p3z1e6 = jgd_t54t3z41vhe ^ ypahzv06s1rdg2;

  wire [2-1:0] bj7ex6wl29354zmz = 
                                   jgd_t54t3z41vhe ? (qb0k_89eoa + {{2-1{1'b0}},1'b1})
                                               : (qb0k_89eoa - {{2-1{1'b0}},1'b1})
                                               ;
  
  ux607_gnrl_dfflr #(2) i4vlss_y0l22e (jflxgnf39_p3z1e6, bj7ex6wl29354zmz, qb0k_89eoa, gf33atgy, ru_wi);
  
  wire dl1e0uq8c1swic = (qb0k_89eoa == 3);

  
  
  
  
  
  wire padw0r9xyxkm36fh = yb5ru177dkq2qb 
                       | nvlcc2cq4xv0339t
                       
                       | o9jixjnak_33vfbl
                       | dl1e0uq8c1swic;

  wire oxqqtcjokpeaecyynig; 
  wire pleylcyovtj6ttr34;  

  wire f56j5y58ce35hwpqbnu16;
  wire nk4gkqhhy_a4hc5n4kin;

  assign oxqqtcjokpeaecyynig = (~padw0r9xyxkm36fh) & t8yi927p43l4; 
  assign niejxpmibm8_c3z9     = (~padw0r9xyxkm36fh) & pleylcyovtj6ttr34;  

  
  
  wire dr91idf72q6degdldki7 = f56j5y58ce35hwpqbnu16;
  wire lb7s03sx7nyfkkndx_y = bpmlbcph7uz4fmydd ? nk4gkqhhy_a4hc5n4kin : 1'b1;

  wire x42fyhas4g32apt7tjeq8 = 1'b1;
  wire hptdr4euu3t87qoy4btzp8 = bpmlbcph7uz4fmydd ? 1'b1 : 1'b0;


  wire p0brv6fqgdvccaui21k8 = oxqqtcjokpeaecyynig & x42fyhas4g32apt7tjeq8 
                         & lb7s03sx7nyfkkndx_y
                         ;

  wire j30h3wzip_eqif46u34tw4 = oxqqtcjokpeaecyynig & hptdr4euu3t87qoy4btzp8
                         & dr91idf72q6degdldki7
                         ;

  assign pleylcyovtj6ttr34 =
                         & dr91idf72q6degdldki7
                         & lb7s03sx7nyfkkndx_y
                         ;

  wire y85uyrjj282xf9p3it0u2wvmixet;
  wire ijsk41ad4tvq4zse7kouzpbxcnck2;
  
  
  
  wire g_wql4uu07mqqw8qgtprsk8xoaul = y85uyrjj282xf9p3it0u2wvmixet;
  wire uzy1lty2609v_xavjbkoacvvkv5 = pn0blb6qozvruaiaccluecd ? ijsk41ad4tvq4zse7kouzpbxcnck2 : 1'b1;

  wire m5xxp4vmnpskm89gjfufm23 = 1'b1;
  wire q966g40h505gzbfbtj9sp392n = pn0blb6qozvruaiaccluecd ? 1'b1 : 1'b0;

  wire hcjwu1jmlbr4k4wahdf0ju;


  wire dq71bajnhqrbc7pjo3ilkqpu00atil = hcjwu1jmlbr4k4wahdf0ju & m5xxp4vmnpskm89gjfufm23 
                         & uzy1lty2609v_xavjbkoacvvkv5
                         ;

  wire jo20b3jp2h86mzvqeae5j3xsu3g3 = hcjwu1jmlbr4k4wahdf0ju & q966g40h505gzbfbtj9sp392n
                         & g_wql4uu07mqqw8qgtprsk8xoaul
                         ;

  wire k71jdwvt1q_yy5a7kzwp8cz =
                         & g_wql4uu07mqqw8qgtprsk8xoaul
                         & uzy1lty2609v_xavjbkoacvvkv5
                         ;

  
  wire f1xe_xx4j29e7277py1p2k9uh;
  wire ra61k0r5_z16sciiz8un534o6w;
  wire ujuhwx1rtmvxjxxpbmlhcttboa3kd;
  
  
  wire zylypzxl2r1asy4_sbdielf_2;
  wire eqce_y4zxdhu7zaz6s2fk7vec = (~zylypzxl2r1asy4_sbdielf_2) ? ra61k0r5_z16sciiz8un534o6w : 1'b1;  
  wire m7frhh6dekyuotcrluw9m36kvn4 = ujuhwx1rtmvxjxxpbmlhcttboa3kd;

  wire v2xjuhisvq_5yd8vq6__k0ijc = (~zylypzxl2r1asy4_sbdielf_2) ? 1'b1 : 1'b0;  
  wire vfjafvqeepaxiqz2w76pl8ds6z = 1'b1;

  wire rguv86jfrc_9hefk7y2yvxn6og4d1 = f1xe_xx4j29e7277py1p2k9uh & v2xjuhisvq_5yd8vq6__k0ijc
                         & m7frhh6dekyuotcrluw9m36kvn4
                         ;

  wire fq6q87ocz4n3eh7tq_8l11kiq3xa = f1xe_xx4j29e7277py1p2k9uh & vfjafvqeepaxiqz2w76pl8ds6z
                         & eqce_y4zxdhu7zaz6s2fk7vec
                         ;

  wire te46hx1x_954f8oaiw8vpfl7 =
                           eqce_y4zxdhu7zaz6s2fk7vec
                         & m7frhh6dekyuotcrluw9m36kvn4
                         ;
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  

  
  
  
  
  wire zla7uqbb3yfvop1ja9 = c4ughu0qm5sfai;
  wire fnjtncb80f_1t9v1mn5;
  wire gf3aiywpsjayl9nw6y_rl_r;
  wire hsv3kgrb3c_k_9x6hb;
  wire syeryna6edz5he27_zgkify;
  
  ux607_gnrl_dffr #(1) k1twmto5d66302213o849gk (zla7uqbb3yfvop1ja9    , fnjtncb80f_1t9v1mn5, gf33atgy, ru_wi);
  ux607_gnrl_dffr #(1) kex7m81u0yuh1l9_kxujrpg3oh (fnjtncb80f_1t9v1mn5, gf3aiywpsjayl9nw6y_rl_r, gf33atgy, ru_wi);
  ux607_gnrl_dffr #(1) sy5z2392vbppdpknt27b1m6oph (gf3aiywpsjayl9nw6y_rl_r, hsv3kgrb3c_k_9x6hb, gf33atgy, ru_wi);
  ux607_gnrl_dffr #(1) uqzb7645ng6kxy8kb_a0knchg (hsv3kgrb3c_k_9x6hb, syeryna6edz5he27_zgkify, gf33atgy, ru_wi);
  

  
  wire raha4wzwsh_g_zg = (~indfp6mwqdqamez0mex) & syeryna6edz5he27_zgkify;
  
  wire nywm0kv90g64r5310wz = 
                 fnjtncb80f_1t9v1mn5 
               | gf3aiywpsjayl9nw6y_rl_r 
               | hsv3kgrb3c_k_9x6hb 
               | syeryna6edz5he27_zgkify ;

  wire eeopomndusb3z83b6;
  wire m1630hoivkgbkir3; 

  assign yb5ru177dkq2qb = 
                 zla7uqbb3yfvop1ja9 
               | nywm0kv90g64r5310wz
               | m1630hoivkgbkir3 
               | eeopomndusb3z83b6;
  


  wire [6-1:0] hequb9pd3bn5;

  wire fma8z0hm6f3uewn_vk = (~eeopomndusb3z83b6) & ( 
      
         raha4wzwsh_g_zg
         );

         
  wire oiagurkoxw3mq8p3y_ = eeopomndusb3z83b6;
  wire m04__f5senmr683gvg = fma8z0hm6f3uewn_vk | oiagurkoxw3mq8p3y_;
  wire [6-1:0] x2bla4_9fo9xl3 = 
                                   fma8z0hm6f3uewn_vk ? {6{1'b0}}
                                 : oiagurkoxw3mq8p3y_ ? (hequb9pd3bn5 + {{6-1{1'b0}},1'b1})
                                 : hequb9pd3bn5;
  
  ux607_gnrl_dfflr #(6) i9k9bvfdrefx9b12s8 (m04__f5senmr683gvg, x2bla4_9fo9xl3, hequb9pd3bn5, gf33atgy, ru_wi);
  
  localparam rjzg5aaa7ljdd2rk2ienn = (64 -1);

  assign m1630hoivkgbkir3 = fma8z0hm6f3uewn_vk;
  wire n81bejf_x7hih4c3m = oiagurkoxw3mq8p3y_ & (hequb9pd3bn5 == rjzg5aaa7ljdd2rk2ienn[6-1:0]);
  wire r59_bpoi9japjgeg = m1630hoivkgbkir3 | n81bejf_x7hih4c3m;
  wire m2ww3p90tivvcm2pxrs = m1630hoivkgbkir3;
  ux607_gnrl_dfflr #(1) qnytnrkz41zpef4ygemn (r59_bpoi9japjgeg, m2ww3p90tivvcm2pxrs, eeopomndusb3z83b6, gf33atgy, ru_wi);
  


  wire xpi9_z9vrvzc7gxt  = eeopomndusb3z83b6;
  
  wire xhumyr_ttpqs1x65 = oiagurkoxw3mq8p3y_;
  wire [6-1:0] eaa95xyq1761at3blmo = hequb9pd3bn5;
  wire [24-1:0] ej2juaulfcpj2lnfeqk6  = {24{1'b0}};
  wire                         f74vx9ulb9ziesmeh5   = 1'b1;

  localparam vf6oxg6vw87fiyq__ = (1 + 6 + 24 + 1);
  localparam t8lzfg9qlh_4kwovv7wj = (1 + 8 + 32 + 4);

  wire zf076ac19ivp1csbq2xy9;
  wire [6-1:0] nh60lylvhz65vcjxjzbsr;
  wire [24-1:0] vr6n0he4tf4xn8efytdl4 ;
  wire                         dma1vzh92la2k0k4944lxc2  ;

  wire lsxxcy5p3dky7il0f141w_b;
  wire [6-1:0] pcqyklmfrk69an1nr4tovexclx;
  wire [24-1:0] f6fhl3nngqjym1_ziugv10k ;
  wire                         hw9v3z65samnclk5dkj61h2  ;



  wire i3r6fyspyh4r6kc73en3;
  wire [r4bbs1l72_cd3t_-1:0] eni2zaouo2xcn1_r;

  wire ywx9or41ehj33tekj = eni2zaouo2xcn1_r[r4bbs1l72_cd3t_-1];


  wire jywzcibo3cb08kg0a; 
  wire soj2j1b62_nupmoszxl45_ip; 
  wire [27-1:0] k70vsrf3p8nx_vdlptr_247ei = erg8nrhaecoc2m5idim8fol1zo25m[(32-1):5];
  wire [6-1:0]    n78vaxm8ocds6eac     = k70vsrf3p8nx_vdlptr_247ei[6-1:0];
  assign zf076ac19ivp1csbq2xy9   = soj2j1b62_nupmoszxl45_ip ? i3r6fyspyh4r6kc73en3 : (i3r6fyspyh4r6kc73en3 & (~ywx9or41ehj33tekj));
  assign lsxxcy5p3dky7il0f141w_b   = soj2j1b62_nupmoszxl45_ip ? i3r6fyspyh4r6kc73en3 : (i3r6fyspyh4r6kc73en3 &   ywx9or41ehj33tekj );
  assign nh60lylvhz65vcjxjzbsr = soj2j1b62_nupmoszxl45_ip ? n78vaxm8ocds6eac : eni2zaouo2xcn1_r[6-1:0];
  assign pcqyklmfrk69an1nr4tovexclx = soj2j1b62_nupmoszxl45_ip ? n78vaxm8ocds6eac : eni2zaouo2xcn1_r[6-1:0];

  assign vr6n0he4tf4xn8efytdl4  = {24{1'b0}};
  assign f6fhl3nngqjym1_ziugv10k  = {24{1'b0}};
  assign dma1vzh92la2k0k4944lxc2   = 1'b0;
  assign hw9v3z65samnclk5dkj61h2   = 1'b0;



        


  
  
  
  
  wire ptmhu5qvej_2kw9w3pdr8;
  wire hgpmlnfjch5bm27n3zz3vd;
  wire nf6dcrwxlcch1sv8kmtkb_ry2;
  wire a3ybha5mrl8xcrr8;
  wire oyd54mosns8enc8c;

  wire [32-1:0] pb5q1jscnh9li4g_e5216b6; 
  assign pb5q1jscnh9li4g_e5216b6[5-1:0] = 5'b0;
  assign pb5q1jscnh9li4g_e5216b6[27+5-1:5] = {{(27-6){1'b0}}, nh60lylvhz65vcjxjzbsr};


  wire   ozi9s_ccjtrq6nogjymw         = (jywzcibo3cb08kg0a    ? qe0x130i0z960a1ld7jru7ma   : 1'b1               );
  wire   oi58e_8xo0iwnmf1b4uh         = (jywzcibo3cb08kg0a    ? z2w73ziehrytb1m0t4jo_jr0ici  : 1'b0               );
  wire   wok_5vlideqa4hy763          = (soj2j1b62_nupmoszxl45_ip ? 1'b1                      : 1'b0               );
  wire   dd_0zg96p33sc6t9l_         = (soj2j1b62_nupmoszxl45_ip ? qmpmjqpq_d69kzu6u9bxjr74w1y  : 1'b0               );
  wire   t02_wbi1amns3jes065sn        = (soj2j1b62_nupmoszxl45_ip ? e09r0m8969cj0sl6_iwpy513ad9kih : 1'b0               );
  wire   jjr4zhwlqoejhrtk6fe          = (soj2j1b62_nupmoszxl45_ip ? 1'b0                      : ywx9or41ehj33tekj    );
  wire   fa05x3xvuufk_8vwgwoazt9      = (soj2j1b62_nupmoszxl45_ip ? 1'b0                      : 1'b1               );

  assign ne3qv25fuqotk2dk5         = 1'b0;
  assign fsqkwjz0sanwked5rfthn       = ptmhu5qvej_2kw9w3pdr8     ;
  assign m5uxjf11e0v1munmybb1n3fv  = hgpmlnfjch5bm27n3zz3vd;
  assign eschp5gtzyhx77wg6jhl4z9ny  = nf6dcrwxlcch1sv8kmtkb_ry2;
  assign ycqmiyj7jekquq0pxuy1uk       = a3ybha5mrl8xcrr8     ;
  assign dryvl0kbql72b720rm       = oyd54mosns8enc8c     ;
  assign wo477hsguadhf4cwa9bbl      = 1'b0;
  assign fsfq1s74k43eb5l          = 1'b0;
  assign yajgwlnlp6hvh354akt3lm        = 1'b0;
  assign gec3f9o0vmsnfdwup7xem       = 64'b0   ;
  assign fy5zq5a7ou_6sownckex       = 8'b0   ;
  assign xopz5es01zuocuhfzv        = 1'b0              ;     
  assign j9ngo4gtwitbihmi5djct        = 1'b0              ;     
  assign hmaam0gy6lvgx07vlp6yo7        = 2'b0              ;
  assign foma9juy1lv_7626wum__ceu    = 1'b1;

  assign pte_y5zn1kqfnzxo5izs        = soj2j1b62_nupmoszxl45_ip ? erg8nrhaecoc2m5idim8fol1zo25m : pb5q1jscnh9li4g_e5216b6;

  
  
  
  wire xmvdvsjqgas1r79t0hvyff = dl1e0uq8c1swic;

  wire qnvhn5s48_vnk2s8ngqvxn6elox; 
  wire acejcdmkjp7hc3zmmmoz2j8;
  wire jhm5p8w5rzdzw1d835xkcnwqxdx0;

  wire dfqgbr7fyq0xiz172uj;

  assign qnvhn5s48_vnk2s8ngqvxn6elox = (~xmvdvsjqgas1r79t0hvyff) & dfqgbr7fyq0xiz172uj; 
  wire   tn9wx9b6b96ayt6kh5znx5     = (~xmvdvsjqgas1r79t0hvyff) & acejcdmkjp7hc3zmmmoz2j8; 

  assign stdkgs3cetkrgnprgzkr = dfqgbr7fyq0xiz172uj & tn9wx9b6b96ayt6kh5znx5;

  wire z1dt_7toi2ljqye_yupzbaffjpwvxqyqn = jhm5p8w5rzdzw1d835xkcnwqxdx0;


  wire jkqj750anrk85f54yke66h0yu_70teh5 = qnvhn5s48_vnk2s8ngqvxn6elox
                         ;

  assign acejcdmkjp7hc3zmmmoz2j8 =
                           jhm5p8w5rzdzw1d835xkcnwqxdx0
                         ;


  
  
  
  
  
  
  
  
  
  
  


  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  

  wire rrw0hjx1by8649e;
  wire eeu1a5x5fakgzef;
  wire u3dek804pblv01rwby3;
  wire nvzb52ltxbr826ffui6;
  wire cbjv6fberut9px0ext ;


  
  wire jkq984ky8fozrzq;
  wire wy8e7v3mv0oudza = (~rrw0hjx1by8649e) & (~cbjv6fberut9px0ext) & (~nvzb52ltxbr826ffui6) & (~u3dek804pblv01rwby3)  & (~jkq984ky8fozrzq);
  wire j1cskt8wmrapwcuwwwjwq = (~rrw0hjx1by8649e) &  (~cbjv6fberut9px0ext) & (~nvzb52ltxbr826ffui6) & (~jkq984ky8fozrzq) ;
  wire i1vah87l1fxh01choeoz2m4 = (~rrw0hjx1by8649e) &  (~nvzb52ltxbr826ffui6) & (~jkq984ky8fozrzq) ;
  wire e30rf6a88vykhuva14zjnu = (~rrw0hjx1by8649e) | jkq984ky8fozrzq; 
  wire i0ccgjn4_vexlacjblx = 1'b1 & (~jkq984ky8fozrzq) ;

  wire shj7yt_dr082bfdo0c6 = rrw0hjx1by8649e & i0ccgjn4_vexlacjblx;
  wire vvvr_o5rv85e56upfg_n = u3dek804pblv01rwby3 & j1cskt8wmrapwcuwwwjwq;
  wire i2cwubtp3ylg1ewfv   = cbjv6fberut9px0ext   & i1vah87l1fxh01choeoz2m4; 
  wire ufe4xjm3p1bk2gw0  = (nvzb52ltxbr826ffui6  & e30rf6a88vykhuva14zjnu) | jkq984ky8fozrzq;
  wire k88qugtn8ofr      = eeu1a5x5fakgzef      & wy8e7v3mv0oudza;   

  wire mkvubuawtidmr0qz =      
                      ( (vvvr_o5rv85e56upfg_n & u3dek804pblv01rwby3)
                      | (i2cwubtp3ylg1ewfv   & cbjv6fberut9px0ext  )
                      | (ufe4xjm3p1bk2gw0  & nvzb52ltxbr826ffui6 )
                      | (shj7yt_dr082bfdo0c6  & rrw0hjx1by8649e )
                      | (k88qugtn8ofr      & eeu1a5x5fakgzef     )); 

  wire had01mmuqyc8tzrxd5;
  wire w0dzgnd8l98an1zx6ijhlbtalpk;

  assign eeu1a5x5fakgzef              = p0brv6fqgdvccaui21k8;
  assign f56j5y58ce35hwpqbnu16 = had01mmuqyc8tzrxd5 & wy8e7v3mv0oudza;

  assign u3dek804pblv01rwby3       = jkqj750anrk85f54yke66h0yu_70teh5;
  assign jhm5p8w5rzdzw1d835xkcnwqxdx0 = had01mmuqyc8tzrxd5 & j1cskt8wmrapwcuwwwjwq;

  assign nvzb52ltxbr826ffui6         = w0dzgnd8l98an1zx6ijhlbtalpk;
  wire   vt1176n4bhzdaz39cel8dhxqwrawhf = had01mmuqyc8tzrxd5 & e30rf6a88vykhuva14zjnu;

  assign cbjv6fberut9px0ext         = dq71bajnhqrbc7pjo3ilkqpu00atil;
  assign y85uyrjj282xf9p3it0u2wvmixet = had01mmuqyc8tzrxd5 & i1vah87l1fxh01choeoz2m4;

  assign rrw0hjx1by8649e         = rguv86jfrc_9hefk7y2yvxn6og4d1;
  assign ra61k0r5_z16sciiz8un534o6w = had01mmuqyc8tzrxd5 & i0ccgjn4_vexlacjblx;

  wire i6z74pebe0ra5htg2uo;
  wire me3trrsw6wqsrh6w4;

  wire [6-1:0] l_0u_48a8iuyaal7qgl;
  wire [6-1:0] rf99quy5w7mi_qa748z;

  wire [24-1:0] o33xxeetwtdlelf04 ;
  wire                         khvu04h61q09inc_6  ;
  wire [24-1:0] mnwvvetpxt3aayw4htb59 ;
  wire                         n0tel4727bjok_zrc  ;



  wire                           e3rxl7mic_dpejl98_ts2;  
  wire  [6-1:0]  dlxukfkm1k19y_gskjb9vnl;
  wire                           sdmu0iskkbwi6blvi5 ;
  wire  [24-1:0]  suwghvh7qn2812e0i1b3he4;          
   
  wire                           ejddc553ql3y8eh4p8zbx9;  
  wire  [6-1:0]  gt8340_0a15il23cs0dyfy; 
  wire                           rocadn0agggbhe8c7k6f ;
  wire  [24-1:0]  wa8alqpvm8_8wqh82v4;          

  wire                           xd358a2nj1otzbd40o73xb;  
  wire  [6-1:0]  mx268wfdr27bxvwnmmo;
  wire                           wftjq44g43xvkg428 ;
  wire  [24-1:0]  dxze5eqmhutphmuxctr;          
   
  wire                           akuzoy0x17uo4jeh1_kpe;  
  wire  [6-1:0]  xtwgwqnfhzoh7z4upxshz6y; 
  wire                           rhlr3nyozzrn6fofxgxji0 ;
  wire  [24-1:0]  or9rw5q8w0eistsrkf;          


  wire                           gg8smz7g8ompdkylfsii;  
  wire  [6-1:0]  y_4c2_1ibmz5t6q3cxlkbc25;
  wire                           bc73rkmzmuniy5r6c7jvi ;
  wire  [24-1:0]  vkqnes_n9nib643hgr;          
   
  wire                           vfwv2h15g194_9vp6v0qj6;  
  wire  [6-1:0]  hy9oy2mo1t8mvphwqkiipyi9; 
  wire                           v12kpdmdljqz6v4yd_fh5p ;
  wire  [24-1:0]  kahkbbr9p728erz9ilfg;          


  wire jgeyki3wp7rzhsh958;
  wire                          nsc0elm1w3m_inebi5nie51  ;
  wire                          kbae6svksx713v4pbhv8  ;
  wire [6-1:0]  hgfb_gwm97sz53betsjyk5;
  wire [6-1:0]  ee18h0eqehcvi043ns32gf;
  wire                          qxdc_js0dtaug304lp11_gu  ;
  wire                          tarnkvmavl9287x895  ;
  wire [24-1:0]  bshid8lzm3x5d3ju1u82v ;
  wire [24-1:0]  wuf4wr1vape2nd15r20p ;
 



  assign { 
           mum8f1rtatle7p_55y84   
         , pn5bpwlp5ijfako9m5ao 
         , a1rl4lmhqp8ydyk07kqkn  
         , g3s0qe2adsxsx8e6z    
         , pmz7e4mgvbnmimqp0nghk   
         , j61algpxjoycxbswhgsuf 
         , fbv1q6sraswzp91zcn  
         , omq1ehm8hp4q9jgp5n5vn    
         } = 
                 k88qugtn8ofr ? 
                            { 
                  i6z74pebe0ra5htg2uo   , l_0u_48a8iuyaal7qgl , o33xxeetwtdlelf04  , khvu04h61q09inc_6  
                , me3trrsw6wqsrh6w4   , rf99quy5w7mi_qa748z , mnwvvetpxt3aayw4htb59  , n0tel4727bjok_zrc  
                } : (
                    (
                      {2*vf6oxg6vw87fiyq__{ufe4xjm3p1bk2gw0}} & {
                                                            e3rxl7mic_dpejl98_ts2 , dlxukfkm1k19y_gskjb9vnl , suwghvh7qn2812e0i1b3he4  , sdmu0iskkbwi6blvi5   
                                                          , ejddc553ql3y8eh4p8zbx9 , gt8340_0a15il23cs0dyfy , wa8alqpvm8_8wqh82v4  , rocadn0agggbhe8c7k6f  
                              }
                    ) | 
                    (
                      {2*vf6oxg6vw87fiyq__{i2cwubtp3ylg1ewfv}} & {
                                                            gg8smz7g8ompdkylfsii , y_4c2_1ibmz5t6q3cxlkbc25 , vkqnes_n9nib643hgr  , bc73rkmzmuniy5r6c7jvi   
                                                          , vfwv2h15g194_9vp6v0qj6 , hy9oy2mo1t8mvphwqkiipyi9 , kahkbbr9p728erz9ilfg  , v12kpdmdljqz6v4yd_fh5p 
                              }
                    ) | 
                    (
                      {2*vf6oxg6vw87fiyq__{shj7yt_dr082bfdo0c6}} & {
                                                            xd358a2nj1otzbd40o73xb   , mx268wfdr27bxvwnmmo , dxze5eqmhutphmuxctr  , wftjq44g43xvkg428   
                                                          , akuzoy0x17uo4jeh1_kpe   , xtwgwqnfhzoh7z4upxshz6y , or9rw5q8w0eistsrkf  , rhlr3nyozzrn6fofxgxji0  
                              }
                    ) |    
                    (
                      {2*vf6oxg6vw87fiyq__{vvvr_o5rv85e56upfg_n}} & {
                                                            zf076ac19ivp1csbq2xy9   , nh60lylvhz65vcjxjzbsr , vr6n0he4tf4xn8efytdl4  , dma1vzh92la2k0k4944lxc2   
                                                          , lsxxcy5p3dky7il0f141w_b   , pcqyklmfrk69an1nr4tovexclx , f6fhl3nngqjym1_ziugv10k  , hw9v3z65samnclk5dkj61h2  
                              }
                    ) |    
                    (
                      {2*vf6oxg6vw87fiyq__{xpi9_z9vrvzc7gxt}} & {
                                                            xhumyr_ttpqs1x65   , eaa95xyq1761at3blmo , ej2juaulfcpj2lnfeqk6  , f74vx9ulb9ziesmeh5   
                                                          , xhumyr_ttpqs1x65   , eaa95xyq1761at3blmo , ej2juaulfcpj2lnfeqk6  , f74vx9ulb9ziesmeh5  
                              }
                    ) |    
                    (
                    
                      {2*vf6oxg6vw87fiyq__{jgeyki3wp7rzhsh958}} & {
                                                            nsc0elm1w3m_inebi5nie51 , hgfb_gwm97sz53betsjyk5, bshid8lzm3x5d3ju1u82v, qxdc_js0dtaug304lp11_gu     
                                                          , kbae6svksx713v4pbhv8 , ee18h0eqehcvi043ns32gf, wuf4wr1vape2nd15r20p, tarnkvmavl9287x895    
                              }
                    )    

                  );

  
  
  
  
  
  
  
  
  
  
  
  
  
  
  

  wire rwqdh9w472dna;
  wire jq7e16ojaaz1ur04t47;
  wire dpwkelsg4w4rf28ny1u9;
  wire vnglpee2kb7x4v3e2b6 ;

  
  wire e4y_8hurgo98x4wemt = (~dpwkelsg4w4rf28ny1u9) & (~jq7e16ojaaz1ur04t47) & (~vnglpee2kb7x4v3e2b6)  & (~jkq984ky8fozrzq); 
  wire t1nuj0z_9rltyuyp0gm = (~dpwkelsg4w4rf28ny1u9) & (~jq7e16ojaaz1ur04t47) & (~jkq984ky8fozrzq) ;
  wire xrat1gwekt44mcw32uw94 = (~jq7e16ojaaz1ur04t47) | jkq984ky8fozrzq;
  wire dof2qdvmkc2rssai2hb1u6 = 1'b1 & (~jkq984ky8fozrzq);


  wire ao36lev_ys2bw97s   = vnglpee2kb7x4v3e2b6   & t1nuj0z_9rltyuyp0gm; 
  wire yeo9u3v77n2dimne  = (dpwkelsg4w4rf28ny1u9  & xrat1gwekt44mcw32uw94) | jkq984ky8fozrzq;
  wire eaux4rpzn5avq66   = jq7e16ojaaz1ur04t47   & dof2qdvmkc2rssai2hb1u6;
  wire btmvep9nehgs      = rwqdh9w472dna      & e4y_8hurgo98x4wemt;   

  wire gw1nu9da4hehn0n1 = 
  
                 had01mmuqyc8tzrxd5 
  
               | (~brfek3hm0m1h_0qdx) 
               ;

  wire kcvmtch763q8ina8s4zil7kyspcf0;

  assign rwqdh9w472dna             = j30h3wzip_eqif46u34tw4;
  assign nk4gkqhhy_a4hc5n4kin = gw1nu9da4hehn0n1 & e4y_8hurgo98x4wemt;

  assign jq7e16ojaaz1ur04t47      = fq6q87ocz4n3eh7tq_8l11kiq3xa;
  assign ujuhwx1rtmvxjxxpbmlhcttboa3kd = gw1nu9da4hehn0n1 & dof2qdvmkc2rssai2hb1u6;

  assign vnglpee2kb7x4v3e2b6               = jo20b3jp2h86mzvqeae5j3xsu3g3;
  assign ijsk41ad4tvq4zse7kouzpbxcnck2 = gw1nu9da4hehn0n1 & t1nuj0z_9rltyuyp0gm;

  assign dpwkelsg4w4rf28ny1u9           = kcvmtch763q8ina8s4zil7kyspcf0;
  wire   wyyj6g00owlp1khb6vv9ycavglf = gw1nu9da4hehn0n1 & xrat1gwekt44mcw32uw94;
  
  wire                            vqk9s6vdwj03b1nk46;  
  wire  [8-1:0]  ftxo1913pi2k8gqfhhzalo; 
  wire  [4-1:0]  kbxf845povp5e5witzqjk;
  wire  [32-1:0]  a7nsr8tm_g5p5yek17ff7i;          
                                  
  wire                            rtl6pef_7afwbyimpdzz;  
  wire  [8-1:0]  n_mnmtuwkqc34kiucl1t5c; 
  wire  [4-1:0]  fuy5xpvy57_bb_r7h_;
  wire  [32-1:0]  x6gmclknmv0wspuem14db76;          
                                 
  wire                            lasdt5zxlelolfv4i;  
  wire  [8-1:0]  ixvdqtu1o_7q05drk9p; 
  wire  [4-1:0]  lvk3p1ksfy64il0ktw2w;
  wire  [32-1:0]  y4v98fdt14u2fg0kn_eiuco;          
                     
  wire                            ce1xag7wxa_l0irqi;  
  wire  [8-1:0]  h8g_w8qo3vwr23j57mitm9o; 
  wire  [4-1:0]  hsx_qko4lqeerbg1jt22jlw;
  wire  [32-1:0]  roczx_v0ys9xuqcq68sa;

  wire                            zffkoq91x2yrt8idy12;  
  wire  [8-1:0]  cw8g0z3xpl_jmzl0bqsr4qz7r; 
  wire  [4-1:0]  c3o9e_kce6dj_oses5ebis;
  wire  [32-1:0]  nl6qyr_h4vq399gjb47;          
                                   
  wire                            ywnbexiz4zyc0xfli8;  
  wire  [8-1:0]  fe0_jbuekwa1u_igwcjrf5; 
  wire  [4-1:0]  ezoxoh6x_6pp3kplit2ipzy;
  wire  [32-1:0]  merrnyoykrdknka8adx1kp;          
                                  
  wire                            g0zewsbtm0xx173b6w3n;  
  wire  [8-1:0]  ks8_k_t4av7jsxfssailx; 
  wire  [4-1:0]  fuqvy5sh_dgu5b6_k5te2;
  wire  [32-1:0]  s5br9ji17fis2ai4t5b257ui;          
                     
  wire                            opg7to8zm4fdk0kbxb;  
  wire  [8-1:0]  xuch6yvcgtv5auc_2s5g32; 
  wire  [4-1:0]  c3es5lys6yhd7wv8lg2ho553;
  wire  [32-1:0]  buo4rvqs58con3m3n965h6a;          

  wire                            gymo5upuuufrkiu0g;  
  wire  [8-1:0]  yfl3z2gjyii2os6js5u7xux; 
  wire  [4-1:0]  l1wuw4784zfpjcxv_tv9f;
  wire  [32-1:0]  nxzxonv_ne6j0bo_bhtel;          
                                  
  wire                            qpdcndj__mjjubf4;  
  wire  [8-1:0]  pd_1u9zwdqqbxjs9ba7g; 
  wire  [4-1:0]  rysv66sonr6uldbb379uf;
  wire  [32-1:0]  gl2h7cy3yftrtcdjqht;          
                                 
  wire                            xhtjh5yqah1skcehze;  
  wire  [8-1:0]  jk41isdbxrtauo9gcxyyo; 
  wire  [4-1:0]  ip8kc5qycn6__tojwd;
  wire  [32-1:0]  ywswe20ycctmqeo1qkgm8a;          
                     
  wire                            bdl_fud5zqzxlabhb2q;  
  wire  [8-1:0]  ythxm8b2m6qm86g5j_4hvbl; 
  wire  [4-1:0]  jihrna79l86fvm3tvhrx;
  wire  [32-1:0]  heqnwxy0x0uw2nv8r;

  wire                            cswt3kuajv3zxjj3royb;  
  wire  [8-1:0]  yt6fnikwf0c8ztaq91rwz; 
  wire  [4-1:0]  yi50g8outdxmqa4e2uo;
  wire  [32-1:0]  zc6u0jmmj3gkj9vgxdgt;          
                                  
  wire                            wtjfz_620cbhzvtnyosm;  
  wire  [8-1:0]  nn9f5y1j5r_u_pwa3ye; 
  wire  [4-1:0]  y44utukerytn8bcnd7cxi3;
  wire  [32-1:0]  iggkgmc7p_70htdrjtf6gv1;          
                                 
  wire                            qyje8_wx1y6nov9nt;  
  wire  [8-1:0]  u4h_rc_dg1scnmq0la4tyyim; 
  wire  [4-1:0]  v8fwqjnng9vhsymrb3jc3p;
  wire  [32-1:0]  qwkfrhebeat5x3r6tdd464;          
                     
  wire                            u9pufmsi7150uxn_9uqxp5;  
  wire  [8-1:0]  yedl9u82iubd5w_uw3zfm9y; 
  wire  [4-1:0]  x3jcl5fq5odurkfmee9ncr0;
  wire  [32-1:0]  lmqzp5jgcehv098rwtxpu;   


  assign { 
           qgl4363n31jx6xjyo05zkn   , zec78nyllxlfwmpsgncluudf , gngmcj5c1jd85csel9ntru  , dwvnjl0vxqkgd8t6dtvg5z   
         , km7co8hqm563od8ga_03_g   , j4mas6g26o63wvnsdquh8c4p , rcy_v3911lf33nza5j  , nniah5mh0cunkhyln9   
         , xzgkclcxsgfuseg87   , djwlah5bo0r6myit6cal0t , dydwz9i6k80alqfarffop  , qu_ju3lv6nvkdbo8h11uf   
         , kp2j8kv1p1cjcg0lerwm   , v4a7g1wh3ivw0esp7dye0oiz , n_h5oz0c5bo5rpevwjcu8  , x9zuk21gpaj58uszvm5   
         } = 
                 btmvep9nehgs ? 
                            { 
                  gymo5upuuufrkiu0g   , yfl3z2gjyii2os6js5u7xux , nxzxonv_ne6j0bo_bhtel  , l1wuw4784zfpjcxv_tv9f 
                , qpdcndj__mjjubf4   , pd_1u9zwdqqbxjs9ba7g , gl2h7cy3yftrtcdjqht  , rysv66sonr6uldbb379uf 
                , xhtjh5yqah1skcehze   , jk41isdbxrtauo9gcxyyo , ywswe20ycctmqeo1qkgm8a  , ip8kc5qycn6__tojwd 
                , bdl_fud5zqzxlabhb2q   , ythxm8b2m6qm86g5j_4hvbl , heqnwxy0x0uw2nv8r  , jihrna79l86fvm3tvhrx 
                } : (
                    (
                      {4*t8lzfg9qlh_4kwovv7wj{eaux4rpzn5avq66}} & {
                                                            vqk9s6vdwj03b1nk46   , ftxo1913pi2k8gqfhhzalo , a7nsr8tm_g5p5yek17ff7i  , kbxf845povp5e5witzqjk 
                                                          , rtl6pef_7afwbyimpdzz   , n_mnmtuwkqc34kiucl1t5c , x6gmclknmv0wspuem14db76  , fuy5xpvy57_bb_r7h_ 
                                                          , lasdt5zxlelolfv4i   , ixvdqtu1o_7q05drk9p , y4v98fdt14u2fg0kn_eiuco  , lvk3p1ksfy64il0ktw2w 
                                                          , ce1xag7wxa_l0irqi   , h8g_w8qo3vwr23j57mitm9o , roczx_v0ys9xuqcq68sa  , hsx_qko4lqeerbg1jt22jlw 
                              }
                    ) |  

                    (
                      {4*t8lzfg9qlh_4kwovv7wj{yeo9u3v77n2dimne}} & {
                                                            zffkoq91x2yrt8idy12 , cw8g0z3xpl_jmzl0bqsr4qz7r , nl6qyr_h4vq399gjb47  , c3o9e_kce6dj_oses5ebis 
                                                          , ywnbexiz4zyc0xfli8 , fe0_jbuekwa1u_igwcjrf5 , merrnyoykrdknka8adx1kp  , ezoxoh6x_6pp3kplit2ipzy 
                                                          , g0zewsbtm0xx173b6w3n , ks8_k_t4av7jsxfssailx , s5br9ji17fis2ai4t5b257ui  , fuqvy5sh_dgu5b6_k5te2 
                                                          , opg7to8zm4fdk0kbxb , xuch6yvcgtv5auc_2s5g32 , buo4rvqs58con3m3n965h6a  , c3es5lys6yhd7wv8lg2ho553 
                              }
                    ) | 
                    (
                      {4*t8lzfg9qlh_4kwovv7wj{ao36lev_ys2bw97s}} & {
                                                            cswt3kuajv3zxjj3royb , yt6fnikwf0c8ztaq91rwz , zc6u0jmmj3gkj9vgxdgt  , yi50g8outdxmqa4e2uo 
                                                          , wtjfz_620cbhzvtnyosm , nn9f5y1j5r_u_pwa3ye , iggkgmc7p_70htdrjtf6gv1  , y44utukerytn8bcnd7cxi3 
                                                          , qyje8_wx1y6nov9nt , u4h_rc_dg1scnmq0la4tyyim , qwkfrhebeat5x3r6tdd464  , v8fwqjnng9vhsymrb3jc3p 
                                                          , u9pufmsi7150uxn_9uqxp5 , yedl9u82iubd5w_uw3zfm9y , lmqzp5jgcehv098rwtxpu  , x3jcl5fq5odurkfmee9ncr0 
                              }
                    )   
                            );

 





  
  
  
  
  

  wire [5-1:0]      wb5io39sh3kw47crv    = a7h_7269eov[4:0];
  wire [27-1:0]   dbcliz7z9p4m24h2c_jr = a7h_7269eov[(32-1):5];
  
  wire [6-1:0]      r1taf2aepfbvol5 = dbcliz7z9p4m24h2c_jr[6-1:0];
  wire [21-1:0]        v1ysponf94idgs4u45 = dbcliz7z9p4m24h2c_jr[27-1:6];
  
  
  assign i6z74pebe0ra5htg2uo  = jo2m0mwneyhm & p0brv6fqgdvccaui21k8;
  assign me3trrsw6wqsrh6w4  = jo2m0mwneyhm & p0brv6fqgdvccaui21k8;
  assign gg8smz7g8ompdkylfsii = u3gm9gusc9log5m42rc & dq71bajnhqrbc7pjo3ilkqpu00atil;
  assign vfwv2h15g194_9vp6v0qj6 = u3gm9gusc9log5m42rc & dq71bajnhqrbc7pjo3ilkqpu00atil;

  wire   dfg63fb5pt1ns8gd = jo2m0mwneyhm & j30h3wzip_eqif46u34tw4 ;
  wire   ty2urjgi6le0cxqumorte = u3gm9gusc9log5m42rc & jo20b3jp2h86mzvqeae5j3xsu3g3 ;


  
  assign l_0u_48a8iuyaal7qgl = r1taf2aepfbvol5;
  assign rf99quy5w7mi_qa748z = r1taf2aepfbvol5;

  assign o33xxeetwtdlelf04  = {24{1'b0}}; 
  assign khvu04h61q09inc_6   = 1'b0;
  assign mnwvvetpxt3aayw4htb59  = {24{1'b0}}; 
  assign n0tel4727bjok_zrc   = 1'b0;


  assign nxzxonv_ne6j0bo_bhtel  = {32{1'b0}}; 
  assign l1wuw4784zfpjcxv_tv9f  = {4{1'b0}};
  assign gl2h7cy3yftrtcdjqht  = {32{1'b0}}; 
  assign rysv66sonr6uldbb379uf  = {4{1'b0}};
  assign ywswe20ycctmqeo1qkgm8a  = {32{1'b0}}; 
  assign ip8kc5qycn6__tojwd  = {4{1'b0}};
  assign heqnwxy0x0uw2nv8r  = {32{1'b0}}; 
  assign jihrna79l86fvm3tvhrx  = {4{1'b0}};


  suzytsmnh3c_jk3y2hekvvubgi ebxzmphnvpg56bv44r0(
    .vhqr9jgt5       (dfg63fb5pt1ns8gd),

    .u4amtcbhq_6g6rx9 (r1taf2aepfbvol5),
    .sm0ktbr6as2sl7ho(wb5io39sh3kw47crv),

    .rl_3d1m7gcc0    (gymo5upuuufrkiu0g),
    .tsdapc3y0fh    (qpdcndj__mjjubf4),
    .mohep6fqp67x    (xhtjh5yqah1skcehze),
    .mmmu7pm6e_uqx    (bdl_fud5zqzxlabhb2q),

    .e_9jhaby2__46fj  (yfl3z2gjyii2os6js5u7xux),
    .lpcj6ymxsst2n  (pd_1u9zwdqqbxjs9ba7g),
    .wdb90nca460cp  (jk41isdbxrtauo9gcxyyo),
    .rin3amuhzyhjgg  (ythxm8b2m6qm86g5j_4hvbl)
  );

  
  
  
  
  
  wire [5-1:0]      wkz_4r2zmdu604l20n79kp    = fwgc_k58kjyp_va[4:0];
  wire [27-1:0]   hl94ul8nkhs8bqdszlda6gb = fwgc_k58kjyp_va[(32-1):5];
  
  wire [6-1:0]      l_gbxjnkkjjvhh5akwe = hl94ul8nkhs8bqdszlda6gb[6-1:0];
  wire [21-1:0]        fc32tw88qkmrzqw2j4alcvi = hl94ul8nkhs8bqdszlda6gb[27-1:6];
  

  
  assign y_4c2_1ibmz5t6q3cxlkbc25 = l_gbxjnkkjjvhh5akwe;
  assign hy9oy2mo1t8mvphwqkiipyi9 = l_gbxjnkkjjvhh5akwe;

  assign vkqnes_n9nib643hgr  = {24{1'b0}}; 
  assign bc73rkmzmuniy5r6c7jvi   = 1'b0;
  assign kahkbbr9p728erz9ilfg  = {24{1'b0}}; 
  assign v12kpdmdljqz6v4yd_fh5p   = 1'b0;


  assign zc6u0jmmj3gkj9vgxdgt  = {32{1'b0}}; 
  assign yi50g8outdxmqa4e2uo  = {4{1'b0}};
  assign iggkgmc7p_70htdrjtf6gv1  = {32{1'b0}}; 
  assign y44utukerytn8bcnd7cxi3  = {4{1'b0}};
  assign qwkfrhebeat5x3r6tdd464  = {32{1'b0}}; 
  assign v8fwqjnng9vhsymrb3jc3p  = {4{1'b0}};
  assign lmqzp5jgcehv098rwtxpu  = {32{1'b0}}; 
  assign x3jcl5fq5odurkfmee9ncr0  = {4{1'b0}};


  suzytsmnh3c_jk3y2hekvvubgi wienzg88s7vmyfqhixj(
    .vhqr9jgt5       (ty2urjgi6le0cxqumorte),

    .u4amtcbhq_6g6rx9 (l_gbxjnkkjjvhh5akwe),
    .sm0ktbr6as2sl7ho(wkz_4r2zmdu604l20n79kp),

    .rl_3d1m7gcc0    (cswt3kuajv3zxjj3royb),
    .tsdapc3y0fh    (wtjfz_620cbhzvtnyosm),
    .mohep6fqp67x    (qyje8_wx1y6nov9nt),
    .mmmu7pm6e_uqx    (u9pufmsi7150uxn_9uqxp5),

    .e_9jhaby2__46fj  (yt6fnikwf0c8ztaq91rwz),
    .lpcj6ymxsst2n  (nn9f5y1j5r_u_pwa3ye),
    .wdb90nca460cp  (u4h_rc_dg1scnmq0la4tyyim),
    .rin3amuhzyhjgg  (yedl9u82iubd5w_uw3zfm9y)
  );

  
  
  
  
  wire                         y4z10x_uk5tx9gjpp;  
  wire [3-1:0] vt4fxo524ecd4y832detyma;  
  wire [32-1:0]   cb39rlyxl60nbkm;  
  wire [64-1:0]      c3h8wzh_yyz3847v; 
  wire [8-1:0]      zz8qhy80jaf147ase;

  wire [5-1:0]      fph7zc9jyjpn03_hd1z04sa04    = cb39rlyxl60nbkm[4:0];
  wire [27-1:0]   a2w11qavrtvinkcl_25iiu_b_ = cb39rlyxl60nbkm[(32-1):5];
  
  wire [6-1:0]      w7q6rcy2teneytmuos7dufv8 = a2w11qavrtvinkcl_25iiu_b_[6-1:0];
  wire [21-1:0]        uibl3zc1u490w_3zyw0 = a2w11qavrtvinkcl_25iiu_b_[27-1:6];
  

  wire lgdhsk7cwbxgrv43;


  uy3gep77czajwdyrmq3ed7su xkraalw_hv78wxnkn213ou(
    .s71tjwwz         (y4z10x_uk5tx9gjpp),
    .vhqr9jgt5       (lgdhsk7cwbxgrv43),
    .mm89bcd_zxeoe1y    (c3h8wzh_yyz3847v),
    .amz4453y8nx6q    (zz8qhy80jaf147ase),

    .u4amtcbhq_6g6rx9 (w7q6rcy2teneytmuos7dufv8),
    .sm0ktbr6as2sl7ho(fph7zc9jyjpn03_hd1z04sa04),

    .rl_3d1m7gcc0    (vqk9s6vdwj03b1nk46),
    .tsdapc3y0fh    (rtl6pef_7afwbyimpdzz),
    .mohep6fqp67x    (lasdt5zxlelolfv4i),
    .mmmu7pm6e_uqx    (ce1xag7wxa_l0irqi),

    .e_9jhaby2__46fj  (ftxo1913pi2k8gqfhhzalo),
    .lpcj6ymxsst2n  (n_mnmtuwkqc34kiucl1t5c),
    .wdb90nca460cp  (ixvdqtu1o_7q05drk9p),
    .rin3amuhzyhjgg  (h8g_w8qo3vwr23j57mitm9o),

    .e6rwnjewsq6s6oro  (a7nsr8tm_g5p5yek17ff7i),
    .u74ed5k2tobo  (x6gmclknmv0wspuem14db76),
    .cthiem_1bgmj  (y4v98fdt14u2fg0kn_eiuco),
    .dg5w1zgjmlq1a4n  (roczx_v0ys9xuqcq68sa),

    .ft2vjq7oh7l1hzqu  (kbxf845povp5e5witzqjk),
    .wbr3gkcxil8f_hgq  (fuy5xpvy57_bb_r7h_),
    .t1ncj092lli  (lvk3p1ksfy64il0ktw2w),
    .vhh7ujoe4fwn_8  (hsx_qko4lqeerbg1jt22jlw)
  );



  
  assign zylypzxl2r1asy4_sbdielf_2 = vt4fxo524ecd4y832detyma[1];

  wire reh5cltwd1u892j7xoky2sp =   y4z10x_uk5tx9gjpp  & lgdhsk7cwbxgrv43;
  wire c6aixo29buw824jvkxx0ylg4 = (~y4z10x_uk5tx9gjpp) & lgdhsk7cwbxgrv43;

  assign xd358a2nj1otzbd40o73xb = reh5cltwd1u892j7xoky2sp & (~zylypzxl2r1asy4_sbdielf_2);  
  assign akuzoy0x17uo4jeh1_kpe = c6aixo29buw824jvkxx0ylg4 & (~zylypzxl2r1asy4_sbdielf_2);  

  assign mx268wfdr27bxvwnmmo = w7q6rcy2teneytmuos7dufv8; 
  assign xtwgwqnfhzoh7z4upxshz6y = w7q6rcy2teneytmuos7dufv8; 

  assign wftjq44g43xvkg428  = 1'b1;
  assign rhlr3nyozzrn6fofxgxji0  = 1'b1;

  wire [24-1:0] rrkco7gwh3mt7saebiigt0ocgs_ = {vt4fxo524ecd4y832detyma, uibl3zc1u490w_3zyw0}; 
  assign dxze5eqmhutphmuxctr = (((24'b010<<21) & {24{1'b1}}) | ((~(24'b010<<21)) & rrkco7gwh3mt7saebiigt0ocgs_));
  assign or9rw5q8w0eistsrkf = (((24'b010<<21) & {24{1'b1}}) | ((~(24'b010<<21)) & rrkco7gwh3mt7saebiigt0ocgs_));


  
  
  
  
  
  
  
  
  
  
  
  
  
  

  localparam hxhz0y3mpud0ey59v = (f16zrowg1s1f5+12);

  wire [hxhz0y3mpud0ey59v-1:0] ukllsj0e1xzeouqnrx;

  wire dbkpihmr6104_e36q4zoxpgy  ;
  wire gxv5oxyuuit9f6lci1p0v22   ;
  wire bfrlc8tog574i131socryaap  ;
  wire v5rjtrkyv236_aeycevjw  ;
  wire v14gd4036xa4fahc_461n ;
  wire ti3tf23yq0i6r0hmenfl6   ;

  assign ukllsj0e1xzeouqnrx = (
                            ( {hxhz0y3mpud0ey59v{k88qugtn8ofr}} & {
                                           1'b1
                                         , 1'b0
                                         , 1'b0
                                         , 1'b0
                                         , 1'b0
                                         , 1'b0
                                         , 1'b0
                                         , 1'b0
                                         , 1'b0
                                         , 1'b0
                                         , 1'b0
                                         , 1'b0
                                         , se0zyj4n4upz  
                                         } 
                            )
                          | ( {hxhz0y3mpud0ey59v{vvvr_o5rv85e56upfg_n}} & {
                                           1'b0
                                         , 1'b1
                                         , 1'b0
                                         , 1'b0
                                         , 1'b0
                                         , ozi9s_ccjtrq6nogjymw  
                                         , wok_5vlideqa4hy763  
                                         , dd_0zg96p33sc6t9l_  
                                         , t02_wbi1amns3jes065sn  
                                         , oi58e_8xo0iwnmf1b4uh  
                                         , jjr4zhwlqoejhrtk6fe  
                                         , fa05x3xvuufk_8vwgwoazt9  
                                         , cdqzid8vpi25lg6fx  
                                         } 
                            )
                          | ( {hxhz0y3mpud0ey59v{ufe4xjm3p1bk2gw0}} & {
                                           1'b0
                                         , 1'b0
                                         , 1'b1
                                         , 1'b0
                                         , 1'b0
                                         , 1'b0
                                         , 1'b0
                                         , 1'b0
                                         , 1'b0
                                         , 1'b0
                                         , 1'b0
                                         , 1'b0
                                         , k8qtf1i196m8bfpmqi  
                                         } 
                            )
                          | ( {hxhz0y3mpud0ey59v{i2cwubtp3ylg1ewfv}} & {
                                           1'b0
                                         , 1'b0
                                         , 1'b0
                                         , 1'b1
                                         , 1'b0
                                         , dbkpihmr6104_e36q4zoxpgy  
                                         , gxv5oxyuuit9f6lci1p0v22  
                                         , v5rjtrkyv236_aeycevjw  
                                         , v14gd4036xa4fahc_461n  
                                         , bfrlc8tog574i131socryaap  
                                         , ti3tf23yq0i6r0hmenfl6  
                                         , v_9kfy4x1fk3adyoz6x2
                                         , ky8zw277b8fa1dq1zk  
                                         } 
                            )
                          | ( {hxhz0y3mpud0ey59v{shj7yt_dr082bfdo0c6}} & {
                                           1'b0
                                         , 1'b0
                                         , 1'b0
                                         , 1'b0
                                         , 1'b1
                                         , 1'b0
                                         , 1'b0
                                         , 1'b0
                                         , 1'b0
                                         , 1'b0
                                         , 1'b0
                                         , 1'b0
                                         , tvypfoh27qvczot  
                                         } 
                            )
                     );

  wire kggnqtwc1ljww3tnze     ; 
  wire mih7nmwcak45d8a2hvfx; 
  wire z_c9c063dzhr5i2tflx1ge ;
  wire gxctvntt6usn533wgnh6  ;
  wire xa74n2vq7asiuic23w  ;

  wire tftxelzlbcv3nmg0ry     ; 
  wire c7l7vyum1z06i355gent; 
  wire d42b0dgiiybnaa647lv9euj ;
  wire rx250nlkrd2m3gkhtzzl  ;

  wire [hxhz0y3mpud0ey59v-1:0] ysoarmlp98243p;

  wire ie6x4201u8jyqlgs    ;  
  wire vfzxxuugm86jff_8iod     ;  
  wire qu2oxvm9fx85hbf    ;
  wire fyqztmgm7gm2uol7   ;
  wire auhnvtbztby6o4qy646    ;
  wire u6xz15_qx1lay5yvg     ;
  wire xj0hdx62yzgvd1qvsf ; 

  assign {
           kggnqtwc1ljww3tnze 
         , mih7nmwcak45d8a2hvfx 
         , z_c9c063dzhr5i2tflx1ge 
         , gxctvntt6usn533wgnh6  
         , xa74n2vq7asiuic23w  
         , ie6x4201u8jyqlgs  
         , vfzxxuugm86jff_8iod  
         , qu2oxvm9fx85hbf  
         , fyqztmgm7gm2uol7  
         , auhnvtbztby6o4qy646  
         , u6xz15_qx1lay5yvg  
         , xj0hdx62yzgvd1qvsf  
         , tv1vy00negaq6kq  
         } = ysoarmlp98243p;

  
  wire dzkf25h87vtefb5g9p;

  ux607_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(hxhz0y3mpud0ey59v)
  ) y6y1rolk1b3j2ohl (
   .i_vld(mkvubuawtidmr0qz),
   .i_rdy(had01mmuqyc8tzrxd5), 
   .i_dat(ukllsj0e1xzeouqnrx),
   .o_vld(c_0qdn252ww1o9nhj4m), 
   .o_rdy(dzkf25h87vtefb5g9p), 
   .o_dat(ysoarmlp98243p),
 
   .clk  (gf33atgy  ),
   .rst_n(ru_wi)  
  );





  
  

  wire xvnxfgnlx05 = apnns9jlj7y3y5bg8ynz[21];
  wire h6yap55ubdbc2 = jv8kv41vzuir6an4iod[21];
  
  wire [5-1:0]      m603xpg5m7bwf6h1d    = dm_t8xh6s80cssm[4:0];
  wire [27-1:0]   nf7a14kdh46q_gb4d27t5o = dm_t8xh6s80cssm[(32-1):5];
  wire [6-1:0]      pkmbkt_zq0yhlemrgi = nf7a14kdh46q_gb4d27t5o[6-1:0];
  wire [21-1:0]        jcbv86t6ccbny9um2sm = nf7a14kdh46q_gb4d27t5o[27-1:6];

  wire apmzaxtau_e4j8y = xvnxfgnlx05 & (jcbv86t6ccbny9um2sm == apnns9jlj7y3y5bg8ynz[21-1:0]);
  wire mrwckdg2xmt_g4e = h6yap55ubdbc2 & (jcbv86t6ccbny9um2sm == jv8kv41vzuir6an4iod[21-1:0]);

  wire cavuvvu8tl9kpn5jta = (~( w1uq15jgugrn3 |  go95at_xv3zz734) & (~ z7yrukhpu2yv7));
  wire turhtksc36s_r8o3 = (~(a7hxr7wh300y3 | dqpjx6e7kt6x2csta) & (~lwq70xytakc30w));
  wire l3829ekia2rl6my8 = (~(g5dm3flv9 | y2yeehopezll49cmf) & (~bqbd1vx7u6p));
  wire xk5o0w8ij4dve8cxrwd22e = (~(n29ai3bkicr4tgyzgk | epi1zu1tfkun1al0l9) & (~etwu6izome4p5cwa0gn));

  wire b293miy3ig80jz = c_0qdn252ww1o9nhj4m & turhtksc36s_r8o3 & apmzaxtau_e4j8y;
  wire yz14ncxfv0 = c_0qdn252ww1o9nhj4m & turhtksc36s_r8o3 & mrwckdg2xmt_g4e;
  



  
 
 
  wire spb80jyq7y69vuz5xkn42;
  wire qregaax7ocnstzw2ho1oqtxfkfe;
  wire moz9tdl4bhiltwpdv96jd;
  wire [8-1:0]  jdklddtcs_yto5;

  wire zweqe8jmwo__bow5j94v68;
  wire s4ivomfr9adc7ty8xl_j;

  wire w9263gaw_lwsqx3wa;
  wire rg73_7zcjcm8e4w403bq;
  wire tgjvwosyypk2bxmb94;

  generate 
    if(64 == 64) begin:fjcbdq
        assign jdklddtcs_yto5 =
                                    (gstkdmb4wbsp8xhi == 2'b00) ? (8'b1 << dm_t8xh6s80cssm[2:0]) : 
                                    (gstkdmb4wbsp8xhi == 2'b01) ? (8'b11 << {dm_t8xh6s80cssm[2:1],1'b0}) : 
                                    (gstkdmb4wbsp8xhi == 2'b10) ? (8'b1111 << {dm_t8xh6s80cssm[2],2'b0}) : 
                                             8'b1111_1111; 
    end
    if(64 == 32) begin:g2z3f
        assign jdklddtcs_yto5 =
                                    (gstkdmb4wbsp8xhi == 2'b00) ? (8'b1 << dm_t8xh6s80cssm[1:0]) : 
                                    (gstkdmb4wbsp8xhi == 2'b01) ? (8'b11 << {dm_t8xh6s80cssm[1],1'b0}) : 
                                             8'b1111; 
    end
  endgenerate

  wire es9c9ezpnvof2_z9nmu;

  wire tmyzm9l_q256dqsxus = (dm_t8xh6s80cssm[32-1:3] == pq05yc_ea9cb[32-1:3]);
  wire unlfnqp2p2q8sa1 = ((jdklddtcs_yto5 & kogy6rrqymszp) == jdklddtcs_yto5);  
  assign tgjvwosyypk2bxmb94  = (~es9c9ezpnvof2_z9nmu) & turhtksc36s_r8o3 & brfek3hm0m1h_0qdx & x0pxzzrure0tp8zh3 & cik9g8nrdjspswqucoa9 & tmyzm9l_q256dqsxus & unlfnqp2p2q8sa1;
  assign rg73_7zcjcm8e4w403bq = (~es9c9ezpnvof2_z9nmu) & turhtksc36s_r8o3 & brfek3hm0m1h_0qdx & x0pxzzrure0tp8zh3 & cik9g8nrdjspswqucoa9 & tmyzm9l_q256dqsxus & (~unlfnqp2p2q8sa1);
  assign w9263gaw_lwsqx3wa  = (~es9c9ezpnvof2_z9nmu) & turhtksc36s_r8o3 & l3829ekia2rl6my8 & x0pxzzrure0tp8zh3 &  
                       (dm_t8xh6s80cssm[32-1:5] == pq05yc_ea9cb[32-1:5]);


 
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  

  wire vldo6rbn;
  wire tlwo81ky1a6b8;
  wire stol5aq_afcmhppp3t;
  wire vajnopldt37ec4kurfj9k;
  wire c8g86vay7y4o8r2d2hoh2e;
  wire jmc66mi6bkws1lwkk6krsjq;
  wire r9hqd030vnyga7o350en;
  wire l9x1ubg9wznb6ixv1i;
  wire kg739ybcd5xc49l6ph;
  wire iilu6o9khdb6tbh;

  wire zj05endwbrothpd7lkjs2qhspzr;
  wire rnlnwebfnqcg8g5oq_2gv0;
  wire y5otpn351odm3mnpnfdshm;
  assign es9c9ezpnvof2_z9nmu = stol5aq_afcmhppp3t;

  wire ero208rbddma5nko = (~(gxctvntt6usn533wgnh6 
                              & ((~rx250nlkrd2m3gkhtzzl) | (~x0pxzzrure0tp8zh3))
                              )
                              ) & (
  
                        (qregaax7ocnstzw2ho1oqtxfkfe) |
                        ( turhtksc36s_r8o3 & vldo6rbn & (
                                               moz9tdl4bhiltwpdv96jd   
                                             | w9263gaw_lwsqx3wa
                                                        )
                        ) |
                        ( turhtksc36s_r8o3 & (
                                             rg73_7zcjcm8e4w403bq |
                                             s4ivomfr9adc7ty8xl_j
                                              )
                        ) |
                       (vajnopldt37ec4kurfj9k ? 
                                    l9x1ubg9wznb6ixv1i : 
                                    (~rnlnwebfnqcg8g5oq_2gv0)
                       ) | 
                       (jmc66mi6bkws1lwkk6krsjq & 
                               kg739ybcd5xc49l6ph    
                       )
                       );

  
  
  
  
  

        
           
           

  wire hy9dltjwgw06uaq8h819ihk = (~xk5o0w8ij4dve8cxrwd22e) | (v_9kfy4x1fk3adyoz6x2);

  wire st7pytysu10a;
  wire mh9ba4wb9dl;
  wire j595qkrfu_okzcv0_4jxww_y_d;
  wire n0ilrfb6r31qw9dkf3mtds9;  
  wire hr3nk64lh9xbbegd9tyynan = 
                   
                       
                    n0ilrfb6r31qw9dkf3mtds9   
                       
                    | iilu6o9khdb6tbh  
                       
                    | j595qkrfu_okzcv0_4jxww_y_d   
                       
                    | tlwo81ky1a6b8  
                       
                    | (
                        hy9dltjwgw06uaq8h819ihk ? 
                                    tlwo81ky1a6b8 : 
                                    (~y5otpn351odm3mnpnfdshm)    
                      )
                    | (st7pytysu10a & gxctvntt6usn533wgnh6)
                    | (mh9ba4wb9dl & rx250nlkrd2m3gkhtzzl)
                    ;

  
  
  
  
  
  
  
  
  wire [64-1:0] zbzcbmwi85_njmfaks63ip;

  wire fxuirt21_3y5v;
  wire zwwbclwkk1c;
      
  wire   gdc31z_ah0g = (b293miy3ig80jz | yz14ncxfv0);
  wire   fknueo = (fxuirt21_3y5v | zwwbclwkk1c);
  assign vldo6rbn = ~gdc31z_ah0g;
  wire   cy0n2ao5wkp = ~fknueo;

  wire r7hgx17o2vo0lp = (
                         tgjvwosyypk2bxmb94 | 
                         zweqe8jmwo__bow5j94v68);
  wire [64-1:0] v_9rsloay1nw9k0k06 = 
                                     tgjvwosyypk2bxmb94 ? rxps0kbgar3hf :  
                                     zbzcbmwi85_njmfaks63ip ; 
  
     

  
  

  localparam l5_clmo2danmz_c19 = (hxhz0y3mpud0ey59v-4 +6 + 64 + 4*32 + 2*24 
                              );

  wire [l5_clmo2danmz_c19-1:0] e9v08zjfihbyxqc0;

  wire [24-1:0] ffb612_2t23r15a6tdgw;
  wire [24-1:0] gx97eig01em1bszuh7we;
  wire [32-1:0] xs8qjjjlfeb8dmez;
  wire [32-1:0] p7r5o9d5_pp1px2c7q;
  wire [32-1:0] b98ju_k45m18z96n0;
  wire [32-1:0] t9ilvhroqjh73dp7txy;

  wire [64-1:0] nnvljks2vlz8;
  wire [64-1:0] w6pgqo55vkzee_4;

  assign nnvljks2vlz8[31:00] = (~pq05yc_ea9cb[3]) ? xs8qjjjlfeb8dmez[31:00] : b98ju_k45m18z96n0[31:00];
  assign nnvljks2vlz8[63:32] = (~pq05yc_ea9cb[3]) ? p7r5o9d5_pp1px2c7q[31:00] : t9ilvhroqjh73dp7txy[31:00];
  assign w6pgqo55vkzee_4[31:00] = (~pq05yc_ea9cb[3]) ? b98ju_k45m18z96n0[31:00] : xs8qjjjlfeb8dmez[31:00];
  assign w6pgqo55vkzee_4[63:32] = (~pq05yc_ea9cb[3]) ? t9ilvhroqjh73dp7txy[31:00] : p7r5o9d5_pp1px2c7q[31:00];

  wire [l5_clmo2danmz_c19-1:0] twu59t94ybyqumq;
  wire teay27atwh1z5v;
  wire [64-1:0] mlnxnudr_2bo818byln;
  wire zklaicjqh98erk8;
  wire dmufi1xaijtfivbu;
  wire twgpc5472_utlu2og7;
  wire jzi3mgmyqego7mgsv81n;
  wire scx29q4wbo88sedwq;
  wire xa6a0counpp0ws7rema;

  wire yoa9z4x73xsc = xvnxfgnlx05 & apnns9jlj7y3y5bg8ynz[22];
  wire x4_cn1tzca1_ne = h6yap55ubdbc2 & jv8kv41vzuir6an4iod[22];
  wire smqoz2oj8ww5don  = xvnxfgnlx05 & apnns9jlj7y3y5bg8ynz[23];
  wire dh_clbn0o20fgf4  = h6yap55ubdbc2 & jv8kv41vzuir6an4iod[23];

  wire afvn9hlpbrsvtyljf6dx = xj0hdx62yzgvd1qvsf ? u6xz15_qx1lay5yvg : yz14ncxfv0;

  wire yng48_s157itc19pk504 = xj0hdx62yzgvd1qvsf ? 
                         (u6xz15_qx1lay5yvg ? h6yap55ubdbc2 : xvnxfgnlx05) 
                         : gdc31z_ah0g 
                         ;

  wire tdx3xfjrbjmmps2ga8p9 = ((yz14ncxfv0 & dh_clbn0o20fgf4) | (b293miy3ig80jz & smqoz2oj8ww5don));

  wire h46ue9w464mbm8tytu2nww = xj0hdx62yzgvd1qvsf ? 
                           (u6xz15_qx1lay5yvg ? (h6yap55ubdbc2 & x4_cn1tzca1_ne) : (xvnxfgnlx05 & yoa9z4x73xsc)) 
                         : ((yz14ncxfv0 & x4_cn1tzca1_ne) | (b293miy3ig80jz & yoa9z4x73xsc))
                         ;

  wire [21-1:0] felvo56_lohlxdcjbu91u = 
                     (u6xz15_qx1lay5yvg ? jv8kv41vzuir6an4iod[21-1:0] : apnns9jlj7y3y5bg8ynz[21-1:0]); 

  assign fzebl49irts00yi4k6c = {
                           ((rnj3s81yxus08gthgj & xj0hdx62yzgvd1qvsf) ? felvo56_lohlxdcjbu91u : jcbv86t6ccbny9um2sm),
                           pkmbkt_zq0yhlemrgi,
                           m603xpg5m7bwf6h1d
                           };  

  
  wire xe1me4zn_lzcyrxb7l = (rnj3s81yxus08gthgj & ie6x4201u8jyqlgs) ? h46ue9w464mbm8tytu2nww : 1'b0;
  
  wire og1dtdfkkbx1ybmy60 = (rnj3s81yxus08gthgj & auhnvtbztby6o4qy646) ? yng48_s157itc19pk504 : 1'b0;



  wire b6zx6289bg21bxi1h4 = ((rnj3s81yxus08gthgj & ie6x4201u8jyqlgs) & h46ue9w464mbm8tytu2nww) 
                          | ((rnj3s81yxus08gthgj & auhnvtbztby6o4qy646) & yng48_s157itc19pk504);

                          
                          
                          
                          
                          
                          
                          
                          
                          
  wire iemcihl0h3gjp = (smqoz2oj8ww5don | dh_clbn0o20fgf4);

  wire wwjqqdj9evzwv7l5b4erq = 
                        
                 gdc31z_ah0g ? ((~tdx3xfjrbjmmps2ga8p9) & iemcihl0h3gjp) : 
                        
                     iemcihl0h3gjp;

  wire vvjh1x6zug_z3vtoji = wwjqqdj9evzwv7l5b4erq | tdx3xfjrbjmmps2ga8p9;
  wire jhpjh6z62fydj9djbf = ~tdx3xfjrbjmmps2ga8p9;
  wire qlu1lged673hkbvh8vh = (rnj3s81yxus08gthgj & (~qu2oxvm9fx85hbf) & (~fyqztmgm7gm2uol7)) ? (~b6zx6289bg21bxi1h4) : 1'b0;
  wire u4l3r6vwoso0zb2tchavbx1_g   = (rnj3s81yxus08gthgj & qu2oxvm9fx85hbf) ?  vvjh1x6zug_z3vtoji : (rnj3s81yxus08gthgj & fyqztmgm7gm2uol7) ? jhpjh6z62fydj9djbf : 1'b0;
  wire wbj6b4bflmlwk6olgu   = xa74n2vq7asiuic23w ? 1'b1 : 1'b0;
  wire e3ldjb4w8w0e = qlu1lged673hkbvh8vh | wbj6b4bflmlwk6olgu | u4l3r6vwoso0zb2tchavbx1_g;

                            
  wire mfc7n7sv4xkc6v10a = yqc55f6txw_pmexi & (jzi3mgmyqego7mgsv81n | scx29q4wbo88sedwq) & fknueo;


  assign e9v08zjfihbyxqc0 = {
                                           apnns9jlj7y3y5bg8ynz 
                                         , jv8kv41vzuir6an4iod 
                                         , tkt93y5lfluzkia5plvksp 
                                         , g4nfgu53_rgc0632w8z97 
                                         , ql1c7hzoj9kf__7r97krm 
                                         , ryid4_99ns1jc83at_88x 
                                         , r7hgx17o2vo0lp
                                         , v_9rsloay1nw9k0k06
                                         , ero208rbddma5nko
                                         , b293miy3ig80jz
                                         , yz14ncxfv0
                                         , kggnqtwc1ljww3tnze 
                                         , mih7nmwcak45d8a2hvfx 
                                         , z_c9c063dzhr5i2tflx1ge 
                                         , gxctvntt6usn533wgnh6  
                                         , xe1me4zn_lzcyrxb7l
                                         , vfzxxuugm86jff_8iod
                                         , og1dtdfkkbx1ybmy60
                                         , qu2oxvm9fx85hbf
                                         , fyqztmgm7gm2uol7
                                         , afvn9hlpbrsvtyljf6dx
                                         , ts27sjuboaf8qsmg  
                     };


  assign {
                                           ffb612_2t23r15a6tdgw 
                                         , gx97eig01em1bszuh7we 
                                         , xs8qjjjlfeb8dmez 
                                         , p7r5o9d5_pp1px2c7q 
                                         , b98ju_k45m18z96n0 
                                         , t9ilvhroqjh73dp7txy 
                                         , teay27atwh1z5v
                                         , mlnxnudr_2bo818byln
                                         , stol5aq_afcmhppp3t
                                         , fxuirt21_3y5v
                                         , zwwbclwkk1c
                                         , tftxelzlbcv3nmg0ry 
                                         , c7l7vyum1z06i355gent 
                                         , d42b0dgiiybnaa647lv9euj 
                                         , rx250nlkrd2m3gkhtzzl  
                                         , zklaicjqh98erk8
                                         , dmufi1xaijtfivbu
                                         , twgpc5472_utlu2og7
                                         , jzi3mgmyqego7mgsv81n
                                         , scx29q4wbo88sedwq
                                         , xa6a0counpp0ws7rema
                                         , gs05ko46ogh5  
                                                          } = twu59t94ybyqumq;

                     

  wire gcsfsfehlyi7d5tcd25;
  wire a86ti3q3r0b3s2a_evs;

  assign gcsfsfehlyi7d5tcd25 = (~e3ldjb4w8w0e) & c_0qdn252ww1o9nhj4m;
  assign dzkf25h87vtefb5g9p =   e3ldjb4w8w0e  | a86ti3q3r0b3s2a_evs;

  wire gq3w46enpc5p1ls = c_0qdn252ww1o9nhj4m & dzkf25h87vtefb5g9p;
  assign ytaw26fvd4q2bkrmzdzc20exc7nofso = gq3w46enpc5p1ls & (qlu1lged673hkbvh8vh | u4l3r6vwoso0zb2tchavbx1_g) ;
  wire fgru0fi7v178lp914d4zbdmqs63z_4 = gq3w46enpc5p1ls & u4l3r6vwoso0zb2tchavbx1_g;
  wire w6m1johuy8qk9wgea0xqv12l_tkgb = gq3w46enpc5p1ls & qlu1lged673hkbvh8vh;
  wire kngugv98d1yeo511y = wwjqqdj9evzwv7l5b4erq & rnj3s81yxus08gthgj & qu2oxvm9fx85hbf;

  wire uvper_b758sow8j9u;

  
  ux607_gnrl_pipe_stage # (
   .CUT_READY(0),
   .DP(1),
   .DW(l5_clmo2danmz_c19)
  ) ftse_79a41hd52 (
   .i_vld(gcsfsfehlyi7d5tcd25),
   .i_rdy(a86ti3q3r0b3s2a_evs), 
   .i_dat(e9v08zjfihbyxqc0),
   .o_vld(x0pxzzrure0tp8zh3), 
   .o_rdy(uvper_b758sow8j9u), 
   .o_dat(twu59t94ybyqumq),
 
   .clk  (gf33atgy  ),
   .rst_n(ru_wi)  
  );

  assign  bpmlbcph7uz4fmydd  = ( cavuvvu8tl9kpn5jta &    n15yjlq97s5vf9  & (~ wzpsauw3j_6xyp0));
  assign brfek3hm0m1h_0qdx  = (turhtksc36s_r8o3 &   io1dzzuksv6fh6w  & (~rnj3s81yxus08gthgj));
  assign t1cqzavxcqpcddy3yhtk  = (l3829ekia2rl6my8 &   jxbtey15c3kkb7  & (~yqc55f6txw_pmexi));
  assign pn0blb6qozvruaiaccluecd  = (xk5o0w8ij4dve8cxrwd22e &   hh6d0ibqo915gqaoole  & (~v_9kfy4x1fk3adyoz6x2));

  assign  dsrz57a4u1pediag = ( cavuvvu8tl9kpn5jta & (~ n15yjlq97s5vf9) & (~ wzpsauw3j_6xyp0));
  assign c5luf4ekdp8uxjd6phdb = (turhtksc36s_r8o3 & (~io1dzzuksv6fh6w) & (~rnj3s81yxus08gthgj));
  assign cik9g8nrdjspswqucoa9 = (l3829ekia2rl6my8 & (~jxbtey15c3kkb7) & (~yqc55f6txw_pmexi));
  assign w3o65s8zjg4wgjw69l7iz58u = (xk5o0w8ij4dve8cxrwd22e & (~hh6d0ibqo915gqaoole) & (~v_9kfy4x1fk3adyoz6x2));
  
  
  wire goqh7apc7a08bj9u = x0pxzzrure0tp8zh3 & uvper_b758sow8j9u;
  assign q6dwr6kors49 = goqh7apc7a08bj9u & (~d42b0dgiiybnaa647lv9euj);
 
  wire irwg_3zavoi9g_a;
  assign uvper_b758sow8j9u = d42b0dgiiybnaa647lv9euj ? 1'b1 : 
                            irwg_3zavoi9g_a;


  wire [64-1:0] vo0toaa76g8ksriet = 
                         (       ({64{fxuirt21_3y5v}} & nnvljks2vlz8) |
                                 ({64{zwwbclwkk1c}} & w6pgqo55vkzee_4)  
                 );

  wire [3-1:0] of351wfep15ud51 = 
                         (       ({3{fxuirt21_3y5v}} & ffb612_2t23r15a6tdgw[(24-1):21]) |
                                 ({3{zwwbclwkk1c}} & gx97eig01em1bszuh7we[(24-1):21])  
                 );

  wire  pt5n0kv5bpa59b31 = 1'b0;

  wire sh76lsmx = fxuirt21_3y5v | zwwbclwkk1c;
  wire rcd3m3rlm8xp = b293miy3ig80jz | yz14ncxfv0;

  wire o1_8jcyxk9tk = rcd3m3rlm8xp | r7hgx17o2vo0lp;
  wire bgt76tmzqwy1 = sh76lsmx | teay27atwh1z5v;
  wire [64-1:0] rark_9btzysdimqacli9_ = teay27atwh1z5v ? mlnxnudr_2bo818byln : vo0toaa76g8ksriet;
  wire f3gvutnvfx6bx6wg = teay27atwh1z5v ? 1'b0 : pt5n0kv5bpa59b31;


  
  assign st7pytysu10a = c_0qdn252ww1o9nhj4m & (~z_c9c063dzhr5i2tflx1ge);
  assign mh9ba4wb9dl = x0pxzzrure0tp8zh3 & (~d42b0dgiiybnaa647lv9euj);
  wire qgppmd2m94otu5uxqbc7hc = x0pxzzrure0tp8zh3 & d42b0dgiiybnaa647lv9euj;

  
  assign r9hqd030vnyga7o350en = (mh9ba4wb9dl & ((t1cqzavxcqpcddy3yhtk & bgt76tmzqwy1) | bqbd1vx7u6p ));
  wire pirp8rqhngzyt0i6     = r9hqd030vnyga7o350en & (~es9c9ezpnvof2_z9nmu); 

  
  assign zj05endwbrothpd7lkjs2qhspzr = (mh9ba4wb9dl & cik9g8nrdjspswqucoa9 & sh76lsmx & (~bqbd1vx7u6p));
  assign jmc66mi6bkws1lwkk6krsjq = (st7pytysu10a & c5luf4ekdp8uxjd6phdb & rcd3m3rlm8xp & (~lwq70xytakc30w));
  wire dayo38p_tlcb6n0ov6qg; 
  wire ud_fiihzz8uhok5wic8ha     = zj05endwbrothpd7lkjs2qhspzr & (~es9c9ezpnvof2_z9nmu);
  wire ecp10s0k_n91ef_jrkaki = q6dwr6kors49 & ud_fiihzz8uhok5wic8ha;

  
  
  
  
  
  assign vajnopldt37ec4kurfj9k = (st7pytysu10a & (~lwq70xytakc30w) & (
                  (brfek3hm0m1h_0qdx & (~o1_8jcyxk9tk)) 
                | (c5luf4ekdp8uxjd6phdb & (~rcd3m3rlm8xp)) 
                | (~turhtksc36s_r8o3) 
                | (rnj3s81yxus08gthgj) 
                )
            );
  assign c8g86vay7y4o8r2d2hoh2e = (mh9ba4wb9dl & (~bqbd1vx7u6p) & (
                  (t1cqzavxcqpcddy3yhtk & (~bgt76tmzqwy1)) 
                | (cik9g8nrdjspswqucoa9 & (~sh76lsmx)) 
                | (~l3829ekia2rl6my8) 
                | (yqc55f6txw_pmexi) 
                )
            );
  wire xn4ip9xr3j5q3rg2n4_8 = c8g86vay7y4o8r2d2hoh2e & (~es9c9ezpnvof2_z9nmu);

  wire qhwwiyjvan775z6uijmq83;

  assign vc0fhfx87dxbgty02yd = mh9ba4wb9dl & es9c9ezpnvof2_z9nmu;
  
    
    
    
    
 
 
 
  wire g_2b1ve9yzm7fl9pmmenkwrstu4882 = cik9g8nrdjspswqucoa9 & (
                             
                           sh76lsmx ? 1'b1 : 
                             
                                 
                           lv2obxi3r4ob ? 1'b0 : 
                                 
                               y5otpn351odm3mnpnfdshm 
                               );

  wire eqdfw7tfoezk75p7hrkkc = ( pirp8rqhngzyt0i6 | 
                         ((mh9ba4wb9dl & g_2b1ve9yzm7fl9pmmenkwrstu4882) & (~es9c9ezpnvof2_z9nmu))
                     );

  wire w0kqiyhky226say_7mo6b5s =
                   yqc55f6txw_pmexi 
                   
                 | g_2b1ve9yzm7fl9pmmenkwrstu4882
                 ;


  assign irwg_3zavoi9g_a = 
                                                     
                                                     
                                                     
                          (eqdfw7tfoezk75p7hrkkc ? dayo38p_tlcb6n0ov6qg : 1'b1)
                        ;




  wire                   r57mgw9ntmg26lxok;
  wire                   cac59gne730vqiq;
  wire                   ypuolenm4dvdg;
  wire                   yu5m552dobcb8gbsq;
  wire  [64-1:0] bo_q_t246zgg3q; 

  assign klkflmsyyf5w7ar = 
             eqdfw7tfoezk75p7hrkkc |

                     r57mgw9ntmg26lxok;

  wire [32-1:0] d4k4iwwrjuzjqt;
  wire [32-1:0] v7q8td8d2htgx9l =   
                           r57mgw9ntmg26lxok ?
                                          d4k4iwwrjuzjqt 
                                        : pq05yc_ea9cb 
                                        ;

  assign h7f6k_ims_9p3 =  
                           r57mgw9ntmg26lxok ?
                                          bo_q_t246zgg3q 
                                        : rark_9btzysdimqacli9_ 
                                        ;
  assign lkjqs6kiuyj   =  
                           r57mgw9ntmg26lxok ? 
                                          ypuolenm4dvdg 
                                        : f3gvutnvfx6bx6wg 
                                        ;
  assign u245it8jnyhc3eqcy0 =  
                           r57mgw9ntmg26lxok ? 
                                          yu5m552dobcb8gbsq 
                                        : 1'b0 
                                        ;


  assign cac59gne730vqiq = wy36iirxspfw56864;
  assign dayo38p_tlcb6n0ov6qg = r57mgw9ntmg26lxok ? 1'b0 : wy36iirxspfw56864;





  
  
  
  
  
  
  
  
  
  
  

  localparam n3bc49qfitvsyfxo = f16zrowg1s1f5 + 6;
  wire pzisij4j58gth_qfo;
  wire fkfwa26f8gf5283f;
  wire [n3bc49qfitvsyfxo-1:0] ss0c22d2fj3oh7;

  assign pzisij4j58gth_qfo = vc0fhfx87dxbgty02yd;
  wire [n3bc49qfitvsyfxo-1:0] nvd_v9290iorcv = {
                                           zklaicjqh98erk8
                                         , dmufi1xaijtfivbu
                                         , twgpc5472_utlu2og7
                                         , jzi3mgmyqego7mgsv81n
                                         , scx29q4wbo88sedwq
                                         , xa6a0counpp0ws7rema
                                         , gs05ko46ogh5
                                         };  

  assign {
                                           dbkpihmr6104_e36q4zoxpgy
                                         , gxv5oxyuuit9f6lci1p0v22
                                         , bfrlc8tog574i131socryaap
                                         , v5rjtrkyv236_aeycevjw
                                         , v14gd4036xa4fahc_461n
                                         , ti3tf23yq0i6r0hmenfl6
                                         , ky8zw277b8fa1dq1zk
                                         } = ss0c22d2fj3oh7;

  
  


  ux607_gnrl_fifo # (
   .CUT_READY(0),
   .DP(3),
   .DW(n3bc49qfitvsyfxo )
  ) jc3hg9nqm17a5u7vt4kbln1 (
   .i_vld(pzisij4j58gth_qfo),
   .i_rdy(fkfwa26f8gf5283f), 
   .i_dat(nvd_v9290iorcv),
   .o_vld(nvlcc2cq4xv0339t), 
   .o_rdy(d8fgkbjcpmd8_4r), 
   .o_dat(ss0c22d2fj3oh7),

   .clk  (gf33atgy  ),
   .rst_n(ru_wi)  
  );


  wire e8qfsi5gi5d6er2yq5s = pzisij4j58gth_qfo & fkfwa26f8gf5283f;
  wire m8vq9bker6sf_h1wgtana6 = ~nvlcc2cq4xv0339t;
     
  assign qregaax7ocnstzw2ho1oqtxfkfe = (~m8vq9bker6sf_h1wgtana6) | e8qfsi5gi5d6er2yq5s;
  assign spb80jyq7y69vuz5xkn42 = (~m8vq9bker6sf_h1wgtana6);

  
  assign hcjwu1jmlbr4k4wahdf0ju = (~hr3nk64lh9xbbegd9tyynan) & nvlcc2cq4xv0339t;
  assign d8fgkbjcpmd8_4r       = (~hr3nk64lh9xbbegd9tyynan) & k71jdwvt1q_yy5a7kzwp8cz;
  


 
  
  
  
  
  
  
  
  
  
  
  


  
  wire oyfo3haj43lmbk8ds = ecp10s0k_n91ef_jrkaki & (~qhwwiyjvan775z6uijmq83);
  wire vhbxz8svsbljbu;
  wire rkx4pzzf1tu01m4j;
  
  
  

  localparam jkw_w4sdw6oadn = (1 +3 +32+64+8);

  wire [jkw_w4sdw6oadn-1:0] r092q73gt_7atlt1a;
  wire [jkw_w4sdw6oadn-1:0] gijtnhz7eo3v_;

  assign r092q73gt_7atlt1a = {
                                           fxuirt21_3y5v
                                         , of351wfep15ud51   
                                         , pq05yc_ea9cb
                                         , rxps0kbgar3hf [64-1:0]
                                         , kogy6rrqymszp [8-1:0]
                     };


  assign {
                                           y4z10x_uk5tx9gjpp
                                         , vt4fxo524ecd4y832detyma   
                                         , cb39rlyxl60nbkm
                                         , c3h8wzh_yyz3847v [64-1:0]
                                         , zz8qhy80jaf147ase [8-1:0]
                                         } = gijtnhz7eo3v_;



  yjm16kn_qwdkfm8if #(
      .xl24j_imhfhfk(jkw_w4sdw6oadn)
)y4i2i8s804fbrib95dab (
   .stbblp081kc9    (oyfo3haj43lmbk8ds),
   .vulpj3pebksw    (vhbxz8svsbljbu), 
   .wbo1zx8iepki     (r092q73gt_7atlt1a),
   .z4qzurty_axomdd    (j55vt_3172gxi8el), 
   .clwlpmx87nqbuq    (rkx4pzzf1tu01m4j), 
   .atl5amsp8tyrm     (gijtnhz7eo3v_),

   .j8kotg18hji        (brfek3hm0m1h_0qdx),
   .gebnakb8ctgri6s   (dm_t8xh6s80cssm),
   .rfdekem29gp7jx0f1   (gstkdmb4wbsp8xhi),
   .krasg_k9_i1zsgbu   (s4ivomfr9adc7ty8xl_j),
   .sf5oaemd1e3k    (zweqe8jmwo__bow5j94v68),
   .ycj5xet5wunw0c  (zbzcbmwi85_njmfaks63ip),

   .pf8rzr1mv        (pn0blb6qozvruaiaccluecd),
   .rj1cfvu3meww   (fwgc_k58kjyp_va),
   .s2fbnn6ekvrsa3j   (xkopv4_km4ey9cihevo2),
   .g_w2g5ygcfsk   (n0ilrfb6r31qw9dkf3mtds9),
   .k4olvo5ol6hvag    (),
   .oivxcjfrvf9efavm  (),

   .x6n2fwiz0cogynnbie (ecp10s0k_n91ef_jrkaki),
   .ncetuvy4lmo       (cik9g8nrdjspswqucoa9),
   .diat9bfkf7mnu  (pq05yc_ea9cb),
   .dn53sr7lydjdo5 (rxps0kbgar3hf),
   .hc79i6u2twxms6ke (kogy6rrqymszp),
   .ybztfzzlexmx9gk   (qhwwiyjvan775z6uijmq83),

   .ahth5hydygfua1j2   (kg739ybcd5xc49l6ph),

   .gf33atgy  (gf33atgy  ),
   .ru_wi(ru_wi)  
  );

  
  assign f1xe_xx4j29e7277py1p2k9uh = (~qhwwiyjvan775z6uijmq83) & j55vt_3172gxi8el;
  assign rkx4pzzf1tu01m4j       = (~qhwwiyjvan775z6uijmq83) & te46hx1x_954f8oaiw8vpfl7;
  

  assign iilu6o9khdb6tbh  = ~vhbxz8svsbljbu;

  assign lgdhsk7cwbxgrv43 = j55vt_3172gxi8el & rkx4pzzf1tu01m4j;














  wire                          g3_8p4g7w5grnl62xy;
  wire                          vqwqaofc8sz_yjccd;


  wire                          tyxs3jzhr2i2gq9dt7 = qgppmd2m94otu5uxqbc7hc;
  wire                          zti98n829owa2p;

  wire [24-1:0]   ye256knohacnaakiw2nqck6 = ffb612_2t23r15a6tdgw;
  wire [24-1:0]   hyxeikuobvxjumz2hibay = gx97eig01em1bszuh7we;
  wire [32-1:0]  zkojor8433oflab2kpvtzi1z9 = xs8qjjjlfeb8dmez;
  wire [32-1:0]  nx6i4o0_cbqmlan1ylpodj9y = p7r5o9d5_pp1px2c7q;
  wire [32-1:0]  tgfv2w2s7qhwkl0pdpf_79v4e = b98ju_k45m18z96n0;
  wire [32-1:0]  qfjl6250hpfb57pxl0t53q6fd = t9ilvhroqjh73dp7txy;

  wire cgnsvvj7srbljqst;
     

  wire [6-1:0]      li2o0fhy6bmhmqeoi6rm;

  assign jgeyki3wp7rzhsh958 = mh9ba4wb9dl & mfc7n7sv4xkc6v10a;
  wire tr_rxyj9lr38m35v2 = xn4ip9xr3j5q3rg2n4_8 & q6dwr6kors49 & mfc7n7sv4xkc6v10a;
  wire vvhwrir0m93lfnd   = xn4ip9xr3j5q3rg2n4_8 & q6dwr6kors49 & (~mfc7n7sv4xkc6v10a);

  assign nsc0elm1w3m_inebi5nie51   = tr_rxyj9lr38m35v2 & fxuirt21_3y5v;  
  assign kbae6svksx713v4pbhv8   = tr_rxyj9lr38m35v2 & zwwbclwkk1c;  
  assign hgfb_gwm97sz53betsjyk5 = li2o0fhy6bmhmqeoi6rm;
  assign ee18h0eqehcvi043ns32gf = li2o0fhy6bmhmqeoi6rm;
  assign qxdc_js0dtaug304lp11_gu   = 1'b1;
  assign tarnkvmavl9287x895   = 1'b1;
  assign bshid8lzm3x5d3ju1u82v  = (((24'b100<<21) & {24{jzi3mgmyqego7mgsv81n}}) | ((~(24'b100<<21)) & ffb612_2t23r15a6tdgw));
  assign wuf4wr1vape2nd15r20p  = (((24'b100<<21) & {24{jzi3mgmyqego7mgsv81n}}) | ((~(24'b100<<21)) & gx97eig01em1bszuh7we));
 


  wire tq5w2fd0flcywep677l;
  wire juwj_oo3r8yt2a4hg;
  wire k6_e3_saw0oup16pudov;
  wire pzfb_24lrjd770iigjx4sm;
  wire [6-1:0] zpq6nysk8b654ynyt4zj9k;
  wire [6-1:0] d2lstp52x9w9900ioarrtfk;


  wire a03er8qo6p0zpb           ;
  wire bzsjo5unerpy5i0e_q_6eqn    ;
  wire z8uuyp_3l6aqut86nkd__vvwgs    ;
  wire ctfhepdgvm53k59kbbe0s0924he0ijd;


  gsmnxrg40o2b1e4gc d6k03s8r61oq7p(


    .hv39pppvbmeqy8b6       (hv39pppvbmeqy8b6       ),
    .t6l88yqbe4wokkhiso9t      (t6l88yqbe4wokkhiso9t      ),
    .hyec__ebnw8lbcssd81      (hyec__ebnw8lbcssd81      ),
    .vs2610q9_on1r996p     (vs2610q9_on1r996p     ),
    .coy3buxdw6yq3duh21azuwflk(coy3buxdw6yq3duh21azuwflk),
    .r_8h5lxb39ug57zli04e_o     (r_8h5lxb39ug57zli04e_o     ),
    .pv7q0ikpayogkay57rgyr     (pv7q0ikpayogkay57rgyr     ),
    .dsq8f3rhmb7yc876v8    (dsq8f3rhmb7yc876v8    ),
    .enu_vumk17eoj1fma5ilz0   (enu_vumk17eoj1fma5ilz0  ),
                                                  
    .ou74jmm5p6th0y0kcdwpqv2ey(ou74jmm5p6th0y0kcdwpqv2ey),
    .adwzzx09c_s_x1seh     (adwzzx09c_s_x1seh     ),
    .zp0aylmm0k4yw4w561bgzh   (zp0aylmm0k4yw4w561bgzh   ),


    .a03er8qo6p0zpb              (a03er8qo6p0zpb           ),
    .bzsjo5unerpy5i0e_q_6eqn       (bzsjo5unerpy5i0e_q_6eqn    ),
    .z8uuyp_3l6aqut86nkd__vvwgs       (z8uuyp_3l6aqut86nkd__vvwgs    ),
    .ctfhepdgvm53k59kbbe0s0924he0ijd(ctfhepdgvm53k59kbbe0s0924he0ijd),

    .tq5w2fd0flcywep677l  (tq5w2fd0flcywep677l  ),
    .juwj_oo3r8yt2a4hg  (juwj_oo3r8yt2a4hg  ),
    .k6_e3_saw0oup16pudov (k6_e3_saw0oup16pudov ),
    .pzfb_24lrjd770iigjx4sm (pzfb_24lrjd770iigjx4sm ),
    .zpq6nysk8b654ynyt4zj9k(zpq6nysk8b654ynyt4zj9k),
    .d2lstp52x9w9900ioarrtfk(d2lstp52x9w9900ioarrtfk),

    .sej7ti3911672ok72k    (vvhwrir0m93lfnd  ),
    .z2s7c4x2upx2k94    (),

    .kix9_o92mst68vescu79v (w0kqiyhky226say_7mo6b5s),
    .hdwldkfk3vetnqg3us     (pq05yc_ea9cb    ),
    .ihkz9tebg3jd5f47z    (io1o8wz_hhx_efhn   ),
    .tu1v8ryo2rv95crsvz    (ar75eg689jsahd   ),
    .ghikvq604upn2v    (lv2obxi3r4ob   ),
    .oodqv7hv99boddj3kk48j    (ntwmchaa8jnutooi3_   ),
    .t4leke6w3uzo3gxu3yhk    (l3i_yp_t5k_ghmdbmvrk4   ),
    .g2x5gi27ly4aw24   (y2yeehopezll49cmf  ),
    .g16len3w2wk22u       (g5dm3flv9      ),
    .vx_fynrmojs7gx     (jxbtey15c3kkb7    ),
    .xpd4oma8mrw21r9b0mc8c (t1cqzavxcqpcddy3yhtk ), 
    .ytx0p13ahjuk751e8crl_0(cik9g8nrdjspswqucoa9), 
    .uacpumgrbwt0fmb    (rxps0kbgar3hf   ),
    .v0uq3fcdfb8eatt3    (kogy6rrqymszp   ),
    .c4otadutq6rav14ed2     (hqchs835s6qbo2wr    ), 
    .mw8uaelv0i5zfav     (kfjijv_31s3    ), 
    .uq0oocqz_ys0no4o_t     (g6qm6ye0l65m    ),
    .ohprpkw231g_f2qqzmq (yqc55f6txw_pmexi),
    .e3l8n6__k56uw5o7jujwibr (zklaicjqh98erk8),
    .rwmac6nity_ikz7xbj_ta1nce  (dmufi1xaijtfivbu ),
    .en9ogfq6nx_uirma3y2jiigbh (twgpc5472_utlu2og7),
    .t9otq6y33fc5qs21p9d2rc3zn (jzi3mgmyqego7mgsv81n),
    .xpbzeko14yty79dehft9e2l (xa6a0counpp0ws7rema),

    .r57mgw9ntmg26lxok    (r57mgw9ntmg26lxok   ),
    .cac59gne730vqiq    (cac59gne730vqiq   ),
    .ypuolenm4dvdg      (ypuolenm4dvdg     ),
    .yu5m552dobcb8gbsq  (yu5m552dobcb8gbsq ),
    .bo_q_t246zgg3q    (bo_q_t246zgg3q   ), 
    .d4k4iwwrjuzjqt     (d4k4iwwrjuzjqt    ), 

    .ktkt_7t0wo1gkg8gormhm    (cv0k9k_ijjnnylw1s7b_0d    ),

    .rjy1ysvx9590bpklijsn0ucgaga  (swpk4h0gei3t_34xogbqncbo4  ),
    .d_933icutbtk8nknxip5t1ds  (u9qmfl3rwx0dhr92z875vx7q  ),
    .a45qubts5uovcopirpl9jxs7uia   (unu_x_i6jmr33nz0yitzk   ),
    .kwbu6olmnnt53fot6kfntm2q7t   (bei3qhdtd0euq2emblogsu_x   ),
    .kq9lkjt85jst7fa5smg1nud  (bf0_ynb648lqi7s93eieo0ln  ),
    .mekhipn8vmxn5adno3jrpek8nkm  (wf8o7p9_qfthhoxs747wyeuwkky  ),
    .wbwviedmyjzfiwi2t1yh0ibf7wv3  (ygro7xue7x7rtdafkj3o4q4  ),
    .h99v8xeu9gkycpsn1wl3lrow7   (drrly3q0ocg8d4pwh3m9o77   ),
    .jvloelo3plm6zwbisesi7fwa   (g654a6a9cesbee7xs6_uu9lu5   ),
    .ecz8u30wtuyonhyfwfrfrc30g   (x7fex0jf9da6a5v1c28upl72t   ),
    .vxwea8jbxv6m5tu7nkqtf6   (ege0_1ufqm8i68zo4il6cwe46d   ),
    .jsswxoezxjsdw154f5xt1omqrup  (ngyxf4n1cpcgks_s2zmgfb260  ),
    .e5cyxxxkg4061gq3_ksqdax_7op  (c7m50uaw8lmp_iv4ci38q2  ),
    .m3pduyvpfh4ximuy0dl6k_wjuc  (m04a1mtbabwezldp1crh4rg6z  ),
    .xhts19tgn12c186fduss6cfjyz (hwjq1ubtaei44lpk609fm2hb8 ),
    .zt7xddfgq3m2nsc8s_3a48r8     (e28p_fu1k484ncul0p85ko     ),

    .s9lcmqjp282zoimy_nw6kv2u    (a0_d_zdz9h9fgk46e8arf    ),

    .pkm6vgcr8iz_el5103gzwdew0hki  (twr9y24wxhs3qj2z9f2hzpaig6  ),
    .vdbkch1krpijvuukam8k5_9g6h4d  (w8b46r9cof57xvd5zo1u4zh8  ),
    .gi8g2jgc5r69ozgg2517f4   (wn1l4cmih7rwce1rb7wk3f9wy   ),
    .nqq4y60r7eh5lbir_nzlqf2q7k   (cgnzbuo_1yz6v42seb25duv   ),
    .rf_rtoowzj9m6zi6taqyqn6ku  (zopev7f487spn9mwvuowqo  ),
    .kqa4ro7t84z342uqr2plzmi1  (p32jk0lb8g31kqlpvmllo75qim  ),
    .d50l6nnxdfj7iuhnqe9gjobewaj4  (g973rcaou05i456suvk_89dm  ),
    .ziqf65e93q9kc_6bj_n4gd2op   (wflv6rhfdwyxttak111v1l   ),
    .lkflakila483fdjdz1hrtobjiz   (ggsmt4nzx8pwlowehinqvk60f   ),
    .zg0qkr8fhe1v0eku3at17q   (xu8494ii8ectqb91224uuer   ),
    .gu2ufdscjjb3hvpwrwu6c8h   (r6rk128ijo839ougen9stbe   ),
    .pn9rf9nl21n4t8clpsygzbo72n  (xo6ciibewn8p8xey97jcsqi5  ),
    .u6t2h_hm580phvwuvdedyagaqg  (evz1w_girwszyfnlcg4mwvtjo  ),
    .h1p8zhyrvirdo9c78wx8cmal83  (ju5f9fb1erjep_bv8gpfn6  ),
    .d11v3v5k967aul6l7_up53azs (hadi1_f3quoaotjv5758x8kksot2 ),
    .tnfd_mhtdr0hw58lveup8w8     (bdi4gjlb0po4ejcztowoqil7     ),

    .fp_qm6eq7380_uydc6pb2sw7  (bvg_3t_ujbpur7b_h7f63jse  ),
    .z9eviza6dmjc6u7jbuzirzh8z1ce  (m5l6wu3uz_jfqasz8e3tsvrm  ),
    .gz2qngl9towiwc_nk48gu38p9    (g9so28ythfl0q7xnk66p1    ),
    .saolr4xnpfm570snrsqk7hazshkz(e66wluxk71p2ldu3a1qk994bq),
    .b85cqul2sjbg0c5ta0bcpgpluvma  (ig2roj0y08x8_ntp3knz9rd  ),

    .me8sa0hl_2m6xmtdm4r_1tn7cer4  (m7tq_t57mr5bovbb9ghffl4k  ),
    .gv_wy8qy9rm50mn4yg66yvagb60l  (gpcgdcri3e6_fxrw8wwtysoqqr  ),
    .byn2o0bi_9ggzegrnvskn    (a6s4kxg1ibr6mntc85jik    ),
    .m12x1nn4kvsdeqofo9rqi8aawa(hizzalmpwr8cqkxqi80wvbt65x),
    .e0xiuuzhk1qbwdjlub9o_cca5  ({64{1'b0}}),

    .jkq984ky8fozrzq             (jkq984ky8fozrzq           ),
    .g3_8p4g7w5grnl62xy          (g3_8p4g7w5grnl62xy        ),
    .vqwqaofc8sz_yjccd          (vqwqaofc8sz_yjccd        ),
    .tyxs3jzhr2i2gq9dt7          (tyxs3jzhr2i2gq9dt7        ),
    .zti98n829owa2p          (zti98n829owa2p        ),
    .ye256knohacnaakiw2nqck6   (ye256knohacnaakiw2nqck6 ),
    .hyxeikuobvxjumz2hibay   (hyxeikuobvxjumz2hibay ),
    .zkojor8433oflab2kpvtzi1z9   (zkojor8433oflab2kpvtzi1z9 ),
    .nx6i4o0_cbqmlan1ylpodj9y   (nx6i4o0_cbqmlan1ylpodj9y ),
    .tgfv2w2s7qhwkl0pdpf_79v4e   (tgfv2w2s7qhwkl0pdpf_79v4e ),
    .qfjl6250hpfb57pxl0t53q6fd   (qfjl6250hpfb57pxl0t53q6fd ),
     
    .j2kcz1faqhvh1ler6j       (e3rxl7mic_dpejl98_ts2  ),
    .a6gdkt5h77dh0mcj8t4gq     (dlxukfkm1k19y_gskjb9vnl),
    .wixbtbeqlhzelg4t       (sdmu0iskkbwi6blvi5  ),
    .uh_ekyw7cw8c3d3xj1      (suwghvh7qn2812e0i1b3he4 ),    
    
    .uf44audysjgtvdnua67       (ejddc553ql3y8eh4p8zbx9  ),
    .qtcasxm90cy0bwaqaxz     (gt8340_0a15il23cs0dyfy),
    .y38seii6ja77q2jy08       (rocadn0agggbhe8c7k6f  ),
    .f42g8ulc2y43ntmai5      (wa8alqpvm8_8wqh82v4 ),    
   
    .rgf8pa4kn20jusruz       (zffkoq91x2yrt8idy12  ),
    .wjwjffxr_4lulivwz     (cw8g0z3xpl_jmzl0bqsr4qz7r),
    .z6udkjbx164gh9yo1o      (c3o9e_kce6dj_oses5ebis ),
    .frkunk72hlttw0ar0np      (nl6qyr_h4vq399gjb47 ),    
  
    .r2tvaf8px0p9vlw4we       (ywnbexiz4zyc0xfli8  ),
    .srfn4smswwo6hbyaa     (fe0_jbuekwa1u_igwcjrf5),
    .a_u2kfmgv2ho357c      (ezoxoh6x_6pp3kplit2ipzy ),
    .svj88sv2u56fepzmg      (merrnyoykrdknka8adx1kp ),    
 
    .rzf167thmprvps0tm62i       (g0zewsbtm0xx173b6w3n  ),
    .lv7fu0hif2n2zhmgtcc     (ks8_k_t4av7jsxfssailx),
    .oj5t3f0lq1n9ae82x      (fuqvy5sh_dgu5b6_k5te2 ),
    .hat38salswlktk821      (s5br9ji17fis2ai4t5b257ui ),    

    .caxkrdjq0tjnnne9       (opg7to8zm4fdk0kbxb  ),
    .qpuk8ry0w9_r7ur4gcnx     (xuch6yvcgtv5auc_2s5g32),
    .v8jl1eh8o0n5g765      (c3es5lys6yhd7wv8lg2ho553 ),
    .c0xnu9p8he2hw10h      (buo4rvqs58con3m3n965h6a ),    


    .cgnsvvj7srbljqst     (cgnsvvj7srbljqst),

    .z8alxhlwgz117      (dm_t8xh6s80cssm), 
    .yafkacaefbdmi3hm6rvuao (moz9tdl4bhiltwpdv96jd),

    .q4j831gvqooep12      (fwgc_k58kjyp_va), 
    .u4frf_hcy8c0dh_aqkgsrp (j595qkrfu_okzcv0_4jxww_y_d),
  
    .tjzl_75hfxv6m          (p7ah58va5_2njbtv     ), 
    .ay20xnz1tx3gv1k     (u981qrwkgi5h0e72b__gg19w),  
    .fyo0ut7e82c         (p0i2i3v3j1tclelx51    ),  
     
    .tlwo81ky1a6b8         (tlwo81ky1a6b8 ),
    .l9x1ubg9wznb6ixv1i     (l9x1ubg9wznb6ixv1i ),
    .y5otpn351odm3mnpnfdshm (y5otpn351odm3mnpnfdshm),
    .rnlnwebfnqcg8g5oq_2gv0 (rnlnwebfnqcg8g5oq_2gv0),
    .bda77mp8zde61a_        (bda77mp8zde61a_),

    .gf33atgy               (gf33atgy       ),
    .ru_wi             (ru_wi     )  
  );



    
  assign k8qtf1i196m8bfpmqi = {f16zrowg1s1f5{1'b0}};

  
  wire mt9lk2yaup7e6ec3wdj77;
  wire mpuf2bhivkznq2s2owa;

  
  wire yvk2y9eyes = 
                     (st7pytysu10a & c5luf4ekdp8uxjd6phdb)
                   | (mh9ba4wb9dl & cik9g8nrdjspswqucoa9)
                   | j55vt_3172gxi8el;

  assign mt9lk2yaup7e6ec3wdj77 = (~yvk2y9eyes) & g3_8p4g7w5grnl62xy    ;
  assign vqwqaofc8sz_yjccd     = (~yvk2y9eyes) & mpuf2bhivkznq2s2owa;

  
  wire m5srj47yuxsm69zoep  = vt1176n4bhzdaz39cel8dhxqwrawhf;
  wire qkqin44n0uemg251 = wyyj6g00owlp1khb6vv9ycavglf;

  assign mpuf2bhivkznq2s2owa = m5srj47yuxsm69zoep & qkqin44n0uemg251
                              ;

  assign w0dzgnd8l98an1zx6ijhlbtalpk      = qkqin44n0uemg251 & mt9lk2yaup7e6ec3wdj77
                                         ;
  assign kcvmtch763q8ina8s4zil7kyspcf0      = m5srj47yuxsm69zoep  & mt9lk2yaup7e6ec3wdj77
                                         ;




  
  
  
  
  
  
  
  
  
  
  
  wire [5-1:0]      sz8s_i7k0mv2jx9rd    = pq05yc_ea9cb[4:0];
  wire [27-1:0]   jc617wq3856ziitfwye = pq05yc_ea9cb[(32-1):5];
  
  assign li2o0fhy6bmhmqeoi6rm = jc617wq3856ziitfwye[6-1:0];
  wire [21-1:0]        tp6b8miyf69e_4aaite = jc617wq3856ziitfwye[27-1:6];
  
  localparam ibwx_oi14egqf43e = 64;
  localparam l94ox50p53qz0lh = 6;
  wire[ibwx_oi14egqf43e-1:0] x61msl7z_lp;
  wire[ibwx_oi14egqf43e-1:0] k_vnkbf2ktlnc6omh;
  wire[ibwx_oi14egqf43e-1:0] i3ldxsak7bodk7;

  wire[ibwx_oi14egqf43e-1:0] cddnqnijha6ty;
  wire[ibwx_oi14egqf43e-1:0] xy1s4lgono9xpus4;
  wire[ibwx_oi14egqf43e-1:0] mrjljz6js9p2f3igcc6uu;
  wire[ibwx_oi14egqf43e-1:0] nn72wjjjexgf6jb2edi546n;
  wire[ibwx_oi14egqf43e-1:0] j23hrtjm_g7b1gs;

  wire[ibwx_oi14egqf43e-1:0] x5r2pynkila07uzj;
  wire[ibwx_oi14egqf43e-1:0] yaiy47p8coiq99;
  wire[ibwx_oi14egqf43e-1:0] vwpctvkryuytc;


  genvar i;

  generate 
      for (i=0; i<ibwx_oi14egqf43e; i=i+1) begin:ehbgy7v5lw63a25dg
    
    
    
    

        
        
        assign cddnqnijha6ty[i] = ecp10s0k_n91ef_jrkaki & (li2o0fhy6bmhmqeoi6rm[l94ox50p53qz0lh-1:0] == i[l94ox50p53qz0lh-1:0]);       
        assign xy1s4lgono9xpus4[i]  = q6dwr6kors49 & pirp8rqhngzyt0i6 & sh76lsmx & (li2o0fhy6bmhmqeoi6rm[l94ox50p53qz0lh-1:0] == i[l94ox50p53qz0lh-1:0]);      
        
        assign mrjljz6js9p2f3igcc6uu[i]  = k6_e3_saw0oup16pudov & (zpq6nysk8b654ynyt4zj9k[l94ox50p53qz0lh-1:0] == i[l94ox50p53qz0lh-1:0]);
        assign nn72wjjjexgf6jb2edi546n[i]  = pzfb_24lrjd770iigjx4sm & (d2lstp52x9w9900ioarrtfk[l94ox50p53qz0lh-1:0] == i[l94ox50p53qz0lh-1:0]);
        assign j23hrtjm_g7b1gs[i]  = mrjljz6js9p2f3igcc6uu[i] | nn72wjjjexgf6jb2edi546n[i];

        assign x5r2pynkila07uzj[i] = zwwbclwkk1c;
        assign yaiy47p8coiq99[i]  = zwwbclwkk1c;
        assign vwpctvkryuytc[i]  = (mrjljz6js9p2f3igcc6uu[i] & tq5w2fd0flcywep677l) | (nn72wjjjexgf6jb2edi546n[i] & juwj_oo3r8yt2a4hg);

        assign k_vnkbf2ktlnc6omh[i] = ( 
                                 cddnqnijha6ty[i]
                               | xy1s4lgono9xpus4[i]
                               | j23hrtjm_g7b1gs[i]
                                );

        assign i3ldxsak7bodk7[i] = ( 
                                 (cddnqnijha6ty[i] & x5r2pynkila07uzj[i])
                               | (xy1s4lgono9xpus4[i]  & yaiy47p8coiq99[i] )
                               | (j23hrtjm_g7b1gs[i]  & vwpctvkryuytc[i] )
                               );

        ux607_gnrl_dfflr #(1) omnwi1803vh2whp35 (k_vnkbf2ktlnc6omh[i], i3ldxsak7bodk7[i], x61msl7z_lp[i], gf33atgy, ru_wi);

      end
  endgenerate
  
  
  
      
  wire qvl0nalt9f5diijr = g3_8p4g7w5grnl62xy & vqwqaofc8sz_yjccd & (~jkq984ky8fozrzq);
  wire [l94ox50p53qz0lh-1:0] x0yljd7scw4jdpdfk3 = dlxukfkm1k19y_gskjb9vnl[l94ox50p53qz0lh-1:0];
  wire [l94ox50p53qz0lh-1:0] sfg4zdt9j_69cvw;

  ux607_gnrl_dfflr #(l94ox50p53qz0lh) sdv6ib_1rvye2bud2_ (qvl0nalt9f5diijr, x0yljd7scw4jdpdfk3, sfg4zdt9j_69cvw, gf33atgy, ru_wi);

  assign cgnsvvj7srbljqst = x61msl7z_lp[sfg4zdt9j_69cvw];






  wire tcbhrc_d0n7nn7r2gp;
  wire ic72uut7dw839dkvic186rezm;


  wire zox0zn2l32xutcve = (~nmqf8r7zm2wfw8pz) & (~b9b7j_s1j6pzebjxovfv6t) & ((j8cjhcuf0m6xjvemdaz & tia1md5dyh6kj4) | ysnexkrvlg2s55ajc5g69tm);

         
  assign i3r6fyspyh4r6kc73en3 = o9jixjnak_33vfbl & stdkgs3cetkrgnprgzkr;
  wire ek5id3cf6gcw0rjq = zox0zn2l32xutcve | i3r6fyspyh4r6kc73en3;
  wire [r4bbs1l72_cd3t_-1:0] uas9yj1olxg_qrsrgead8 = 
                                   zox0zn2l32xutcve ? {r4bbs1l72_cd3t_{1'b0}}
                                 : i3r6fyspyh4r6kc73en3 ? (eni2zaouo2xcn1_r + {{r4bbs1l72_cd3t_-1{1'b0}},1'b1})
                                 : eni2zaouo2xcn1_r;
  
  ux607_gnrl_dfflr #(r4bbs1l72_cd3t_) n6fd1wd9p_vg0xh6gy (ek5id3cf6gcw0rjq, uas9yj1olxg_qrsrgead8, eni2zaouo2xcn1_r, gf33atgy, ru_wi);
  
  wire dk56zdjblla1bkrom4cnnz6 = ysnexkrvlg2s55ajc5g69tm & (~oithmqsqi28np858lo1dztmf);
  wire w_cwdb_bx0n9qfjuj  = ysnexkrvlg2s55ajc5g69tm & oithmqsqi28np858lo1dztmf;
  wire ujmy3k2vmouuvq0    = (~ysnexkrvlg2s55ajc5g69tm) & j8cjhcuf0m6xjvemdaz & tia1md5dyh6kj4;

  wire w4krn94a6edmbd00u62h;

  wire lv8cgj36z2pwp2craly7bcjot;
  assign jywzcibo3cb08kg0a = lv8cgj36z2pwp2craly7bcjot | soj2j1b62_nupmoszxl45_ip;

  wire [r4bbs1l72_cd3t_-1:0] oii43c7aof50jnhvgi = 
      soj2j1b62_nupmoszxl45_ip ? {r4bbs1l72_cd3t_{1'b0}} : {r4bbs1l72_cd3t_{1'b1}}; 

  wire ak62trpnt64_2hcidbu83d = zox0zn2l32xutcve;
  wire j53ncrxv9wwr1z4_g3tpd8o = i3r6fyspyh4r6kc73en3 & (eni2zaouo2xcn1_r == oii43c7aof50jnhvgi);
  wire mhjh_wppzi2f0zswc4y = ak62trpnt64_2hcidbu83d | j53ncrxv9wwr1z4_g3tpd8o;
  wire pjwczzivvaeeb8nxavr = ak62trpnt64_2hcidbu83d;
  ux607_gnrl_dfflr #(1) nt6qvwy9b9gz8dgdfvjmx4vz (mhjh_wppzi2f0zswc4y, pjwczzivvaeeb8nxavr, o9jixjnak_33vfbl, gf33atgy, ru_wi);

  ux607_gnrl_dfflr #(1) tr1nngtvvdbisd_n_bd9unle04cd (ak62trpnt64_2hcidbu83d, dk56zdjblla1bkrom4cnnz6, lv8cgj36z2pwp2craly7bcjot, gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1) gnj011oqayj6nszfntmew8wcwv  (ak62trpnt64_2hcidbu83d, w_cwdb_bx0n9qfjuj , soj2j1b62_nupmoszxl45_ip , gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1) h94vsrz0oqjipt5qots7tujhjp2   (ak62trpnt64_2hcidbu83d, ujmy3k2vmouuvq0   , w4krn94a6edmbd00u62h   , gf33atgy, ru_wi);

  wire b_jq_m0xxmv006fkw6 = ysnexkrvlg2s55ajc5g69tm ? axgfwdkn0nyose7m3bwgcx92jc5gl61 : q7ru87fmzxczveihcxcwh;
  wire wabdz2q0q0gbkugcbjm = ysnexkrvlg2s55ajc5g69tm ? dyw1ymrkp8_lbpgb36w25d8fef1 : umc_2tn6um_9xaiy7_ksg0w;
  wire r8w8fpxoi98xpv8i = ysnexkrvlg2s55ajc5g69tm ? gq9tfy8ozjrgv8isn05omqqolwzip : uiyh4da4134sjv7gnmc;
  wire n2skbhe6fxja59uj659 = ysnexkrvlg2s55ajc5g69tm ? pvt527iyu2jjdtrzg1dhd0zi084q0nmww : 1'b0;
  wire r1px82knng5k016ja2ctpe_t = ysnexkrvlg2s55ajc5g69tm ? n3vgs5xww30vllhavnnqse8w0t8mrph : 1'b0;

  ux607_gnrl_dfflr #(1) g6nlqievu2w0y82q7ir9 (ak62trpnt64_2hcidbu83d, b_jq_m0xxmv006fkw6, ptmhu5qvej_2kw9w3pdr8, gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1) z3jgz6m3po5_7vapjk_8j1 (ak62trpnt64_2hcidbu83d, wabdz2q0q0gbkugcbjm, a3ybha5mrl8xcrr8, gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1) yehyzan9n_uyw7kt219h8b (ak62trpnt64_2hcidbu83d, r8w8fpxoi98xpv8i, oyd54mosns8enc8c, gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1) dlkr1ykfl_703kikpyzjlmv44r0_o (ak62trpnt64_2hcidbu83d, n2skbhe6fxja59uj659, hgpmlnfjch5bm27n3zz3vd, gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1) l60q2ijfga240b6ktdjsjlzhyjif (ak62trpnt64_2hcidbu83d, r1px82knng5k016ja2ctpe_t, nf6dcrwxlcch1sv8kmtkb_ry2, gf33atgy, ru_wi);
  
  assign dfqgbr7fyq0xiz172uj = o9jixjnak_33vfbl;


  wire m1hsvute2jmck3xkskdltq = j53ncrxv9wwr1z4_g3tpd8o;
  wire hbhowkp3zlgxun4o47j_ = tcbhrc_d0n7nn7r2gp & (~s_fxmgzl8pdoycnrftl7z7wz);
  wire nnz0wxl29fm83qt6b_v2o = m1hsvute2jmck3xkskdltq | hbhowkp3zlgxun4o47j_;
  wire fi84sb8q355o726aej = m1hsvute2jmck3xkskdltq;
  ux607_gnrl_dfflr #(1) zsh8gvijcrw277iif3fj (nnz0wxl29fm83qt6b_v2o, fi84sb8q355o726aej, tcbhrc_d0n7nn7r2gp, gf33atgy, ru_wi);

  
  wire ncrw4y6z8hn7qukcacrz3kolaehn = hbhowkp3zlgxun4o47j_;
  wire rmxclsditqfp46lc2sk_mkawky = ic72uut7dw839dkvic186rezm;
  wire sv36lgobs857ary_7vllugu8 = ncrw4y6z8hn7qukcacrz3kolaehn |   rmxclsditqfp46lc2sk_mkawky;
  wire w3hqhg874twer3vyyeb4i5iu = ncrw4y6z8hn7qukcacrz3kolaehn;
  ux607_gnrl_dfflr #(1) em2qu5v0cto_jky_8bu269css (sv36lgobs857ary_7vllugu8, w3hqhg874twer3vyyeb4i5iu, ic72uut7dw839dkvic186rezm, gf33atgy, ru_wi);
  

  wire pvz52yy2vzokr2ohsawza_egs;
  wire uytinyubmf6_8jxws4jpwztpa2 = j8cjhcuf0m6xjvemdaz & (~tia1md5dyh6kj4) & (~pvz52yy2vzokr2ohsawza_egs) & (~b9b7j_s1j6pzebjxovfv6t) ;
  wire gt7oixk8kvnp90dpbloevmn = pvz52yy2vzokr2ohsawza_egs;
  wire nu1742fz7syj4sm8p6hsskf = uytinyubmf6_8jxws4jpwztpa2 |   gt7oixk8kvnp90dpbloevmn;
  wire f74ck6k9z7iphg_0xjcuu7465i1 = uytinyubmf6_8jxws4jpwztpa2;
  ux607_gnrl_dfflr #(1) q777pd7iggzy9eqalwyg7ah0a6ezw (nu1742fz7syj4sm8p6hsskf, f74ck6k9z7iphg_0xjcuu7465i1, pvz52yy2vzokr2ohsawza_egs, gf33atgy, ru_wi);

  assign s_eowfyzlvx7gjv542upo = (ic72uut7dw839dkvic186rezm & w4krn94a6edmbd00u62h) | pvz52yy2vzokr2ohsawza_egs;


  assign nmqf8r7zm2wfw8pz = o9jixjnak_33vfbl | tcbhrc_d0n7nn7r2gp | ic72uut7dw839dkvic186rezm; 

  wire nve927ga5xugfv_y8aa6;
  wire dpwukg0syhkslzt657qf2c;
  wire ndslkzbikd36kmsxsxswgloxx77;
  wire oua72bcqsl0t2xpuadsbh97pazd3s;
  
  

  wire k1rq2k70b8y1eqkfccs5wuj = lv8cgj36z2pwp2craly7bcjot ? ncrw4y6z8hn7qukcacrz3kolaehn : 
                                               (  nve927ga5xugfv_y8aa6 
                                                | dpwukg0syhkslzt657qf2c
                                                ); 

  wire szf9ii2083hi9beh4zwln      = lv8cgj36z2pwp2craly7bcjot ? 1'b0 : nve927ga5xugfv_y8aa6 ? ndslkzbikd36kmsxsxswgloxx77      : 1'b0;
  wire r71c091gej74dwl__6brwtifoxm93dk = lv8cgj36z2pwp2craly7bcjot ? 1'b0 : nve927ga5xugfv_y8aa6 ? oua72bcqsl0t2xpuadsbh97pazd3s : 1'b0;
  


  assign nve927ga5xugfv_y8aa6      = fgru0fi7v178lp914d4zbdmqs63z_4 | tr_rxyj9lr38m35v2 | a03er8qo6p0zpb; 
  assign dpwukg0syhkslzt657qf2c  = w6m1johuy8qk9wgea0xqv12l_tkgb | bzsjo5unerpy5i0e_q_6eqn; 

  assign ndslkzbikd36kmsxsxswgloxx77 = (fgru0fi7v178lp914d4zbdmqs63z_4 & kngugv98d1yeo511y) | (a03er8qo6p0zpb & z8uuyp_3l6aqut86nkd__vvwgs);
  assign oua72bcqsl0t2xpuadsbh97pazd3s = (a03er8qo6p0zpb & z8uuyp_3l6aqut86nkd__vvwgs);
  

  
  
  

  ux607_gnrl_dfflr #(1) svgx7qzxb1c_2mpp5k74g    (1'b1              , k1rq2k70b8y1eqkfccs5wuj   , t1xtkdoie_8djygqlt1br56pwt   , gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1) klj0e05e9o016qoindm_n779z (k1rq2k70b8y1eqkfccs5wuj, szf9ii2083hi9beh4zwln, w33zvryieg8hhgy58581ny437h9, gf33atgy, ru_wi);
  
  ux607_gnrl_dfflr #(1) cp8bbseh7ij49p9rmh_cq4q5jlq_x_cg7 (k1rq2k70b8y1eqkfccs5wuj, r71c091gej74dwl__6brwtifoxm93dk, lv96t6re1w44borcb7do83ndua3vjy, gf33atgy, ru_wi);










  d7stl61zflp21cls1tg tm9w0cgdh85kersg7vk9 (
      .sxvvsxtbhyvt    (sxvvsxtbhyvt),
      .pcr4upio7_tx37     (pcr4upio7_tx37   ), 
      .uzklqlncpqqm1rav  (uzklqlncpqqm1rav),
      .ortueunvnkx_l5m_j  (ortueunvnkx_l5m_j),
      .hwuhtb7ucto_utk56  (hwuhtb7ucto_utk56),
      .i1env2kmns7qvvuuc  (i1env2kmns7qvvuuc),
      .g3s3vpafvy3i  (g3s3vpafvy3i),

      .rm1dxjejhq7dh3q5m  (rm1dxjejhq7dh3q5m ),

      .xatytj_r0fv14q  (coy3buxdw6yq3duh21azuwflk),
      .oily7           (hyec__ebnw8lbcssd81),
      .ly3dor8           (vs2610q9_on1r996p),
      .p1m           (1'b0),
      .u2k4dyp52s_m       (r_8h5lxb39ug57zli04e_o  ),
      .bktu0z1mk56       (pv7q0ikpayogkay57rgyr  ),
      .e98zc_xde8d        (t6l88yqbe4wokkhiso9t  ),

      .foj6m18         (dsq8f3rhmb7yc876v8  )
  );
      assign enu_vumk17eoj1fma5ilz0 = 1'b0;




      assign zp0aylmm0k4yw4w561bgzh = 1'b0;



endmodule
























module yjm16kn_qwdkfm8if #(
    parameter xl24j_imhfhfk = 64 
)(
    
  input                           stbblp081kc9,
  output                          vulpj3pebksw,
  input  [xl24j_imhfhfk      -1:0]    wbo1zx8iepki, 

  output                          z4qzurty_axomdd,
  input                           clwlpmx87nqbuq,
  output [xl24j_imhfhfk      -1:0]    atl5amsp8tyrm, 
  
  input                           j8kotg18hji,
  input  [32-1:0]    gebnakb8ctgri6s, 
  input  [1:0]                    rfdekem29gp7jx0f1, 
  output                          krasg_k9_i1zsgbu,
  output                          sf5oaemd1e3k,
  output reg [64-1:0]   ycj5xet5wunw0c,

  input                           pf8rzr1mv,
  input  [32-1:0]    rj1cfvu3meww, 
  input  [1:0]                    s2fbnn6ekvrsa3j, 
  output                          g_w2g5ygcfsk,
  output                          k4olvo5ol6hvag,
  output reg [64-1:0]   oivxcjfrvf9efavm,


  input                           x6n2fwiz0cogynnbie,
  input                           ncetuvy4lmo,
  input  [32-1:0]    diat9bfkf7mnu ,
  input  [64-1:0]       dn53sr7lydjdo5,
  input  [8-1:0]       hc79i6u2twxms6ke,
  output                          ybztfzzlexmx9gk,

  output ahth5hydygfua1j2,

  input  gf33atgy,
  input  ru_wi
);

  localparam bz6vmwhs94 = 4;
  localparam hermkomdto5zh1163m = (4-1);

  
  

  
  wire [4-1:0] d35brwhbkm;
  wire [4-1:0] xlzi7_mjg;
  wire [4-1:0] xayqet0sd;
  wire [4-1:0] d0x7t39v;
  wire [4-1:0] ycgzbt;

  wire [4-1:0] frdp1srjq7wfkr5pbrmm;
  wire [4-1:0] q0hvc42xv2;

  wire [64-1:0] c2daa2ko5tc1kr[4-1:0];
  wire [8-1:0] aju5nub5w4pdzi[4-1:0];
  wire [64-1:0] cdoijb57xe[4-1:0];
  wire [8-1:0] y5_ic3xhdy69h[4-1:0];

  wire [4-1:0] kuahmh7s6_xqs2foe43x;
  wire [4-1:0] junxbp4zh_8sbnuhivg;
  wire [4-1:0] k6h8pvd5a_4lon9b;
  wire [4-1:0] vfdzxjfvy8r0a;
  wire [4-1:0] kq41uyak08dennf9u0hjz7;
  wire [4-1:0] hmi_2i70n9b00b5ai_5;
  wire [4-1:0] tczedru9o1w;
  wire [4-1:0] pnqu6hzdxgr3tzg;
  wire [4-1:0] jewyarertntl;

  wire [64-1:0] h96b0cpofuouc122qnl_nu;

  

  wire  nkgylnugdg02yt;
  wire  [3-1:0] bwwdolbmwyxwyxwgwo;
  wire  [32-1:0] y0extssobeqgv;
  wire  [64   -1:0] oiq72xcdyk9;
  wire  [8   -1:0] fejl08khwu6;

  wire  a9sylku3twkk                     ;
  wire  [3-1:0] ze1rhnlau2i_0pibby9;
  wire  [32-1:0] ifvinhzxvs ;
  wire  [64   -1:0] y7bezxcu0bihmj1;
  wire  [8   -1:0] fabu73o9b99e6u;

  assign {
           nkgylnugdg02yt
         , bwwdolbmwyxwyxwgwo
         , y0extssobeqgv
         , oiq72xcdyk9
         , fejl08khwu6
        } = wbo1zx8iepki;

  assign atl5amsp8tyrm = {
           a9sylku3twkk
         , ze1rhnlau2i_0pibby9
         , ifvinhzxvs
         , y7bezxcu0bihmj1
         , fabu73o9b99e6u
        };

  wire                        xc9nkzc0ylsp[4-1:0]; 
  wire  [3-1:0] xijb062z22fxf026o50  [4-1:0]; 
  wire  [32-1:0] i00quc3x43h  [4-1:0]; 
  wire  [64   -1:0] esmp6teq31 [4-1:0]; 
  wire  [8   -1:0] po7c9zrn [4-1:0]; 
  
  
  wire [2-1:0] klzlbzxf9k70;

  
  wire [2-1:0] oyd91wgthmz3b;


  wire l0kqs5qujoo = stbblp081kc9 & vulpj3pebksw;
  wire f8fvunfazuj5_ = z4qzurty_axomdd & clwlpmx87nqbuq;

  
  
  wire s2roq9roe5is258;
  wire lvs4u7g1bwtxpvtjs5ip = ~s2roq9roe5is258;
  wire daabtq8vpy8e9ysdyler = (klzlbzxf9k70 == hermkomdto5zh1163m[2-1:0]) & l0kqs5qujoo;
  
  ux607_gnrl_dfflr #(1) w__bu901_di1711if (daabtq8vpy8e9ysdyler, lvs4u7g1bwtxpvtjs5ip, s2roq9roe5is258, gf33atgy, ru_wi);
  
  wire [2-1:0] wenl_o0vzxw21; 
  
  assign wenl_o0vzxw21 = daabtq8vpy8e9ysdyler ? 2'b0 : (klzlbzxf9k70 + {{2-1{1'b0}},1'b1});
  
  ux607_gnrl_dfflr #(2) zcv9x2s5ku87ej (l0kqs5qujoo, wenl_o0vzxw21, klzlbzxf9k70, gf33atgy, ru_wi);
      

  
  wire l1n5t8iv0_vlbjd5zd;
  wire y3afem4lrnejnhp = ~l1n5t8iv0_vlbjd5zd;
  wire zhp697t12otd9bwfzm = (oyd91wgthmz3b == hermkomdto5zh1163m[2-1:0]) & f8fvunfazuj5_;
  
  ux607_gnrl_dfflr #(1) n16_5zxk07a0qcr6mhm8 (zhp697t12otd9bwfzm, y3afem4lrnejnhp, l1n5t8iv0_vlbjd5zd, gf33atgy, ru_wi);
  
  wire [2-1:0] ntnwjp6se52b; 
  
  assign ntnwjp6se52b = zhp697t12otd9bwfzm ? 2'b0 : (oyd91wgthmz3b + {{2-1{1'b0}},1'b1});

  ux607_gnrl_dfflr #(2) tbxo_34b0860av (f8fvunfazuj5_, ntnwjp6se52b, oyd91wgthmz3b, gf33atgy, ru_wi);

  wire z8cy652mi3r = (oyd91wgthmz3b == klzlbzxf9k70) &   (l1n5t8iv0_vlbjd5zd == s2roq9roe5is258);
  wire yn5im8g4q1q  = (oyd91wgthmz3b == klzlbzxf9k70) & (~(l1n5t8iv0_vlbjd5zd == s2roq9roe5is258));


  wire [2-1:0] nfpvh8kxawm = f8fvunfazuj5_ ? ntnwjp6se52b : oyd91wgthmz3b;
  wire [2-1:0] vcs61nqhoxgn = l0kqs5qujoo ? wenl_o0vzxw21 : klzlbzxf9k70;
  wire zqcutsvzb_gemc83n = daabtq8vpy8e9ysdyler ? lvs4u7g1bwtxpvtjs5ip : s2roq9roe5is258;
  wire v54xzfv9t09t7zx41 = zhp697t12otd9bwfzm ? y3afem4lrnejnhp : l1n5t8iv0_vlbjd5zd;
  assign ahth5hydygfua1j2  = (nfpvh8kxawm == vcs61nqhoxgn) & (~(v54xzfv9t09t7zx41 == zqcutsvzb_gemc83n));

  wire [8-1:0] v7bd_280i0ax6zgyif;
  wire [8-1:0] nelwc61day117q;

  genvar i;
  generate 
      for (i=0; i<bz6vmwhs94; i=i+1) begin:tz9npc7nthu18o8k3
  
        assign d35brwhbkm[i] = l0kqs5qujoo & (klzlbzxf9k70 == i[2-1:0]);
        assign xlzi7_mjg[i] = f8fvunfazuj5_ & (oyd91wgthmz3b == i[2-1:0]);
        assign xayqet0sd[i] = d35brwhbkm[i] |   xlzi7_mjg[i];
        assign d0x7t39v[i] = d35brwhbkm[i];
  
        ux607_gnrl_dfflr #(1) hdti_6iaq (xayqet0sd[i], d0x7t39v[i], ycgzbt[i], gf33atgy, ru_wi);

        
        ux607_gnrl_dfflr #(32) c3x_7a0gzdh083r  (d35brwhbkm[i], y0extssobeqgv, i00quc3x43h[i], gf33atgy, ru_wi);
        ux607_gnrl_dfflr #(3) mx66bo7c6g17z4wydvajk3  (d35brwhbkm[i], bwwdolbmwyxwyxwgwo, xijb062z22fxf026o50[i], gf33atgy, ru_wi);
        ux607_gnrl_dfflr #(1) l9l0w_szl5rbp4  (d35brwhbkm[i], nkgylnugdg02yt, xc9nkzc0ylsp[i], gf33atgy, ru_wi);

        
        assign frdp1srjq7wfkr5pbrmm[i] = x6n2fwiz0cogynnbie & jewyarertntl[i];
        assign c2daa2ko5tc1kr[i] = (esmp6teq31[i] & (~h96b0cpofuouc122qnl_nu)) | (dn53sr7lydjdo5 & h96b0cpofuouc122qnl_nu);
        assign aju5nub5w4pdzi[i] = (po7c9zrn[i] | hc79i6u2twxms6ke);
        assign q0hvc42xv2[i] = d35brwhbkm[i] | frdp1srjq7wfkr5pbrmm[i];
        assign cdoijb57xe[i] = d35brwhbkm[i] ? oiq72xcdyk9 : c2daa2ko5tc1kr[i];
        assign y5_ic3xhdy69h[i] = d35brwhbkm[i] ? fejl08khwu6 : aju5nub5w4pdzi[i];
        ux607_gnrl_dfflr #(64) qe0462bbwrbueuv (q0hvc42xv2[i], cdoijb57xe[i], esmp6teq31[i], gf33atgy, ru_wi);
        ux607_gnrl_dfflr #(8) ju5da9jomeiuaoh3 (q0hvc42xv2[i], y5_ic3xhdy69h[i], po7c9zrn[i], gf33atgy, ru_wi);

      assign kuahmh7s6_xqs2foe43x[i] = (gebnakb8ctgri6s[32-1:3] == i00quc3x43h[i][32-1:3]) & ycgzbt[i];
      assign junxbp4zh_8sbnuhivg[i] = ((v7bd_280i0ax6zgyif & po7c9zrn[i]) == v7bd_280i0ax6zgyif) & ycgzbt[i];  

      assign vfdzxjfvy8r0a[i] = j8kotg18hji & kuahmh7s6_xqs2foe43x[i] & (~(junxbp4zh_8sbnuhivg[i]));  
      assign k6h8pvd5a_4lon9b [i] = j8kotg18hji & kuahmh7s6_xqs2foe43x[i] &   (junxbp4zh_8sbnuhivg[i]) ;  

      assign kq41uyak08dennf9u0hjz7[i] = (rj1cfvu3meww[32-1:3] == i00quc3x43h[i][32-1:3]) & ycgzbt[i];
      assign hmi_2i70n9b00b5ai_5[i] = ((nelwc61day117q & po7c9zrn[i]) == nelwc61day117q) & ycgzbt[i];  

      assign pnqu6hzdxgr3tzg[i] = pf8rzr1mv & kq41uyak08dennf9u0hjz7[i] & (~(hmi_2i70n9b00b5ai_5[i]));  
      assign tczedru9o1w [i] = pf8rzr1mv & kq41uyak08dennf9u0hjz7[i] &   (hmi_2i70n9b00b5ai_5[i]) ;  

      assign jewyarertntl[i] = x6n2fwiz0cogynnbie & ncetuvy4lmo & 
          (diat9bfkf7mnu[32-1:3] == i00quc3x43h[i][32-1:3]) & ycgzbt[i];

  
      end
  endgenerate

  assign sf5oaemd1e3k = (| k6h8pvd5a_4lon9b);
  assign krasg_k9_i1zsgbu = (| vfdzxjfvy8r0a);
  assign k4olvo5ol6hvag = (| tczedru9o1w);
  assign g_w2g5ygcfsk = (| pnqu6hzdxgr3tzg);
  assign ybztfzzlexmx9gk = (| jewyarertntl);

  assign ze1rhnlau2i_0pibby9 = xijb062z22fxf026o50[oyd91wgthmz3b];
  assign a9sylku3twkk = xc9nkzc0ylsp[oyd91wgthmz3b];
  assign ifvinhzxvs   = i00quc3x43h  [oyd91wgthmz3b];
  assign y7bezxcu0bihmj1  = esmp6teq31 [oyd91wgthmz3b];
  assign fabu73o9b99e6u  = po7c9zrn [oyd91wgthmz3b];

  assign z4qzurty_axomdd  = ~z8cy652mi3r;
  assign vulpj3pebksw  = ~yn5im8g4q1q;

  integer j;

  always @ * begin: mksbtsddhz
    ycj5xet5wunw0c = 64'b0;
    oivxcjfrvf9efavm = 64'b0;
    for (j=0; j<bz6vmwhs94; j=j+1) begin
      ycj5xet5wunw0c = (ycj5xet5wunw0c | ({64{k6h8pvd5a_4lon9b[j]}} & esmp6teq31[j])); 
      oivxcjfrvf9efavm = (oivxcjfrvf9efavm | ({64{tczedru9o1w[j]}} & esmp6teq31[j])); 
    end
  end


  generate 
      if(64 == 64) begin:fjcbdq
                assign v7bd_280i0ax6zgyif =
                                      (rfdekem29gp7jx0f1 == 2'b00) ? (8'b1 << gebnakb8ctgri6s[2:0]) : 
                                      (rfdekem29gp7jx0f1 == 2'b01) ? (8'b11 << {gebnakb8ctgri6s[2:1],1'b0}) : 
                                      (rfdekem29gp7jx0f1 == 2'b10) ? (8'b1111 << {gebnakb8ctgri6s[2],2'b0}) : 
                                               8'b1111_1111; 
                assign nelwc61day117q =
                                      (s2fbnn6ekvrsa3j == 2'b00) ? (8'b1 << rj1cfvu3meww[2:0]) : 
                                      (s2fbnn6ekvrsa3j == 2'b01) ? (8'b11 << {rj1cfvu3meww[2:1],1'b0}) : 
                                      (s2fbnn6ekvrsa3j == 2'b10) ? (8'b1111 << {rj1cfvu3meww[2],2'b0}) : 
                                               8'b1111_1111; 
            assign h96b0cpofuouc122qnl_nu = {
                           {8{hc79i6u2twxms6ke[7]}},
                           {8{hc79i6u2twxms6ke[6]}},
                           {8{hc79i6u2twxms6ke[5]}},
                           {8{hc79i6u2twxms6ke[4]}},
                           {8{hc79i6u2twxms6ke[3]}},
                           {8{hc79i6u2twxms6ke[2]}},
                           {8{hc79i6u2twxms6ke[1]}},
                           {8{hc79i6u2twxms6ke[0]}}
                    };
      end
      if(64 == 32) begin:g2z3f
                assign v7bd_280i0ax6zgyif =
                                      (rfdekem29gp7jx0f1 == 2'b00) ? (8'b1 << gebnakb8ctgri6s[1:0]) : 
                                      (rfdekem29gp7jx0f1 == 2'b01) ? (8'b11 << {gebnakb8ctgri6s[1],1'b0}) : 
                                               8'b1111; 
                assign nelwc61day117q =
                                      (s2fbnn6ekvrsa3j == 2'b00) ? (8'b1 << rj1cfvu3meww[1:0]) : 
                                      (s2fbnn6ekvrsa3j == 2'b01) ? (8'b11 << {rj1cfvu3meww[1],1'b0}) : 
                                               8'b1111; 
            assign h96b0cpofuouc122qnl_nu = {
                           {8{hc79i6u2twxms6ke[3]}},
                           {8{hc79i6u2twxms6ke[2]}},
                           {8{hc79i6u2twxms6ke[1]}},
                           {8{hc79i6u2twxms6ke[0]}}
                    };
      end
  endgenerate


endmodule





















module neplroszbk3r28 (

  input                          f5jobxqu5r8tdcgp9dz_,
  input                          hfh_n8b2_6ltn5lve4_271m, 
  output                         xiy2xcok2j1vz3hdn21fq8us4e, 
  input  [32-1:0]   ezq9pnmedz815gxhjrvk5x, 
  input                          gs8s9g8gtij6u619m3tcdcvnd,   
  input                          i36cd1y8_65k09dz0thns,   
  input                          wb6ynztvqw_c7jt0r60z0a3,   
  input                          rykqnjd3sew6zqm077moncthemet9, 
  input                          z2oi9osh3p0wy7vb2sr69u07, 
  input                          n1ko5ud3mahcu4f2t8,
  input                          k250aa9_7n16_xye3p__d4ew7, 
  input                          p4_cbhjumvsd2_nee5pbvt1, 
  input                          m63kr3yu_6uz_m3_yti5_e9,
  input  [64-1:0]        at3xavrqfa9vpvz2wfl28m2, 
  input  [8-1:0]     zawrb3vcmuri8b2986t8n2f, 
  input  [1:0]                   y_nw0z1jiz_z1j47b284ciw,
  input                          sxokdo7nllqwvltwlem22uf5,
  input  [4 -1:0] z_l3eykrjali3v1mh46uf5mt,
  input                          jis_avsh9dp0zny0zshz7,
  input  [4:0]                   tudsip00rgu_1pit8jhrmcjt35cbx,
  input                          z_rab_1o8tf_6vir         ,
  input                          as_mlum8anvtnrny9tls     ,
  input                          fd8f2gq4oaalsv4p_j     ,


  input                           y5qvboneeuu7u9c6ex2k32,
  input                           r0b984qp4dbimt7m049jn,
  input [4-1:0]    eq0u1926xaldb_6z8t8xdam,

  input                           vhfqvbg0i9tkhk8b7_1xw94s_n3h,
  input [4-1:0]    hn6ha7kpsoxids4i7ilrw,
  input                           o4tmdwuwe0a_icm5c4xc3pnm0,
  input [64-1:0]          qelk6ys1izwqop2178az43,  

  input                           pdl18ljotymfj543wtjh49b_r,
  input [4-1:0]    kavx5xx6zd8f9hqjq1s,
  input                           wt6jy410rpokxn04lscbst6uo7,
  input [64-1:0]          z8hscmi55sjt_ufebya9e, 


  input                           slk31s106jz ,


  output                          o21b8ypt1xiu5ml63d,
  output                          vrsqde4muadsevgpemk, 
  output                          badsf4ksbp3k6p_p5hnj2i, 
  input                           ed4kcy8s9nrisftgx_q, 
  output  [32-1:0]   bdqo1tgw2_bpi2e8alini, 
  output                          jp5nha2l14e7kx2jzpke,   
  output                          za9xg3zsqni_aeqmke,   
  output                          c1gmncmorg16sachdas,   
  output                          p648zxn2luyxy8mt992a, 
  output                          uxlldm0w_h7kicit8gvhqv2, 
  output                          yvu98r_7ji4o250r_u,
  output                          zdpamqgv7ddf1n3x5t2q, 
  output                          wpsukhyqhl92dzoam7cm, 
  output                          v3oo69y614hgiemyyld,
  output  [64-1:0]        a4a48egkdkec8d9b_9, 
  output  [8-1:0]     xwfmltfzahuj4qfn4qf2, 
  output  [1:0]                   ggxoqcj7ytp1a4pjf7ee,
  output                          l3c127qdc9a2mfc13,
  output  [4 -1:0] oq9b5zfhza9yvdoj,
  output  [4:0]                   szrgf24or2mbt7w_yleh_vt,
  output  yixt0a_xmh    ,
  output  fgnb7mhn1254le9     ,
  output  okt7c24tca9ji6pw     ,
  output                          sg33s7pt45jp_,
  output                          g9i9mf8jq7sc699j,

  output  f0jwv0n5olimpf4vnvqpb4hs,

  input                           gf33atgy,
  input                           ru_wi
);


  wire a7ysdemx0o8a;

  wire zoqg7ispio42di7;
  wire km6b8_2zng1v1727ro7r16p9w40;
  wire [32-1:0]   xlr6euqcclj1jbf65vsoh;

  wire ax49i75tk  =  gs8s9g8gtij6u619m3tcdcvnd;
  wire fzs1etb5tv44 = ~gs8s9g8gtij6u619m3tcdcvnd;

  wire n5ekwdb0o5itvvs8ue5 = (ezq9pnmedz815gxhjrvk5x[32-1:3] == xlr6euqcclj1jbf65vsoh[32-1:3]);
  wire s51qsmhp1c_b7z9dj  = (z2oi9osh3p0wy7vb2sr69u07 && km6b8_2zng1v1727ro7r16p9w40);




  wire hgs200wa1m8dtm_w;
  wire zwi7ocpler3zip7ma6;
  wire j50h2yer70l    = f5jobxqu5r8tdcgp9dz_ & ax49i75tk;
  wire gvipokeyosuvmdnu  = hfh_n8b2_6ltn5lve4_271m & ax49i75tk;
  wire x6n2fwiz0cogynnbie = hfh_n8b2_6ltn5lve4_271m & fzs1etb5tv44;
  assign xiy2xcok2j1vz3hdn21fq8us4e = ax49i75tk ? hgs200wa1m8dtm_w : zwi7ocpler3zip7ma6;


  wire bt9shzgcqycs6o193 = (n5ekwdb0o5itvvs8ue5 | s51qsmhp1c_b7z9dj) & zoqg7ispio42di7;


  wire vk7jhl80iumbqk_3;
  wire icu69kziufvljht01;
  wire   vswwz4xrpct   =  j50h2yer70l & (~bt9shzgcqycs6o193);
  assign vk7jhl80iumbqk_3 =  gvipokeyosuvmdnu & (~bt9shzgcqycs6o193);
  assign  hgs200wa1m8dtm_w = icu69kziufvljht01 & (~bt9shzgcqycs6o193);


  wire gwcyc814yd2z3f_yac;
  wire dfrmcobjfbgcscnbwb;
  assign gwcyc814yd2z3f_yac =  x6n2fwiz0cogynnbie & (~slk31s106jz);
  assign  zwi7ocpler3zip7ma6 = dfrmcobjfbgcscnbwb;
  wire ggidb_bkj8keqqas0e = gwcyc814yd2z3f_yac & dfrmcobjfbgcscnbwb;


  wire   t3wgx9jv4z1;
  wire   wlx00s9xnmgqyit2;
  wire   wmxaigx2sgoy8itlh4eb;
  assign wlx00s9xnmgqyit2  = a7ysdemx0o8a & zoqg7ispio42di7;
  assign t3wgx9jv4z1      = a7ysdemx0o8a & wmxaigx2sgoy8itlh4eb;


  wire   bvjm3irn;
  wire   rqvv9111 = ~bvjm3irn; 
  assign wmxaigx2sgoy8itlh4eb = (~rqvv9111) ? ed4kcy8s9nrisftgx_q : 1'b0; 
  assign icu69kziufvljht01   =   rqvv9111  ? ed4kcy8s9nrisftgx_q : 1'b0; 

  assign badsf4ksbp3k6p_p5hnj2i = (~rqvv9111) ? wlx00s9xnmgqyit2 : vk7jhl80iumbqk_3;
  assign o21b8ypt1xiu5ml63d   = (~rqvv9111) ? wlx00s9xnmgqyit2 : f5jobxqu5r8tdcgp9dz_;






  wire h9ug7pjno9e97phd4i6dqm9a;
  wire kq2tv38wrsn8rl6io2zinvji;
  wire [4 -1:0]qb4t55busoetvxyb1ooe0_ork;



   wire p9_84ph0rjoughfop3hoar  = (eq0u1926xaldb_6z8t8xdam == hn6ha7kpsoxids4i7ilrw);
   wire crcgb75c2p1m4uf2_1r_i_4yrkoi = p9_84ph0rjoughfop3hoar 
                                & hfh_n8b2_6ltn5lve4_271m 
                                & vhfqvbg0i9tkhk8b7_1xw94s_n3h 
                                & o4tmdwuwe0a_icm5c4xc3pnm0 
                                ;

   wire ahanzmie8jevvv7dc6ns = (eq0u1926xaldb_6z8t8xdam == kavx5xx6zd8f9hqjq1s);
   wire f3fhpzgqn9xwyeotqxgl_rv9q2v = ahanzmie8jevvv7dc6ns 
                                & hfh_n8b2_6ltn5lve4_271m 
                                & pdl18ljotymfj543wtjh49b_r 
                                & wt6jy410rpokxn04lscbst6uo7 
                                ;

   wire ocx7icyptl8yx45bth  = (qb4t55busoetvxyb1ooe0_ork == hn6ha7kpsoxids4i7ilrw);
   wire o601g4iirycoggsgoakybqixpbt = ocx7icyptl8yx45bth 
                                & zoqg7ispio42di7 
                                & vhfqvbg0i9tkhk8b7_1xw94s_n3h 
                                & o4tmdwuwe0a_icm5c4xc3pnm0 
                                ;

   wire v3hx0p8qlgg1fxhefr8 = (qb4t55busoetvxyb1ooe0_ork == kavx5xx6zd8f9hqjq1s);
   wire ny986k5uwa4ks78avxt35c5g = v3hx0p8qlgg1fxhefr8 
                                & zoqg7ispio42di7 
                                & pdl18ljotymfj543wtjh49b_r 
                                & wt6jy410rpokxn04lscbst6uo7 
                                ;

   wire [64-1:0] xv5to55_4wd = 

                               ({64{crcgb75c2p1m4uf2_1r_i_4yrkoi}} & qelk6ys1izwqop2178az43)
                             | ({64{f3fhpzgqn9xwyeotqxgl_rv9q2v}} & z8hscmi55sjt_ufebya9e)
                             ; 
   wire [64-1:0] e_bpogyelz0h = 

                               ({64{o601g4iirycoggsgoakybqixpbt}} & qelk6ys1izwqop2178az43)
                             | ({64{ny986k5uwa4ks78avxt35c5g}} & z8hscmi55sjt_ufebya9e)
                             ; 


   wire [64-1:0] awpq068vos = y5qvboneeuu7u9c6ex2k32   ? {xv5to55_4wd} : at3xavrqfa9vpvz2wfl28m2; 
   wire [64-1:0] k67tywvm9gpl = e_bpogyelz0h; 
   wire [64-1:0] swbwo112tnd = ggidb_bkj8keqqas0e ? awpq068vos : k67tywvm9gpl; 

   wire aortxa8s4madvjc4hl0k = crcgb75c2p1m4uf2_1r_i_4yrkoi | f3fhpzgqn9xwyeotqxgl_rv9q2v;
   wire ndxvcg8tfubzpvch6k1 = o601g4iirycoggsgoakybqixpbt | ny986k5uwa4ks78avxt35c5g;
   wire w36v74h15xbskqsaro = aortxa8s4madvjc4hl0k & y5qvboneeuu7u9c6ex2k32;
   wire agtf8ysq1jyhkuqgf = ndxvcg8tfubzpvch6k1 & h9ug7pjno9e97phd4i6dqm9a;

   wire yy95v2lcrr0n8sm = ggidb_bkj8keqqas0e ? w36v74h15xbskqsaro : agtf8ysq1jyhkuqgf;
   wire n2e11ebegn = ((~y5qvboneeuu7u9c6ex2k32) & ggidb_bkj8keqqas0e) 
                | (y5qvboneeuu7u9c6ex2k32 & (yy95v2lcrr0n8sm))
                ; 
   wire wxdjral4lf5c2fx7hq7  = ggidb_bkj8keqqas0e | yy95v2lcrr0n8sm;


   wire pupx4lmyufv2tqr =((~w36v74h15xbskqsaro) & y5qvboneeuu7u9c6ex2k32);
   wire h5mmt5uzjkl0fo7t3 = (~agtf8ysq1jyhkuqgf) & h9ug7pjno9e97phd4i6dqm9a;
   wire cy4nzm6_1ruro5f0 = ggidb_bkj8keqqas0e ? pupx4lmyufv2tqr : h5mmt5uzjkl0fo7t3;
   wire p9y5qthv_fd9v02 = ggidb_bkj8keqqas0e | yy95v2lcrr0n8sm;
   ux607_gnrl_dfflr #(1) hkc07ites1nqbtb9hnb9a (p9y5qthv_fd9v02, cy4nzm6_1ruro5f0  , h9ug7pjno9e97phd4i6dqm9a, gf33atgy, ru_wi);
   ux607_gnrl_dfflr #(1) ttmzrwajq_oy8lrw9(ggidb_bkj8keqqas0e, r0b984qp4dbimt7m049jn  , kq2tv38wrsn8rl6io2zinvji, gf33atgy, ru_wi);

   ux607_gnrl_dfflr #(4) in087sdgbxzqur (ggidb_bkj8keqqas0e, eq0u1926xaldb_6z8t8xdam , qb4t55busoetvxyb1ooe0_ork, gf33atgy, ru_wi);


   assign a7ysdemx0o8a   =  
                             (~h9ug7pjno9e97phd4i6dqm9a) 
                           ; 

   assign bvjm3irn = wlx00s9xnmgqyit2 & (~vswwz4xrpct);





  wire                         umlpb7ug9u9ws19jrwdxs;
  wire                         xzlbb89vuod_lc4_xarf4kej;
  wire                         xlusu5ifu2aflibdjuhicwm0x;
  wire                         tq5sx_z9_t4jpv208g5ng9vlm;
  wire                         j50743oeax1_3gfxf2vz5;
  wire                         gyru72xtej7h4shu14x_z5j5;
  wire                         yb86l7sjetx5cim3w8idgxwq4;
  wire                         f1f7nvfc7fb60khqq2wug;
  wire [64-1:0]        zd0o_ghc5adq6b1dd1ptlg4k7c;
  wire [8-1:0]     jdx5ia6o5r3ij075yytcemij1b;
  wire [1:0]                   fge8n71ryohm7_z0f1qo;
  wire                         kay0p1u7ais56ny_dmxpw56x;
  wire [4 -1:0] u3pt6klbfknzseuthp55i;
  wire                         ndkzxobymtej5hw5fq729     ;

  wire                         ybn66n27s68gu2t ;
  wire                         hf5x5xai5qs00i_3wv ;



  wire [64-1:0]        uinxud0ci62m6byypbsensjbv6p;

  ux607_gnrl_dfflr #(32)  kc73g02c3fp4pncc2p     (ggidb_bkj8keqqas0e, ezq9pnmedz815gxhjrvk5x    , xlr6euqcclj1jbf65vsoh    , gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1              )  u1wbplrusswlrozp37wxn33     (ggidb_bkj8keqqas0e, gs8s9g8gtij6u619m3tcdcvnd    , umlpb7ug9u9ws19jrwdxs    , gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1              )  g16_6j1ez5ouo4b72ym     (ggidb_bkj8keqqas0e, i36cd1y8_65k09dz0thns    , xzlbb89vuod_lc4_xarf4kej    , gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1              )  yd8di2zz3nu2fmmfx7s8j     (ggidb_bkj8keqqas0e, wb6ynztvqw_c7jt0r60z0a3    , xlusu5ifu2aflibdjuhicwm0x    , gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1)                frojz68z7q4l7gbl7796553 (ggidb_bkj8keqqas0e, rykqnjd3sew6zqm077moncthemet9, tq5sx_z9_t4jpv208g5ng9vlm, gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1)                kbpl85ej20rnc7mhkwrzkmj   (ggidb_bkj8keqqas0e, z2oi9osh3p0wy7vb2sr69u07  , km6b8_2zng1v1727ro7r16p9w40  , gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1)                v3cca17fbqfhpm8pd3w       (ggidb_bkj8keqqas0e, n1ko5ud3mahcu4f2t8      , j50743oeax1_3gfxf2vz5      , gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1)                s1k1ser9ux9jn07ht322j4w    (ggidb_bkj8keqqas0e, k250aa9_7n16_xye3p__d4ew7   , gyru72xtej7h4shu14x_z5j5   , gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1)                nj0mvrxuniqzed96az1f377b    (ggidb_bkj8keqqas0e, p4_cbhjumvsd2_nee5pbvt1   , yb86l7sjetx5cim3w8idgxwq4   , gf33atgy, ru_wi);

  ux607_gnrl_dfflr #(1)                tpz9_j1mrt3j7o_macr6    (ggidb_bkj8keqqas0e, m63kr3yu_6uz_m3_yti5_e9   , f1f7nvfc7fb60khqq2wug   , gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(8)    exdu6cdbfgag8rv6lodfx    (ggidb_bkj8keqqas0e, zawrb3vcmuri8b2986t8n2f   , jdx5ia6o5r3ij075yytcemij1b   , gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(2)                eirxg5_7u7k84liplcxc     (ggidb_bkj8keqqas0e, y_nw0z1jiz_z1j47b284ciw    , fge8n71ryohm7_z0f1qo    , gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1)                kb6yatwrucex308a0vap    (ggidb_bkj8keqqas0e, sxokdo7nllqwvltwlem22uf5   , kay0p1u7ais56ny_dmxpw56x   , gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(4) qv3xrjok_6e09ykbiz7pn7     (ggidb_bkj8keqqas0e, z_l3eykrjali3v1mh46uf5mt    , u3pt6klbfknzseuthp55i    , gf33atgy, ru_wi);
  assign ndkzxobymtej5hw5fq729     =  1'b0;

  ux607_gnrl_dfflr #(1)                bt4jptciakzbxyc096l4s(ggidb_bkj8keqqas0e, as_mlum8anvtnrny9tls        , ybn66n27s68gu2t    , gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1)                vfmtjxlg5snc75cbzp1(ggidb_bkj8keqqas0e, fd8f2gq4oaalsv4p_j        , hf5x5xai5qs00i_3wv    , gf33atgy, ru_wi);

  ux607_gnrl_dfflr #(64)       n7h24daextrh0sys0fur_d8    (wxdjral4lf5c2fx7hq7, swbwo112tnd                 , zd0o_ghc5adq6b1dd1ptlg4k7c   , gf33atgy, ru_wi);

     ux607_gnrl_pipe_stage # (
      .CUT_READY(0),
      .DP(1),
      .DW(1)
     ) rahye864u7dz0uqw_ (
       .i_vld(gwcyc814yd2z3f_yac), 
       .i_rdy(dfrmcobjfbgcscnbwb), 
       .i_dat(1'b0 ),
       .o_vld(zoqg7ispio42di7), 
       .o_rdy(t3wgx9jv4z1), 
       .o_dat( ),

       .clk  (gf33atgy  ),
       .rst_n(ru_wi)  
      );



   assign vrsqde4muadsevgpemk     = bvjm3irn ? 1'b0                           : slk31s106jz;
   assign bdqo1tgw2_bpi2e8alini      = bvjm3irn ? xlr6euqcclj1jbf65vsoh           : ezq9pnmedz815gxhjrvk5x    ;
   assign jp5nha2l14e7kx2jzpke      = bvjm3irn ? umlpb7ug9u9ws19jrwdxs           : gs8s9g8gtij6u619m3tcdcvnd    ;
   assign za9xg3zsqni_aeqmke      = bvjm3irn ? xzlbb89vuod_lc4_xarf4kej           : i36cd1y8_65k09dz0thns    ;
   assign c1gmncmorg16sachdas      = bvjm3irn ? xlusu5ifu2aflibdjuhicwm0x           : wb6ynztvqw_c7jt0r60z0a3    ;
   assign p648zxn2luyxy8mt992a  = bvjm3irn ? tq5sx_z9_t4jpv208g5ng9vlm       : rykqnjd3sew6zqm077moncthemet9;
   assign uxlldm0w_h7kicit8gvhqv2    = bvjm3irn ? km6b8_2zng1v1727ro7r16p9w40         : z2oi9osh3p0wy7vb2sr69u07  ;
   assign yvu98r_7ji4o250r_u        = bvjm3irn ? j50743oeax1_3gfxf2vz5             : n1ko5ud3mahcu4f2t8   ;                   
   assign zdpamqgv7ddf1n3x5t2q     = bvjm3irn ? gyru72xtej7h4shu14x_z5j5          : k250aa9_7n16_xye3p__d4ew7; 
   assign wpsukhyqhl92dzoam7cm     = bvjm3irn ? yb86l7sjetx5cim3w8idgxwq4          : p4_cbhjumvsd2_nee5pbvt1; 
   assign v3oo69y614hgiemyyld     = bvjm3irn ? f1f7nvfc7fb60khqq2wug          : m63kr3yu_6uz_m3_yti5_e9; 
   assign ggxoqcj7ytp1a4pjf7ee      = bvjm3irn ? fge8n71ryohm7_z0f1qo           : y_nw0z1jiz_z1j47b284ciw ;
   assign l3c127qdc9a2mfc13     = bvjm3irn ? kay0p1u7ais56ny_dmxpw56x          : sxokdo7nllqwvltwlem22uf5;
   assign oq9b5zfhza9yvdoj      = bvjm3irn ? u3pt6klbfknzseuthp55i           : z_l3eykrjali3v1mh46uf5mt ;

   assign a4a48egkdkec8d9b_9     = uinxud0ci62m6byypbsensjbv6p  ;
   assign xwfmltfzahuj4qfn4qf2     = jdx5ia6o5r3ij075yytcemij1b       ;

  assign  yixt0a_xmh =   z_rab_1o8tf_6vir ; 
  assign fgnb7mhn1254le9     = bvjm3irn ? ybn66n27s68gu2t  : as_mlum8anvtnrny9tls;
  assign okt7c24tca9ji6pw     = bvjm3irn ? hf5x5xai5qs00i_3wv  : fd8f2gq4oaalsv4p_j;










   assign sg33s7pt45jp_          = zoqg7ispio42di7 | jis_avsh9dp0zny0zshz7 ;

   assign szrgf24or2mbt7w_yleh_vt = 5'b0;



   assign uinxud0ci62m6byypbsensjbv6p = 
            ({64{fge8n71ryohm7_z0f1qo == 2'b00}} & {8{zd0o_ghc5adq6b1dd1ptlg4k7c[ 7:0]}})
          | ({64{fge8n71ryohm7_z0f1qo == 2'b01}} & {4{zd0o_ghc5adq6b1dd1ptlg4k7c[15:0]}})
          | ({64{fge8n71ryohm7_z0f1qo == 2'b10}} & {2{zd0o_ghc5adq6b1dd1ptlg4k7c[31:0]}})
          | ({64{fge8n71ryohm7_z0f1qo == 2'b11}} &    zd0o_ghc5adq6b1dd1ptlg4k7c[63:0])
          ;









  assign f0jwv0n5olimpf4vnvqpb4hs = zoqg7ispio42di7;
  assign g9i9mf8jq7sc699j = zoqg7ispio42di7;

endmodule



















module urpfdi55wfwmmi3i (


  input                         k8qtud5yr1e98g, 
  output                        mw1zdgavbul7ic, 
  input [64-1:0]        covjtr51ggzngufqow,
  input [4 -1:0] qfhwjs9ygxr4e0rg86a,
  input                         r86mhhg0562g6n9sah0z , 
  input                         drgmlg58l2czwg2ijhc,
  input                         hvgjjhizbfp9km9dd,
  input [64 -1:0]  nd1hj8zlmdgys5obof18pe,
  input [64 -1:0]  oe3uwa3e_ggymrc7ri,
  input                         aqz_nh46x0w0rdwc83s7c , 
  input                         oor8acg0u_d09e0moah , 
  input [4:0]                   a51im30isjous61asad1lrg5,



  input                         eapsrdy52u,
  input                         slk31s106jz,

  output                         vz63qkw5s3m8urb9, 
  output [64-1:0]        iojqlhtwx45_siz,
  output [4 -1:0] ydtm1yuxqj7fmxvqc,

  output                         jfsrn6g5wjvu1s, 
  input                          a726ykhkw2fkfxd, 
  output [64-1:0]        sml00v8pmuueefw,
  output [4 -1:0] ewg8titgu69y7lmx0j,
  output                         hz3c9eiwgzw2hb , 
  output                         xbzkx8ucmech,
  output                         ehkpciu6l7p,
  output [64 -1:0]  jm0nv8cdtqhyk5t2ddht,
  output [64 -1:0]  oo04o1rrd2a,
  output                         mxu7x8rtlq0kewjvcl , 
  output                         p4pen8le4jxeud_b , 
  output [4:0]                   eqedamf6p97lmc2ywq,

  output                         b0ylmw5xa8oytsw3j6n,


  input                           gf33atgy,
  input                           ru_wi
);


  wire          mgjqsgpiza1dr;


  wire qqlfmnnkeewqaepmyz6;
  wire ifpwpn9cje7ts6ay7bl42;
  wire ld9r25q2ljqxxvw743hecl;
  wire zpzhpz0yx4dz0z6ce12tc8o;


  wire          zvyiwdpyvt;
  wire          o0ozobxf1oc2t5;
  wire          jf92hqkj0cxz;
  wire          qos62pcur8;
  wire          jae1i1kz83d2c; 

  wire uv0i532o = jae1i1kz83d2c;


  wire nusxc051gyf44jr4o =  drgmlg58l2czwg2ijhc & (~uv0i532o);
  assign qqlfmnnkeewqaepmyz6   = k8qtud5yr1e98g & (~nusxc051gyf44jr4o);




  assign mw1zdgavbul7ic    = (nusxc051gyf44jr4o | ifpwpn9cje7ts6ay7bl42) ;






  assign vz63qkw5s3m8urb9   = k8qtud5yr1e98g & uv0i532o ;
  assign iojqlhtwx45_siz    = covjtr51ggzngufqow ;
  assign ydtm1yuxqj7fmxvqc    = qfhwjs9ygxr4e0rg86a ;



  wire vtrh64t_ilwd_7kg1 = eapsrdy52u;

  wire c36vprtr19jh3 = drgmlg58l2czwg2ijhc & (k8qtud5yr1e98g & mw1zdgavbul7ic); 

  assign  zvyiwdpyvt  = vtrh64t_ilwd_7kg1;

  assign  jf92hqkj0cxz = ~slk31s106jz;

  assign  qos62pcur8 = c36vprtr19jh3;

   ux607_gnrl_fifo # (
         .DP(8+1),
         .DW(1),
         .CUT_READY(0) 
    ) t70bb97y4ddu44l9r5v0b(
      .i_vld   (zvyiwdpyvt),
      .i_rdy   (o0ozobxf1oc2t5),
      .i_dat   (jf92hqkj0cxz),
      .o_vld   (mgjqsgpiza1dr),
      .o_rdy   (qos62pcur8),
      .o_dat   (jae1i1kz83d2c),
      .clk     (gf33atgy  ),
      .rst_n   (ru_wi)
    );


  assign b0ylmw5xa8oytsw3j6n =  mgjqsgpiza1dr; 



  localparam epef6ura = 
                       64                
                     + 4          
                     + 1                         
                     + 1                         
                     + 1                         
                     + 5                         
                     + 64           
                     + 64           
                     + 1                         
                     + 1                         
                     ;
  wire [epef6ura-1:0] t6rrba8f52_htbc39, yqwvj28rv36_pyx4;
  assign t6rrba8f52_htbc39 = {
                             covjtr51ggzngufqow  ,
                             qfhwjs9ygxr4e0rg86a  ,
                             r86mhhg0562g6n9sah0z   ,
                             drgmlg58l2czwg2ijhc     ,
                             hvgjjhizbfp9km9dd     ,
                             a51im30isjous61asad1lrg5 , 
                             nd1hj8zlmdgys5obof18pe,
                             oe3uwa3e_ggymrc7ri     ,
                             aqz_nh46x0w0rdwc83s7c , 
                             oor8acg0u_d09e0moah  
                            };

    assign {
            sml00v8pmuueefw,
            ewg8titgu69y7lmx0j,
            hz3c9eiwgzw2hb ,
            xbzkx8ucmech  ,
            ehkpciu6l7p  ,
            eqedamf6p97lmc2ywq,
            jm0nv8cdtqhyk5t2ddht,
            oo04o1rrd2a     ,
            mxu7x8rtlq0kewjvcl , 
            p4pen8le4jxeud_b  
           } = yqwvj28rv36_pyx4;



      ux607_gnrl_pipe_stage # (
       .CUT_READY(0),
       .DP(1),
       .DW(epef6ura)
      ) h6fpifhw62e2gmr (
        .i_vld(qqlfmnnkeewqaepmyz6), 
        .i_rdy(ifpwpn9cje7ts6ay7bl42), 
        .i_dat(t6rrba8f52_htbc39 ),
        .o_vld(ld9r25q2ljqxxvw743hecl), 
        .o_rdy(zpzhpz0yx4dz0z6ce12tc8o), 
        .o_dat(yqwvj28rv36_pyx4 ),

        .clk  (gf33atgy  ),
        .rst_n(ru_wi)  
       );


  assign jfsrn6g5wjvu1s     = ld9r25q2ljqxxvw743hecl ;
  assign zpzhpz0yx4dz0z6ce12tc8o = a726ykhkw2fkfxd;

endmodule


















module upb8yfyhriv8e (

  input dn8riluj40uunvq5,
  input w92a5o09fp9dg6, 
  input eglor15f7p2ivpny5dc, 


  output bhjn0b8ydp0vfsiy,
  input [32-1:0] yh9n8rxd7xt9w6cyy9,
  input [32-1:0] r0bsza4vt3629icr,




  output o4qff84vfbn, 
  input  x74_jhmpouk, 
  output [64-1:0] z5tnbveujliw633sxlb8,
  output [4 -1:0] l8ng5e_pa1fg07__37,
  output erdoc9bbdnq8065yw , 
  output ro93aearv5754gz9w, 
  output [64 -1:0] y9389ymcyh2ia2082yx1_,
  output [64 -1:0] uiu4_g7j41kz,
  output zqx1cj9lvt0e,
  output zsxgccndqw2suf6,
  output [4:0] ytp8_jsqr2sjmu08gdn,





  input                          qzarx9bid_hex85cnt,
  input                          wg5jouh0rdnsnk8kgtlq,
  input                          i0o9d6dhf5giw4uln5c,
  input  [4:0]                   szrgf24or2mbt7w_yleh_vt,
  input                          o21b8ypt1xiu5ml63d, 

  input                          badsf4ksbp3k6p_p5hnj2i, 
  input                          vrsqde4muadsevgpemk, 
  output                         ed4kcy8s9nrisftgx_q, 
  input  [32-1:0]   bdqo1tgw2_bpi2e8alini, 
  input                          jp5nha2l14e7kx2jzpke,   
  input                          uxlldm0w_h7kicit8gvhqv2,
  input                          yvu98r_7ji4o250r_u,
  input                          zdpamqgv7ddf1n3x5t2q,
  input                          wpsukhyqhl92dzoam7cm,
  input                          v3oo69y614hgiemyyld,
  input  [64-1:0]        a4a48egkdkec8d9b_9, 
  input  [8-1:0]     xwfmltfzahuj4qfn4qf2, 
  input                          za9xg3zsqni_aeqmke,
  input                          c1gmncmorg16sachdas,
  input  [1:0]                   ggxoqcj7ytp1a4pjf7ee,
  input                          p648zxn2luyxy8mt992a, 
  input                          l3c127qdc9a2mfc13,
  input  [4 -1:0] oq9b5zfhza9yvdoj,
  input                          sg33s7pt45jp_,

  input                          g9i9mf8jq7sc699j,


  output                         flcopog5zzpohfautwy, 
  input                          gtb8f_h0g28itdr8k, 
  output                         wf15djwi2hw25nz_  , 
  output                         t1q5qmk9jzpf6glng4y,
  output [64-1:0]        xsmx4zoewhbt07jxq,


  
  
  
  
  input                          cxrbvs1hde7j8ziudd4ar,
  output                         dmzxpdd5dgmp_2ip6h3_6,
  input  [32-1:0]     piv1ndd8n8dlaqx9, 
  input                          r3rgwuaokuw68zin, 
  input                          m2aue5rcrjkbzdwbqvlzvr, 
  input                          u7a8_cbg_zi4w4b4slc08, 
  input                          fd_1f891ni339pnyzw63mg, 
  input                          zqnzorh6g9hnwsot5zr, 
  input                          wic6t212ob4tfa, 
  input  [64-1:0]      p1g5jbgswdsx9v1j01103,
  input  [8-1:0]      zmrmpw_9vyme3rakn8br8e,
  input                          sp2wnouu73ujsanhkn0,
  input                          n5w05rcecv47nvnfkkw5,
  input  [1:0]                   dycy3iz66xw6yj5ea,

  
  output                         ro76scx3ggmfi4xp2bjx,
  input                          t9yh0n7ay27ft001vimu6,
  output                         gpjxeoxkmf35ldn  ,
  output                         owde01ai01h2x5kn3_ng,
  output [64-1:0]      atur2zwqwk4mnbtz68l2,

  
  
  
  
  input                          fkm9up63o1aeauaqhjb,
  output                         to_1lv9wnb3vmu6tvz5rc,
  input  [32-1:0]   ju1kbeplcqy314lfj4, 
  input                          r985fbe5k7hgzaq9i, 
  input                          bb04gpwotp2s6c7_p1gqkq, 
  input                          sqmey185cu3mtixhl, 
  input                          rffcsd1o699ytclmx,
  input                          roa7ljysjukna1_f_rh5l, 
  input                          swz29iuutp9bjf_, 
  input  [64-1:0]        lbr88vbqtg8rht7320frde,
  input  [8-1:0]     g7qq38mx3d58n1b15kcia,
  input                          demg_fwfkmaeawq30t,
  input                          grtb6ypa0px2gi1c,
  input  [1:0]                   f128d8ws0seoihu1,
  
  output                         m2r7mfmq3afdd1ine,
  input                          nhafiywg3hg_52kogwh,
  output                         xrqayy6vigrw66z8a  ,
  output                         jyy72ywt9nbo10f2jxupacld,
  output [64-1:0]        drz92qecqx_qtxwro,































  output                         k5t515v6aa4oilq98cy6lrd8,
  output                         nbgnnsuqy2oogaz89vmbl1,
  input                          lkdpdaxvpxpy8w8hpchiph,
  output [32-1:0]   c1_3zcfvbhkc9cf7jgm7x, 
  output                         sk43hkjk_z2mer7becad, 
  output                         cki2l53v3p6py9awsecgj, 
  output                         ddjl2wsfh12b286nsrl3m5z, 
  output                         y09wfhff_yx31yoe7cxv, 
  output                         zn80vi7_hafilb62kh72jx5d6, 
  output                         e1wmvmyg_x8tobsfzpo, 
  output [64-1:0]        lo0fo8wk5o04f7ezwv474,
  output [8-1:0]     zutoko8hik1j9pa64jmpuw,
  output                         xqdmvgffpmzj6n0l23o,
  output                         of_yab2i0nf9xv_tek5r,
  output [1:0]                   i1pzsd21aml3amhex3sf,


  input                          ltzq1n1rg2b9lrt8j0bs__wa,
  output                         qui4zelf64bknwchxnz6,
  input                          qf_hxpj8b9rdyabqx8q7l  ,
  input                          pqfnz7dk2f2khe5zxq0081lzv,
  input  [64-1:0]        j3gop6yag94s712e_mipwr484,


  
  
  
  
  
  output                         hr7la0400ty0hiwk5d0,
  input                          y1ipzdhzcfq282ups6ja,
  output [32-1:0]   lqv5bv6hq78ov_prb97v5z, 
  output                         uarhtvlb5te5hc2g3, 
  output                         o15lm7no18top00l32ra, 
  output                         ly1y__c5rzaa9xv_9_m1ppr, 
  output                         f1msmreidlchd7rf9w625, 
  output [64-1:0]        g9ayxf51lhjl44vvw62u3,
  output [8-1:0]      qfoijjxktg6dht3klxhyw5g,
  output                         gao2lzva86gawlwp2,
  output                         xpt7vgmhw7tamcpv2l,
  output [1:0]                   lrh4lctjvrz1rhm6b9oh,
  output                         krh62hs2scfnb76m67a,
  output                         pyfc_rgr3cwwvo34pf,
  output                         u6xj18ku9lj1890n7,
  output                         s3lwpy5def9adgbbvx9ct,
  output                         q96vjidg4x6ohxl7,
  
  
  input                          b6m1vcd7bmemxnu99_zke,
  output                         vqld30a8qt13mzhwoc,
  input                          jpa5gwkjwqz_j0a3cy1  ,
  input                          kjxe2fpsacp9bx2_0fah36ij,
  input  [64-1:0]        xsw8oz2ni13z6vac1tn61,




  
  
  
  output                         c0x_72w8ddbpt17fn,
  
  
  output                         tw0yf9aln_vu06k8l,
  input                          q84eo09gg53r2jj5a5xn,
  output [16-1:0]   ss4cm882613f24kdjqsyl, 
  output                         oefdpb9h9kx627r_0y5, 
  output                         zm9uosdggg7ntkh97elw, 
  output                         g_ahl2zik6mj75atnp_hej, 
  output                         bjl40q8m35dwdn_mn9, 
  output [64-1:0]        fh1jm1za5zvqmvdloi,
  output [8-1:0]      sp_0hv_ae5rrl9vagusi,
  output                         b4oh48a9a0g269ybrm,
  output                         r5s3ykb7_xkl6t12oucf,
  output [1:0]                   ssswxj_bpfx_ebsbj,
  
  
  input                          fsj22rallxmhdrvuwenpq,
  output                         yign8d_dhrow0i5wjts4bd,
  input                          hhlfu4md9k5v7naf1qt  ,
  input                          j8m9s_du9fk99idlbh80  ,
  input  [64-1:0]        aapsfpke41r7dyya4ah,


  
  
  
  output                         y1rlahaedj99shvl6uc,
  
  
  output                         rqf8b5xxbw0n1_qaw,
  input                          ocwcf75wgxfb1bawe,
  output [16-1:0]   holgl43_yucp7f7l, 
  output                         gy2sgn_1bpkac7msq3, 
  output                         oyev1ipmdflkvxygwr, 
  output                         ihknw7_lm_572tv6s, 
  output                         o31l03k34sdhwt4lkazfa5, 
  output [64-1:0]        r_1u6q2lzkfus3o9nfl,
  output [8-1:0]      yff7wf8wth2vjkdjpr,
  output                         lppjhpov_5lgvx7n7fm4g,
  output                         sdfg9zykj79rz_7thf9k,
  output [1:0]                   wt4e4tlh0u_4cljr2j5f9,
  
  
  input                          o4wuryrcvw13y2v5m6b6u,
  output                         bt4howrm5xnf6u4fuwrum6,
  input                          vnqegbzme0jutvf  ,
  input                          jdj122rbumyogtin6xpg97  ,
  input  [64-1:0]        p9mcc6npaw32uigcp6,


  input  gf33atgy,
  input  ru_wi
  );

  wire [32-1:0] r480zryu00zrqkrbk = 32'h00000000;
  wire [32-1:0] zys87dxafg7t5ll4o9 = 32'h0c000000;
  wire [32-1:0] o4f5s69ex_fk0k7q13x = 32'h08000000;
  wire [32-1:0] rqbq0wq0_ojyw61v5 = 32'h02000000;
  wire [32-1:0] dak283_f21dou11_grfkt = 32'h10000000;










          localparam y7fi7kw8i180nr4b   = 3;
          localparam senagm_wgrp66rwiuyf1d = 2;










  wire                  c0l6w8lh_td7pzkcpdfp0ir_t;
  wire                  a_pr26ts5th7p3ziyczhdy;
  wire                  r22ymekw52k08rw4tm0  ;
  wire                  zdg2ytmoa2dqi_9xntu0hld3fx;
  wire [64-1:0] wsxqohy8uxi3mw1ruq9o5z2;

  wire                         af66zf64p_pphlj9uy240vtnsz; 
  wire                         gt923cnjxl9zc1kavj6ay3l6vo6; 
  wire                         y3cb9jdvssvccg6b1mqbt7jl_;
  wire                         gx8_jfgud1t_azz9c19jh;
  wire                         g1au1uuxkz40lxd494d7ma;
  wire [2-1:0]                 nxjbs9v14ld33363ewcmdo1;
  wire [4 -1:0] uyma7dg_jtxevl8vmljt;
  wire [32-1:0]   jqxmjq8am07ckn333alfaky1b;
  wire cf_fu13q7n0up5qevsfiq5xf788; 
  wire l0aco1cxtoml1g4byoibwl; 
  wire zs25fw9ohsy43_e2z409h0jq;
  wire dant527kjskp0aikp8_70;
  wire desv6k9j3glnmlfx0hu30ots6i;
  wire xedpt5e1vonpdv78parohexbw;
  wire bzjsole_y2xxo6diyfseg;
  wire [4:0] vh0mg3miltnw_b4o_ga66yzvjx;


  localparam s3xvyho = (4+9+32+1+5+1+1)
                     + 1
                     + 1 
                     ;
  localparam q_ldd1waoilf7q1 = 3;
  localparam ale66u8k_50s8h4vdf4 = 2;
  localparam a69a9ho1_kmpwc58n = 1;
  localparam y61y499cunmtec = 0;
  localparam au8wnhbd2ozhfnnm = q_ldd1waoilf7q1+1;
  localparam qn77zdua2lv05_ = au8wnhbd2ozhfnnm+1;

  localparam bvma5mx5x4uqrf = s3xvyho-1; 
  wire [s3xvyho-1:0] m8adyck2et7e0qcwg_ =
      {
         vrsqde4muadsevgpemk  
        ,p648zxn2luyxy8mt992a  
        ,l3c127qdc9a2mfc13
        ,jp5nha2l14e7kx2jzpke
        ,ggxoqcj7ytp1a4pjf7ee
        ,oq9b5zfhza9yvdoj 
        ,bdqo1tgw2_bpi2e8alini 
        ,qzarx9bid_hex85cnt 
        ,i0o9d6dhf5giw4uln5c 
        ,szrgf24or2mbt7w_yleh_vt 
        ,wpsukhyqhl92dzoam7cm
        ,yvu98r_7ji4o250r_u
        ,c1gmncmorg16sachdas 
        ,uxlldm0w_h7kicit8gvhqv2 
        ,zdpamqgv7ddf1n3x5t2q 
        ,v3oo69y614hgiemyyld 
      };


  wire [s3xvyho-1:0] nhyv494899nv6d2 =
      {
         1'b0 
        ,1'b0
        ,1'b0
        ,r985fbe5k7hgzaq9i
        ,f128d8ws0seoihu1
        ,4'b0
        ,ju1kbeplcqy314lfj4 
        ,1'b0 
        ,5'b0 
        ,sqmey185cu3mtixhl 
        ,swz29iuutp9bjf_
        ,grtb6ypa0px2gi1c 
        ,roa7ljysjukna1_f_rh5l 
        ,bb04gpwotp2s6c7_p1gqkq 
        ,rffcsd1o699ytclmx 
      };

  wire [s3xvyho-1:0] t3ysg7mwfhqy_9hje;
  wire [s3xvyho-1:0] n1lhs71oc209opa;

  wire [s3xvyho-1:0] hlhiqyobvyaycq770rym =
      {
         1'b0
        ,1'b0
        ,1'b0
        ,r3rgwuaokuw68zin
        ,dycy3iz66xw6yj5ea
        ,4'b0
        ,piv1ndd8n8dlaqx9 
        ,1'b0
        ,1'b0
        ,4'b0
        ,u7a8_cbg_zi4w4b4slc08
        ,wic6t212ob4tfa
        ,n5w05rcecv47nvnfkkw5 
        ,zqnzorh6g9hnwsot5zr 
        ,m2aue5rcrjkbzdwbqvlzvr 
        ,fd_1f891ni339pnyzw63mg 
      };



  wire [s3xvyho-1:0]      zxgpsirnmn33k29fvgm;
  assign 
      {
         af66zf64p_pphlj9uy240vtnsz  
        ,gt923cnjxl9zc1kavj6ay3l6vo6  
        ,y3cb9jdvssvccg6b1mqbt7jl_
        ,gx8_jfgud1t_azz9c19jh
        ,nxjbs9v14ld33363ewcmdo1
        ,uyma7dg_jtxevl8vmljt 
        ,jqxmjq8am07ckn333alfaky1b
        ,xedpt5e1vonpdv78parohexbw
        ,bzjsole_y2xxo6diyfseg
        ,vh0mg3miltnw_b4o_ga66yzvjx
        ,dant527kjskp0aikp8_70
        ,l0aco1cxtoml1g4byoibwl
        ,g1au1uuxkz40lxd494d7ma 
        ,cf_fu13q7n0up5qevsfiq5xf788 
        ,zs25fw9ohsy43_e2z409h0jq
        ,desv6k9j3glnmlfx0hu30ots6i
      } = zxgpsirnmn33k29fvgm;


  wire ouat_m1vwjc0l5igzo2z4g;
  wire sw9511te5wakyzkx_xdo;

  wire gyja61p9t197hw65hvyi63g;
  wire [32-1:0] v10jhardhhvft6w6t3u;
  wire mrrzsfopopzgqr_nro5;
  wire [64-1:0] pp5egelk49dgurfb3w;
  wire [8-1:0] n9sl3nl16qlprh9ocn6trcs;
  wire l1368lp6updfhsbebtzpc;
  wire rvqfn2hxjfeh8egdvsc;
  wire [1:0] c55olxxsckol_k4eb9fyu;
  wire [2:0] g3iy6vml027o3gv9wt;
  wire [1:0] z0y5vk22vnz94pcxx;
  wire [s3xvyho-1:0] jmo524gyok0abs1u1;

  wire k8aii0cb2ywh7xvp5ud9 = jmo524gyok0abs1u1[a69a9ho1_kmpwc58n]; 
  wire vyaut44yc_lmxpxuhm = jmo524gyok0abs1u1[qn77zdua2lv05_]; 
  wire t06t7flkpby01affnv56x64 = jmo524gyok0abs1u1[y61y499cunmtec];

  wire n0wp_tjsit08gjo9ggcxe_a;
  wire ebnc6trwg85shv8_iz8qpa2;
  wire n93c2nog4f68lktvd0;
  wire uezhv2clc8f9woh7dc5ss1;
  wire [64-1:0] j2p0ug10na1wztrfj39;
  wire [s3xvyho-1:0] guqjz9gxv28q8f719;

  wire qywrqdqbkmyeridmga5k;
  wire ya7at6mg3adjqzbi1c6;
  wire l8ymtznl9hcobcfqg;
  wire ybmlc9yctmeh5ymbek57;
  wire [64-1:0] z4lyw1_nvshizqbim5x;
  wire [s3xvyho-1:0] s_s052pc2p3r_9o280580;


  wire [y7fi7kw8i180nr4b*1-1:0] ccxw7l8izxzjj14ozqkgvvyd6;

  wire [y7fi7kw8i180nr4b*1-1:0] k1_j5ubhqqpfrl3p0bi186va9;
  wire [y7fi7kw8i180nr4b*1-1:0] w0hjg2xow0ymilw7bcxpm2l;
  wire [y7fi7kw8i180nr4b*32-1:0] xzpsiztjmn62eb967x1xkc6;
  wire [y7fi7kw8i180nr4b*1-1:0] a_dm6kd_qbw2cv84wtboltif01;
  wire [y7fi7kw8i180nr4b*64-1:0] ae00o9ay050qc5d5zxf18282b92;
  wire [y7fi7kw8i180nr4b*8-1:0] puxr8jzij0m30qcwmdz2sufl51;
  wire [y7fi7kw8i180nr4b*1-1:0] s6vj39lt1yt7f1ytk3pr3;
  wire [y7fi7kw8i180nr4b*1-1:0] wspjbjcpf459zy17qhyz8jmqy7;
  wire [y7fi7kw8i180nr4b*2-1:0] y7jg1o7n3jl52fxr0isdv8;
  wire [y7fi7kw8i180nr4b*s3xvyho-1:0] w8o2oxw46tp1zf4rujrx4zyxw;
  wire [y7fi7kw8i180nr4b*3-1:0] sxjmcdip1m7ighns0k5aue59fj;
  wire [y7fi7kw8i180nr4b*2-1:0] noyjdh392j1x0s9g1b_lk;

  wire [y7fi7kw8i180nr4b*1-1:0] qkiytqsa_fo9x5ls7yb_x1k2;
  wire [y7fi7kw8i180nr4b*1-1:0] idw2i93am7m9wy_5hzipgymj5k3;
  wire [y7fi7kw8i180nr4b*1-1:0] wzmdtyq65i82w_tt0juwqle;
  wire [y7fi7kw8i180nr4b*1-1:0] kz10yoaxkacgm38dwv37tl2ixfv;
  wire [y7fi7kw8i180nr4b*64-1:0] fyvkbec2dn4rlcslyiyttfrx;
  wire [y7fi7kw8i180nr4b*s3xvyho-1:0] od5a1yudx9bmyqpwleexh4h9;

  wire rsugt_kl1l2oy2_snu6nd; 
  wire j5xn5cw86bpa3g6q9k_ly7;

  assign rsugt_kl1l2oy2_snu6nd = (~g9i9mf8jq7sc699j) & cxrbvs1hde7j8ziudd4ar    ;
  assign dmzxpdd5dgmp_2ip6h3_6     = (~g9i9mf8jq7sc699j) & j5xn5cw86bpa3g6q9k_ly7;


  assign k1_j5ubhqqpfrl3p0bi186va9 =
                           {
                             badsf4ksbp3k6p_p5hnj2i
                           , fkm9up63o1aeauaqhjb
                           , rsugt_kl1l2oy2_snu6nd
                           } ;


  wire jivto5soso7t2shjdzdtpo3 = 1'b0;
  wire nv8nvom_0jskth8 = 1'b0;

  wire rx5ecsbhut83vs55c   = 1'b0;

  assign ccxw7l8izxzjj14ozqkgvvyd6 =

                           {

                             (o21b8ypt1xiu5ml63d | sg33s7pt45jp_)
                           , fkm9up63o1aeauaqhjb
                           , (rsugt_kl1l2oy2_snu6nd)
                           } ;



  assign xzpsiztjmn62eb967x1xkc6 =
                           {
                             bdqo1tgw2_bpi2e8alini
                           , ju1kbeplcqy314lfj4
                           , piv1ndd8n8dlaqx9
                           } ;

  assign a_dm6kd_qbw2cv84wtboltif01 =
                           {
                             jp5nha2l14e7kx2jzpke
                           , r985fbe5k7hgzaq9i
                           , r3rgwuaokuw68zin
                           } ;

  assign ae00o9ay050qc5d5zxf18282b92 =
                           {
                             a4a48egkdkec8d9b_9
                           , lbr88vbqtg8rht7320frde
                           , p1g5jbgswdsx9v1j01103
                           } ;

  assign puxr8jzij0m30qcwmdz2sufl51 =
                           {
                             xwfmltfzahuj4qfn4qf2
                           , g7qq38mx3d58n1b15kcia
                           , zmrmpw_9vyme3rakn8br8e
                           } ;

  assign s6vj39lt1yt7f1ytk3pr3 =
                           {
                             za9xg3zsqni_aeqmke
                           , demg_fwfkmaeawq30t
                           , sp2wnouu73ujsanhkn0
                           } ;

  assign sxjmcdip1m7ighns0k5aue59fj =
                           {
                             3'b0
                           , 3'b0
                           , 3'b0
                           } ;

  assign noyjdh392j1x0s9g1b_lk =
                           {
                             2'b0
                           , 2'b0
                           , 2'b0
                           } ;

  assign wspjbjcpf459zy17qhyz8jmqy7 =
                           {
                             c1gmncmorg16sachdas
                           , grtb6ypa0px2gi1c
                           , n5w05rcecv47nvnfkkw5
                           } ;

  assign y7jg1o7n3jl52fxr0isdv8 =
                           {
                             ggxoqcj7ytp1a4pjf7ee
                           , f128d8ws0seoihu1
                           , dycy3iz66xw6yj5ea
                           } ;

  assign w8o2oxw46tp1zf4rujrx4zyxw =
                           {
                             m8adyck2et7e0qcwg_
                           , nhyv494899nv6d2
                           , hlhiqyobvyaycq770rym
                           } ;


  assign                   {
                             ed4kcy8s9nrisftgx_q
                           , to_1lv9wnb3vmu6tvz5rc
                           , j5xn5cw86bpa3g6q9k_ly7
                           } = w0hjg2xow0ymilw7bcxpm2l;




  assign                   {
                             c0l6w8lh_td7pzkcpdfp0ir_t
                           , m2r7mfmq3afdd1ine
                           , ro76scx3ggmfi4xp2bjx
                           } = qkiytqsa_fo9x5ls7yb_x1k2;

  assign                   {
                             r22ymekw52k08rw4tm0
                           , xrqayy6vigrw66z8a
                           , gpjxeoxkmf35ldn
                           } = wzmdtyq65i82w_tt0juwqle;

  assign                   {
                             zdg2ytmoa2dqi_9xntu0hld3fx
                           , jyy72ywt9nbo10f2jxupacld
                           , owde01ai01h2x5kn3_ng
                           } = kz10yoaxkacgm38dwv37tl2ixfv;


  assign                   {
                             wsxqohy8uxi3mw1ruq9o5z2
                           , drz92qecqx_qtxwro
                           , atur2zwqwk4mnbtz68l2
                           } = fyvkbec2dn4rlcslyiyttfrx;

  assign                   {
                             zxgpsirnmn33k29fvgm
                           , t3ysg7mwfhqy_9hje
                           , n1lhs71oc209opa
                           } = od5a1yudx9bmyqpwleexh4h9;

  assign idw2i93am7m9wy_5hzipgymj5k3 = {
                             a_pr26ts5th7p3ziyczhdy
                           , nhafiywg3hg_52kogwh
                           , t9yh0n7ay27ft001vimu6
                           };

  wire l0_5x2ohgu6m77k54mg;

  localparam tcebpmbl7g = 0;

  ux607_gnrl_icb_arbt # (
  .ARBT_SCHEME (3),
  .ALLOW_0CYCL_RSP (0),


  .FIFO_OUTS_NUM   (8),
  .FIFO_CUT_READY  (tcebpmbl7g),
  .ARBT_NUM   (y7fi7kw8i180nr4b),
  .ARBT_PTR_W (senagm_wgrp66rwiuyf1d),
  .USR_W      (s3xvyho),
  .AW         (32),
  .DW         (64) 
  ) og6hyji4910900wl8nl(
  .arbt_active            (l0_5x2ohgu6m77k54mg )     ,

  .o_icb_cmd_valid        (ouat_m1vwjc0l5igzo2z4g )     ,
  .o_icb_cmd_ready        (gyja61p9t197hw65hvyi63g )     ,
  .o_icb_cmd_read         (mrrzsfopopzgqr_nro5 )      ,
  .o_icb_cmd_addr         (v10jhardhhvft6w6t3u )      ,
  .o_icb_cmd_wdata        (pp5egelk49dgurfb3w )     ,
  .o_icb_cmd_wmask        (n9sl3nl16qlprh9ocn6trcs)      ,
  .o_icb_cmd_burst        (g3iy6vml027o3gv9wt)     ,
  .o_icb_cmd_beat         (z0y5vk22vnz94pcxx )     ,
  .o_icb_cmd_excl         (rvqfn2hxjfeh8egdvsc )     ,
  .o_icb_cmd_lock         (l1368lp6updfhsbebtzpc )     ,
  .o_icb_cmd_size         (c55olxxsckol_k4eb9fyu )     ,
  .o_icb_cmd_usr          (jmo524gyok0abs1u1  )     ,

  .o_icb_rsp_valid        (n0wp_tjsit08gjo9ggcxe_a )     ,
  .o_icb_rsp_ready        (ebnc6trwg85shv8_iz8qpa2 )     ,
  .o_icb_rsp_err          (n93c2nog4f68lktvd0)        ,
  .o_icb_rsp_excl_ok      (uezhv2clc8f9woh7dc5ss1)    ,
  .o_icb_rsp_rdata        (j2p0ug10na1wztrfj39 )     ,
  .o_icb_rsp_usr          (guqjz9gxv28q8f719   )     ,

  .i_bus_icb_cmd_sel_vec  (ccxw7l8izxzjj14ozqkgvvyd6) ,

  .i_bus_icb_cmd_ready    (w0hjg2xow0ymilw7bcxpm2l ) ,
  .i_bus_icb_cmd_valid    (k1_j5ubhqqpfrl3p0bi186va9 ) ,
  .i_bus_icb_cmd_read     (a_dm6kd_qbw2cv84wtboltif01 )  ,
  .i_bus_icb_cmd_addr     (xzpsiztjmn62eb967x1xkc6 )  ,
  .i_bus_icb_cmd_wdata    (ae00o9ay050qc5d5zxf18282b92 ) ,
  .i_bus_icb_cmd_wmask    (puxr8jzij0m30qcwmdz2sufl51)  ,
  .i_bus_icb_cmd_burst    (sxjmcdip1m7ighns0k5aue59fj)  ,
  .i_bus_icb_cmd_beat     (noyjdh392j1x0s9g1b_lk )  ,
  .i_bus_icb_cmd_excl     (wspjbjcpf459zy17qhyz8jmqy7 )  ,
  .i_bus_icb_cmd_lock     (s6vj39lt1yt7f1ytk3pr3 )  ,
  .i_bus_icb_cmd_size     (y7jg1o7n3jl52fxr0isdv8 )  ,
  .i_bus_icb_cmd_usr      (w8o2oxw46tp1zf4rujrx4zyxw  )  ,

  .i_bus_icb_rsp_valid    (qkiytqsa_fo9x5ls7yb_x1k2 ) ,
  .i_bus_icb_rsp_ready    (idw2i93am7m9wy_5hzipgymj5k3 ) ,
  .i_bus_icb_rsp_err      (wzmdtyq65i82w_tt0juwqle)    ,
  .i_bus_icb_rsp_excl_ok  (kz10yoaxkacgm38dwv37tl2ixfv),
  .i_bus_icb_rsp_rdata    (fyvkbec2dn4rlcslyiyttfrx ) ,
  .i_bus_icb_rsp_usr      (od5a1yudx9bmyqpwleexh4h9) ,

  .clk                    (gf33atgy  ),
  .rst_n                  (ru_wi)
  );


  wire qf94s1s_bj_13_s82dlk = jmo524gyok0abs1u1[ale66u8k_50s8h4vdf4];
  wire c0cdxb8nf4_hmdmd1 = jmo524gyok0abs1u1[au8wnhbd2ozhfnnm];
  assign sw9511te5wakyzkx_xdo = jmo524gyok0abs1u1[bvma5mx5x4uqrf];
















  wire v2xw59pj55k_pw75  = t06t7flkpby01affnv56x64 & (v10jhardhhvft6w6t3u[32-1:12]  ==  r480zryu00zrqkrbk[32-1:12]);
  


  wire sroawsxne_wyc5t9omb6g = (v10jhardhhvft6w6t3u[32-1:16] ==  zys87dxafg7t5ll4o9[32-1:16]);
  wire vb7n7hs52iurv9_q6u2e = (v10jhardhhvft6w6t3u[32-1:26] ==  o4f5s69ex_fk0k7q13x[32-1:26])
                         & (sroawsxne_wyc5t9omb6g ? (~dn8riluj40uunvq5) : 1'b1);

  wire u45laizt1rdqmikfe670x8 = sroawsxne_wyc5t9omb6g & (~vb7n7hs52iurv9_q6u2e);

  wire xyky68zzrw4t0pfg = (v10jhardhhvft6w6t3u[32-1:16] ==  rqbq0wq0_ojyw61v5[32-1:16]) 
                        & (~u45laizt1rdqmikfe670x8)
                        & (~vb7n7hs52iurv9_q6u2e)
                        ;

  wire zg0b0ylwoqa1pzq5j65hk = 1'b0;

  wire c1ypfhh0xys78m38 = (v10jhardhhvft6w6t3u[32-1:20] ==  dak283_f21dou11_grfkt[32-1:20])
                        & (~xyky68zzrw4t0pfg)
                        & (~zg0b0ylwoqa1pzq5j65hk)
                        & (~u45laizt1rdqmikfe670x8)
                        & (~vb7n7hs52iurv9_q6u2e)
                        ;

  wire w1d8q0oe30kyhyhea2mkjp = ( 1'b0
                              | u45laizt1rdqmikfe670x8 
                              | vb7n7hs52iurv9_q6u2e 
                              | xyky68zzrw4t0pfg
                              | c1ypfhh0xys78m38
                              );

  wire pc2v5tjqs_vfqeytpe1bag5 = (v2xw59pj55k_pw75 | w1d8q0oe30kyhyhea2mkjp);









  wire w0cy4kal0ptfu_q6ras9 = 1'b0;

  wire dipozqx7k9625g2y = w92a5o09fp9dg6 & (v10jhardhhvft6w6t3u[32-1:16] ==  yh9n8rxd7xt9w6cyy9[32-1:16]) 
                         & (~pc2v5tjqs_vfqeytpe1bag5)
                         ;

  wire l42_x3lfhhdlhfh8 = eglor15f7p2ivpny5dc & (v10jhardhhvft6w6t3u[32-1:16] ==  r0bsza4vt3629icr[32-1:16]) 
                         & (~pc2v5tjqs_vfqeytpe1bag5)
                         & (~dipozqx7k9625g2y)
                         ;









  wire jt63n99bmn85_0e5y = 1'b0;

  wire ftduj_ksv07krso1v7qzo = ((~dipozqx7k9625g2y) & 
                              (~l42_x3lfhhdlhfh8) & 
                              (~w0cy4kal0ptfu_q6ras9) &
                              (~w1d8q0oe30kyhyhea2mkjp) &
                              (~jt63n99bmn85_0e5y) 
                             ) | v2xw59pj55k_pw75;


  wire x8500k3hem57qn56o = ouat_m1vwjc0l5igzo2z4g & gyja61p9t197hw65hvyi63g;

  wire pmsmdo76nri60l5ki = n0wp_tjsit08gjo9ggcxe_a & ebnc6trwg85shv8_iz8qpa2;



  wire x6zj3owgdax6mcbmtv5;
  wire ocjwpiw30_43eoiw7 = x8500k3hem57qn56o;
  wire qamh5ghinc961fix    = (~x6zj3owgdax6mcbmtv5);
  wire t9l7jv54spo1znips46v;
  wire xzkey22ytu89qx4rj = pmsmdo76nri60l5ki;
  wire gcakj3d_zfb_gif5obck   = (~t9l7jv54spo1znips46v);

  wire gsyk9gdmaaouvjl_mbdk;
  wire cp0pw7bsoc5xossrw8_mmy;
  wire ypafrfh_6tx3_ko9y_051b;
  wire eayxi7s4oo1wauen02a6;
  wire m6udccm1itc8_lrhm;
  wire lu_vj80qwl1wd7npuppw6;

  localparam kcxtq1kcall = (s3xvyho+6);
  wire [8-1:0] rt9r3il3zsa8jwi9hg1gkb8t = n9sl3nl16qlprh9ocn6trcs;

  wire [kcxtq1kcall-1:0] ge2aenpez66yjs20td;
  wire [kcxtq1kcall-1:0] pkz7kx2s1o0eumk;

  assign ge2aenpez66yjs20td =  {
          ftduj_ksv07krso1v7qzo,
          jt63n99bmn85_0e5y,
          w1d8q0oe30kyhyhea2mkjp,
          w0cy4kal0ptfu_q6ras9,
          dipozqx7k9625g2y,
          l42_x3lfhhdlhfh8,
          jmo524gyok0abs1u1 
          };

  assign   
      {
          gsyk9gdmaaouvjl_mbdk,
          cp0pw7bsoc5xossrw8_mmy,
          ypafrfh_6tx3_ko9y_051b,
          eayxi7s4oo1wauen02a6,
          m6udccm1itc8_lrhm,
          lu_vj80qwl1wd7npuppw6,
          s_s052pc2p3r_9o280580 
          } = pkz7kx2s1o0eumk & {kcxtq1kcall{t9l7jv54spo1znips46v}};



  assign guqjz9gxv28q8f719 = s_s052pc2p3r_9o280580;

  ux607_gnrl_fifo # (
    .CUT_READY (tcebpmbl7g),
    .MSKO      (0),
    
    .DP  (8),
    .DW  (kcxtq1kcall)
  ) g2lmqduagxiq4m8v6qmmn (
    .i_vld  (ocjwpiw30_43eoiw7),
    .i_rdy  (x6zj3owgdax6mcbmtv5),
    .i_dat  (ge2aenpez66yjs20td ),
    .o_vld  (t9l7jv54spo1znips46v),
    .o_rdy  (xzkey22ytu89qx4rj),  
    .o_dat  (pkz7kx2s1o0eumk ),  
    .clk  (gf33atgy),
    .rst_n(ru_wi)
  );
















  wire lv1gcem_88yah80x5kf = (~gcakj3d_zfb_gif5obck) & 
        (~({ftduj_ksv07krso1v7qzo, w1d8q0oe30kyhyhea2mkjp, jt63n99bmn85_0e5y, w0cy4kal0ptfu_q6ras9, dipozqx7k9625g2y, l42_x3lfhhdlhfh8}
        == {gsyk9gdmaaouvjl_mbdk, ypafrfh_6tx3_ko9y_051b, cp0pw7bsoc5xossrw8_mmy, eayxi7s4oo1wauen02a6, m6udccm1itc8_lrhm, lu_vj80qwl1wd7npuppw6}));

  wire csr6ull36_jpsgz3o2al = qf94s1s_bj_13_s82dlk ? lv1gcem_88yah80x5kf : 1'b0;


  wire x34gbidn7gdc04sv3xob7gtiyg8 = (~qamh5ghinc961fix) & (~csr6ull36_jpsgz3o2al);
  wire s0dndzoayazaep13ud5wy8_miu7;

  wire u3812fgbq7igezs8_j_umg5lzx = x34gbidn7gdc04sv3xob7gtiyg8 & ouat_m1vwjc0l5igzo2z4g;
  assign gyja61p9t197hw65hvyi63g     = x34gbidn7gdc04sv3xob7gtiyg8 & s0dndzoayazaep13ud5wy8_miu7;

  wire tnol4dhc571tkxhbu;
  wire edca7mfhfghe2olz2pb5yxyg093xy4;
  wire n658pzyddgw113gth7puctgz6ajb82g_2;
  wire ekmsh07qax_1w3x07vrccw_ftm941;
  wire kkxaswsip67h0jf4nu1xi2feika6d;
  wire ekxmo4ahsqfwqjhg6mytoug_gm3j7mzp;
  wire poo39net46fse3ohh15meqrxmkk;
  wire qwe3beh7gwnvqjd0sg1jglxn63xrit;

  assign k5t515v6aa4oilq98cy6lrd8 = u3812fgbq7igezs8_j_umg5lzx & ftduj_ksv07krso1v7qzo & n658pzyddgw113gth7puctgz6ajb82g_2;
  assign nbgnnsuqy2oogaz89vmbl1 = sw9511te5wakyzkx_xdo; 
  assign c1_3zcfvbhkc9cf7jgm7x  = v10jhardhhvft6w6t3u ; 
  assign cki2l53v3p6py9awsecgj = k8aii0cb2ywh7xvp5ud9; 
  assign ddjl2wsfh12b286nsrl3m5z = vyaut44yc_lmxpxuhm; 
  assign y09wfhff_yx31yoe7cxv = t06t7flkpby01affnv56x64; 
  assign sk43hkjk_z2mer7becad  = mrrzsfopopzgqr_nro5 ; 
  assign zn80vi7_hafilb62kh72jx5d6= qf94s1s_bj_13_s82dlk ; 
  assign e1wmvmyg_x8tobsfzpo    = c0cdxb8nf4_hmdmd1 ; 
  assign lo0fo8wk5o04f7ezwv474 = pp5egelk49dgurfb3w;
  assign zutoko8hik1j9pa64jmpuw = rt9r3il3zsa8jwi9hg1gkb8t;
  assign xqdmvgffpmzj6n0l23o  = l1368lp6updfhsbebtzpc ;
  assign of_yab2i0nf9xv_tek5r  = rvqfn2hxjfeh8egdvsc ;
  assign i1pzsd21aml3amhex3sf  = c55olxxsckol_k4eb9fyu ;















  assign hr7la0400ty0hiwk5d0 = u3812fgbq7igezs8_j_umg5lzx & w1d8q0oe30kyhyhea2mkjp & kkxaswsip67h0jf4nu1xi2feika6d;
  assign lqv5bv6hq78ov_prb97v5z  = v10jhardhhvft6w6t3u;
  assign o15lm7no18top00l32ra = k8aii0cb2ywh7xvp5ud9; 
  assign ly1y__c5rzaa9xv_9_m1ppr = vyaut44yc_lmxpxuhm; 
  assign f1msmreidlchd7rf9w625 = t06t7flkpby01affnv56x64; 
  assign uarhtvlb5te5hc2g3  = mrrzsfopopzgqr_nro5 ; 
  assign g9ayxf51lhjl44vvw62u3 = pp5egelk49dgurfb3w;
  assign qfoijjxktg6dht3klxhyw5g = rt9r3il3zsa8jwi9hg1gkb8t;
  assign gao2lzva86gawlwp2  = l1368lp6updfhsbebtzpc ;
  assign xpt7vgmhw7tamcpv2l  = rvqfn2hxjfeh8egdvsc ;
  assign lrh4lctjvrz1rhm6b9oh  = c55olxxsckol_k4eb9fyu ;
  assign pyfc_rgr3cwwvo34pf   = xyky68zzrw4t0pfg;
  assign u6xj18ku9lj1890n7  = u45laizt1rdqmikfe670x8;
  assign s3lwpy5def9adgbbvx9ct  = vb7n7hs52iurv9_q6u2e;
  assign q96vjidg4x6ohxl7   = zg0b0ylwoqa1pzq5j65hk;
  assign krh62hs2scfnb76m67a   = c1ypfhh0xys78m38;


  assign tw0yf9aln_vu06k8l = u3812fgbq7igezs8_j_umg5lzx & dipozqx7k9625g2y & poo39net46fse3ohh15meqrxmkk;
  assign ss4cm882613f24kdjqsyl  = v10jhardhhvft6w6t3u [16-1:0]; 
  assign zm9uosdggg7ntkh97elw = k8aii0cb2ywh7xvp5ud9; 
  assign g_ahl2zik6mj75atnp_hej = vyaut44yc_lmxpxuhm; 
  assign bjl40q8m35dwdn_mn9 = t06t7flkpby01affnv56x64; 
  assign oefdpb9h9kx627r_0y5  = mrrzsfopopzgqr_nro5 ; 
  assign fh1jm1za5zvqmvdloi = pp5egelk49dgurfb3w;
  assign sp_0hv_ae5rrl9vagusi = rt9r3il3zsa8jwi9hg1gkb8t;
  assign b4oh48a9a0g269ybrm  = l1368lp6updfhsbebtzpc ;
  assign r5s3ykb7_xkl6t12oucf  = rvqfn2hxjfeh8egdvsc ;
  assign ssswxj_bpfx_ebsbj  = c55olxxsckol_k4eb9fyu ;

  assign rqf8b5xxbw0n1_qaw = u3812fgbq7igezs8_j_umg5lzx & l42_x3lfhhdlhfh8 & qwe3beh7gwnvqjd0sg1jglxn63xrit;
  assign holgl43_yucp7f7l  = v10jhardhhvft6w6t3u [16-1:0]; 
  assign oyev1ipmdflkvxygwr = k8aii0cb2ywh7xvp5ud9; 
  assign ihknw7_lm_572tv6s = vyaut44yc_lmxpxuhm; 
  assign o31l03k34sdhwt4lkazfa5 = t06t7flkpby01affnv56x64; 
  assign gy2sgn_1bpkac7msq3  = mrrzsfopopzgqr_nro5 ; 
  assign r_1u6q2lzkfus3o9nfl = pp5egelk49dgurfb3w;
  assign yff7wf8wth2vjkdjpr = rt9r3il3zsa8jwi9hg1gkb8t;
  assign lppjhpov_5lgvx7n7fm4g  = l1368lp6updfhsbebtzpc ;
  assign sdfg9zykj79rz_7thf9k  = rvqfn2hxjfeh8egdvsc ;
  assign wt4e4tlh0u_4cljr2j5f9  = c55olxxsckol_k4eb9fyu ;









  assign y1rlahaedj99shvl6uc = (|ccxw7l8izxzjj14ozqkgvvyd6);
  assign c0x_72w8ddbpt17fn = (|ccxw7l8izxzjj14ozqkgvvyd6) & dipozqx7k9625g2y;



























  assign tnol4dhc571tkxhbu =  
            (lkdpdaxvpxpy8w8hpchiph) 
          & (y1ipzdhzcfq282ups6ja) 
          & (q84eo09gg53r2jj5a5xn) 
          & (ocwcf75wgxfb1bawe) 
             ;

  assign edca7mfhfghe2olz2pb5yxyg093xy4 =  
            1'b1
          & (lkdpdaxvpxpy8w8hpchiph) 
          & (y1ipzdhzcfq282ups6ja) 
          & (q84eo09gg53r2jj5a5xn) 
          & (ocwcf75wgxfb1bawe) 
             ;

  assign n658pzyddgw113gth7puctgz6ajb82g_2 =  
            1'b1
          & (y1ipzdhzcfq282ups6ja) 
          & (q84eo09gg53r2jj5a5xn) 
          & (ocwcf75wgxfb1bawe) 
             ;
  assign ekmsh07qax_1w3x07vrccw_ftm941 =  
            (lkdpdaxvpxpy8w8hpchiph) 
          & (y1ipzdhzcfq282ups6ja) 
          & (q84eo09gg53r2jj5a5xn) 
          & (ocwcf75wgxfb1bawe) 
             ;

 assign kkxaswsip67h0jf4nu1xi2feika6d =  
            (lkdpdaxvpxpy8w8hpchiph) 
          & 1'b1
          & (q84eo09gg53r2jj5a5xn) 
          & (ocwcf75wgxfb1bawe) 
             ;

 assign ekxmo4ahsqfwqjhg6mytoug_gm3j7mzp =  
            (lkdpdaxvpxpy8w8hpchiph) 
          & (y1ipzdhzcfq282ups6ja) 
          & (q84eo09gg53r2jj5a5xn) 
          & (ocwcf75wgxfb1bawe) 
             ;

 assign poo39net46fse3ohh15meqrxmkk =  
            (lkdpdaxvpxpy8w8hpchiph) 
          & (y1ipzdhzcfq282ups6ja) 
          & 1'b1
          & (ocwcf75wgxfb1bawe) 
             ;

 assign qwe3beh7gwnvqjd0sg1jglxn63xrit =  
            (lkdpdaxvpxpy8w8hpchiph) 
          & (y1ipzdhzcfq282ups6ja) 
          & (q84eo09gg53r2jj5a5xn) 
          & 1'b1
             ;


  assign s0dndzoayazaep13ud5wy8_miu7 = tnol4dhc571tkxhbu;  



  localparam mp26klefy4v2f = (2+64);
  wire [mp26klefy4v2f-1:0] i2pk7kg6dmy2u8yk = {
                                 l8ymtznl9hcobcfqg,
                                 ybmlc9yctmeh5ymbek57,
                                 z4lyw1_nvshizqbim5x  
                                 };

  wire [mp26klefy4v2f-1:0] pq28r_0p1z8tuc;

  assign {
                                 n93c2nog4f68lktvd0,
                                 uezhv2clc8f9woh7dc5ss1,
                                 j2p0ug10na1wztrfj39  
                                 } = pq28r_0p1z8tuc;

  ux607_gnrl_bypbuf # (
    .DP  (1),
    .DW  (mp26klefy4v2f)
  ) vd71zpjbwqqln4dju_sreu8cz7 (
    .i_vld(qywrqdqbkmyeridmga5k),
    .i_rdy(ya7at6mg3adjqzbi1c6),
    .i_dat(i2pk7kg6dmy2u8yk ),
    .o_vld(n0wp_tjsit08gjo9ggcxe_a),
    .o_rdy(ebnc6trwg85shv8_iz8qpa2),  
    .o_dat(pq28r_0p1z8tuc ),  
  
    .clk  (gf33atgy),
    .rst_n(ru_wi)
  );








  assign {
          qywrqdqbkmyeridmga5k 
        , l8ymtznl9hcobcfqg 
        , ybmlc9yctmeh5ymbek57 
        , z4lyw1_nvshizqbim5x 
         } =
            ({64+3{gsyk9gdmaaouvjl_mbdk}} &
                        { ltzq1n1rg2b9lrt8j0bs__wa 
                        , qf_hxpj8b9rdyabqx8q7l 
                        , pqfnz7dk2f2khe5zxq0081lzv 
                        , j3gop6yag94s712e_mipwr484 
                        }
            ) 
          | ({64+3{ypafrfh_6tx3_ko9y_051b}} &
                        { b6m1vcd7bmemxnu99_zke 
                        , jpa5gwkjwqz_j0a3cy1 
                        , kjxe2fpsacp9bx2_0fah36ij 
                        , xsw8oz2ni13z6vac1tn61 
                        }
            ) 
          | ({64+3{m6udccm1itc8_lrhm}} &
                        { fsj22rallxmhdrvuwenpq 
                        , hhlfu4md9k5v7naf1qt 
                        , j8m9s_du9fk99idlbh80 
                        , aapsfpke41r7dyya4ah 
                        }
            ) 
          | ({64+3{lu_vj80qwl1wd7npuppw6}} &
                        { o4wuryrcvw13y2v5m6b6u 
                        , vnqegbzme0jutvf 
                        , jdj122rbumyogtin6xpg97 
                        , p9mcc6npaw32uigcp6 
                        }
            ) 
             ;

  assign qui4zelf64bknwchxnz6 = gsyk9gdmaaouvjl_mbdk & ya7at6mg3adjqzbi1c6;
  assign vqld30a8qt13mzhwoc   = ypafrfh_6tx3_ko9y_051b   & ya7at6mg3adjqzbi1c6;
  assign yign8d_dhrow0i5wjts4bd   = m6udccm1itc8_lrhm   & ya7at6mg3adjqzbi1c6;
  assign bt4howrm5xnf6u4fuwrum6   = lu_vj80qwl1wd7npuppw6   & ya7at6mg3adjqzbi1c6;




  assign o4qff84vfbn       = c0l6w8lh_td7pzkcpdfp0ir_t & (~gt923cnjxl9zc1kavj6ay3l6vo6);
  assign flcopog5zzpohfautwy = c0l6w8lh_td7pzkcpdfp0ir_t &   gt923cnjxl9zc1kavj6ay3l6vo6;

  assign a_pr26ts5th7p3ziyczhdy =
      gt923cnjxl9zc1kavj6ay3l6vo6 ?  gtb8f_h0g28itdr8k : x74_jhmpouk; 

  assign wf15djwi2hw25nz_   = r22ymekw52k08rw4tm0  ;
  assign t1q5qmk9jzpf6glng4y = zdg2ytmoa2dqi_9xntu0hld3fx  ;
  assign xsmx4zoewhbt07jxq = wsxqohy8uxi3mw1ruq9o5z2;

  assign l8ng5e_pa1fg07__37   = uyma7dg_jtxevl8vmljt;


  assign ytp8_jsqr2sjmu08gdn = 5'b0;


  wire  afxrizdnkg3         = bzjsole_y2xxo6diyfseg;






















  wire c5oh1h2z = (nxjbs9v14ld33363ewcmdo1 == 2'b00) & (y3cb9jdvssvccg6b1mqbt7jl_ == 1'b1);
  wire nfljtz5q  = (nxjbs9v14ld33363ewcmdo1 == 2'b00) & (y3cb9jdvssvccg6b1mqbt7jl_ == 1'b0);
  wire e3pjnc5fbdsc = (nxjbs9v14ld33363ewcmdo1 == 2'b01) & (y3cb9jdvssvccg6b1mqbt7jl_ == 1'b1);
  wire wath3r5wcu  = (nxjbs9v14ld33363ewcmdo1 == 2'b01) & (y3cb9jdvssvccg6b1mqbt7jl_ == 1'b0);
  wire lx2n9_iy = (nxjbs9v14ld33363ewcmdo1 == 2'b10) & (y3cb9jdvssvccg6b1mqbt7jl_ == 1'b1);
  wire hi_tkvoa  = (nxjbs9v14ld33363ewcmdo1 == 2'b10) & (y3cb9jdvssvccg6b1mqbt7jl_ == 1'b0) 
                   & (~afxrizdnkg3) 
                 ;
    wire f2_q9t25qj  = (nxjbs9v14ld33363ewcmdo1 == 2'b10) & (y3cb9jdvssvccg6b1mqbt7jl_ == 1'b0) & afxrizdnkg3;
  wire v3kxw7  = (nxjbs9v14ld33363ewcmdo1 == 2'b11);

  wire [64-1:0] qo6_c4yxtkeo = 
      (wsxqohy8uxi3mw1ruq9o5z2 >> {jqxmjq8am07ckn333alfaky1b[2:0],3'b0});

  assign z5tnbveujliw633sxlb8   = 
            ({64{c5oh1h2z}} & {{64- 8{          1'b0}}, qo6_c4yxtkeo[ 7:0]})
          | ({64{nfljtz5q }} & {{64- 8{qo6_c4yxtkeo[ 7]}}, qo6_c4yxtkeo[ 7:0]})
          | ({64{e3pjnc5fbdsc}} & {{64-16{          1'b0}}, qo6_c4yxtkeo[15:0]})
          | ({64{wath3r5wcu }} & {{64-16{qo6_c4yxtkeo[15]}}, qo6_c4yxtkeo[15:0]}) 
          | ({64{lx2n9_iy}} & {{64-32{          1'b0}}, qo6_c4yxtkeo[31:0]}) 
          | ({64{hi_tkvoa }} & {{64-32{qo6_c4yxtkeo[31]}}, qo6_c4yxtkeo[31:0]}) 
          | ({64{f2_q9t25qj}} & {{32{1'b1}}, qo6_c4yxtkeo[31:0]})
          | ({64{v3kxw7 }} & qo6_c4yxtkeo[63:0])  
          ;




























  assign erdoc9bbdnq8065yw    = r22ymekw52k08rw4tm0;
  assign ro93aearv5754gz9w  = r22ymekw52k08rw4tm0;
  assign y9389ymcyh2ia2082yx1_ = {{64-32{1'b0}},jqxmjq8am07ckn333alfaky1b};
  assign uiu4_g7j41kz      = 64'b0;
  assign zqx1cj9lvt0e      =  gx8_jfgud1t_azz9c19jh;
  assign zsxgccndqw2suf6      = ~gx8_jfgud1t_azz9c19jh;



  assign bhjn0b8ydp0vfsiy = (|ccxw7l8izxzjj14ozqkgvvyd6) | t9l7jv54spo1znips46v | l0_5x2ohgu6m77k54mg;

endmodule



















module dkh50cge16y( 

  input  rm1dxjejhq7dh3q5m,
  input sxvvsxtbhyvt,

  input [8*32-1:0] pcr4upio7_tx37, 
  input [8*1-1:0] uzklqlncpqqm1rav,
  input [8*1-1:0] ortueunvnkx_l5m_j,
  input [8*1-1:0] hwuhtb7ucto_utk56,
  input [8*2-1:0] i1env2kmns7qvvuuc,
  input [8*1-1:0] g3s3vpafvy3i,
  input  rvr30vvllni,



  input dn8riluj40uunvq5,
  input w92a5o09fp9dg6, 
  input eglor15f7p2ivpny5dc, 


  input  qo5p9t6s74zxpo,
  output umnrzb6pv8dzc,








  output o4qff84vfbn, 
  input  x74_jhmpouk, 
  output [64-1:0] z5tnbveujliw633sxlb8,
  output [4 -1:0] l8ng5e_pa1fg07__37,
  output erdoc9bbdnq8065yw , 
  output zqx1cj9lvt0e,
  output zsxgccndqw2suf6,
  output [64 -1:0] y9389ymcyh2ia2082yx1_,
  output [64 -1:0] uiu4_g7j41kz,
  output ro93aearv5754gz9w , 
  output rqy9v1_k_o74etonfc , 
  output [4:0] ytp8_jsqr2sjmu08gdn,

  output                         flcopog5zzpohfautwy, 
  input                          gtb8f_h0g28itdr8k, 
  output                         wf15djwi2hw25nz_  , 
  output                         t1q5qmk9jzpf6glng4y,
  output [64-1:0]      xsmx4zoewhbt07jxq,




  input                          o21b8ypt1xiu5ml63d,

  input                          badsf4ksbp3k6p_p5hnj2i, 
  input                          vrsqde4muadsevgpemk, 
  output                         ed4kcy8s9nrisftgx_q, 
  input  [32-1:0]   bdqo1tgw2_bpi2e8alini, 
  input                          jp5nha2l14e7kx2jzpke,   
  input                          za9xg3zsqni_aeqmke,   
  input                          c1gmncmorg16sachdas,   
  input                          p648zxn2luyxy8mt992a, 
  input                          uxlldm0w_h7kicit8gvhqv2, 
  input                         yvu98r_7ji4o250r_u,
  input                          zdpamqgv7ddf1n3x5t2q, 
  input                          wpsukhyqhl92dzoam7cm, 
  input                          v3oo69y614hgiemyyld,

  input  [64-1:0]        a4a48egkdkec8d9b_9, 
  input  [8-1:0]      xwfmltfzahuj4qfn4qf2, 
  input  [1:0]                   ggxoqcj7ytp1a4pjf7ee,
  input                          l3c127qdc9a2mfc13,
  input  [4 -1:0] oq9b5zfhza9yvdoj,
  input                          sg33s7pt45jp_,
  input                          g9i9mf8jq7sc699j,
  input  [4:0]                   szrgf24or2mbt7w_yleh_vt,

  input  yixt0a_xmh    ,
  input  fgnb7mhn1254le9     ,
  input  okt7c24tca9ji6pw     ,


  
  
  
  
  input                          fkm9up63o1aeauaqhjb,
  output                         to_1lv9wnb3vmu6tvz5rc,
  input  [32-1:0]   ju1kbeplcqy314lfj4, 
  input                          r985fbe5k7hgzaq9i, 
  input                          bb04gpwotp2s6c7_p1gqkq, 
  input                          sqmey185cu3mtixhl, 
  input                          rffcsd1o699ytclmx,
  input  [64-1:0]        lbr88vbqtg8rht7320frde,
  input  [8-1:0]     g7qq38mx3d58n1b15kcia,
  input                          demg_fwfkmaeawq30t,
  input                          grtb6ypa0px2gi1c,
  input  [1:0]                   f128d8ws0seoihu1,
  
  output                         m2r7mfmq3afdd1ine,
  input                          nhafiywg3hg_52kogwh,
  output                         xrqayy6vigrw66z8a  ,
  output                         jyy72ywt9nbo10f2jxupacld,
  output [64-1:0]        drz92qecqx_qtxwro,

  
  
  
  
  input                          cxrbvs1hde7j8ziudd4ar,
  output                         dmzxpdd5dgmp_2ip6h3_6,
  input  [32-1:0]     piv1ndd8n8dlaqx9, 
  input                          r3rgwuaokuw68zin, 
  input                          m2aue5rcrjkbzdwbqvlzvr, 
  input                          u7a8_cbg_zi4w4b4slc08, 
  input                          fd_1f891ni339pnyzw63mg,
  input  [64-1:0]      p1g5jbgswdsx9v1j01103,
  input  [8-1:0]      zmrmpw_9vyme3rakn8br8e,
  input                          sp2wnouu73ujsanhkn0,
  input                          n5w05rcecv47nvnfkkw5,
  input  [1:0]                   dycy3iz66xw6yj5ea,
  input                          wic6t212ob4tfa,
  input                          zqnzorh6g9hnwsot5zr,
  
  output                         ro76scx3ggmfi4xp2bjx,
  input                          t9yh0n7ay27ft001vimu6,
  output                         gpjxeoxkmf35ldn  ,
  output                         owde01ai01h2x5kn3_ng,
  output [64-1:0]      atur2zwqwk4mnbtz68l2,




  
  
  
  
  output                         c0x_72w8ddbpt17fn,
  
  output                         tw0yf9aln_vu06k8l,
  input                          q84eo09gg53r2jj5a5xn,
  output [16-1:0]   ss4cm882613f24kdjqsyl, 
  output                         zm9uosdggg7ntkh97elw, 
  output                         g_ahl2zik6mj75atnp_hej, 
  output                         bjl40q8m35dwdn_mn9,
  output                         oefdpb9h9kx627r_0y5, 
  output [64-1:0]        fh1jm1za5zvqmvdloi,
  output [8-1:0]      sp_0hv_ae5rrl9vagusi,
  output                         b4oh48a9a0g269ybrm,
  output                         r5s3ykb7_xkl6t12oucf,
  output [1:0]                   ssswxj_bpfx_ebsbj,
  
  
  input                          fsj22rallxmhdrvuwenpq,
  output                         yign8d_dhrow0i5wjts4bd,
  input                          hhlfu4md9k5v7naf1qt  ,
  input                          j8m9s_du9fk99idlbh80  ,
  input  [64-1:0]        aapsfpke41r7dyya4ah,

  
  
  
  output                         y1rlahaedj99shvl6uc,
  
  
  output                         rqf8b5xxbw0n1_qaw,
  input                          ocwcf75wgxfb1bawe,
  output [16-1:0]   holgl43_yucp7f7l, 
  output                         oyev1ipmdflkvxygwr, 
  output                         ihknw7_lm_572tv6s, 
  output                         o31l03k34sdhwt4lkazfa5,
  output                         gy2sgn_1bpkac7msq3, 
  output [64-1:0]        r_1u6q2lzkfus3o9nfl,
  output [8-1:0]      yff7wf8wth2vjkdjpr,
  output                         lppjhpov_5lgvx7n7fm4g,
  output                         sdfg9zykj79rz_7thf9k,
  output [1:0]                   wt4e4tlh0u_4cljr2j5f9,
  
  
  input                          o4wuryrcvw13y2v5m6b6u,
  output                         bt4howrm5xnf6u4fuwrum6,
  input                          vnqegbzme0jutvf  ,
  input                          jdj122rbumyogtin6xpg97  ,
  input  [64-1:0]        p9mcc6npaw32uigcp6,


  
  
  
  
  
  output                         hr7la0400ty0hiwk5d0,
  input                          y1ipzdhzcfq282ups6ja,
  output [32-1:0]   lqv5bv6hq78ov_prb97v5z, 
  output                         o15lm7no18top00l32ra, 
  output                         ly1y__c5rzaa9xv_9_m1ppr, 
  output                         f1msmreidlchd7rf9w625,
  output                         uarhtvlb5te5hc2g3, 
  output [32-1:0]        g9ayxf51lhjl44vvw62u3,
  output [4-1:0]      qfoijjxktg6dht3klxhyw5g,
  output                         gao2lzva86gawlwp2,
  output                         xpt7vgmhw7tamcpv2l,
  output [1:0]                   lrh4lctjvrz1rhm6b9oh,
  output                         krh62hs2scfnb76m67a,
  output                         pyfc_rgr3cwwvo34pf,
  output                         u6xj18ku9lj1890n7,
  output                         s3lwpy5def9adgbbvx9ct,
  output                         q96vjidg4x6ohxl7,
  
  
  input                          b6m1vcd7bmemxnu99_zke,
  output                         vqld30a8qt13mzhwoc,
  input                          jpa5gwkjwqz_j0a3cy1  ,
  input                          kjxe2fpsacp9bx2_0fah36ij  ,
  input  [32-1:0]        xsw8oz2ni13z6vac1tn61,








  output                         cv0k9k_ijjnnylw1s7b_0d,

  output                         swpk4h0gei3t_34xogbqncbo4,

  input                          u9qmfl3rwx0dhr92z875vx7q,
  output [32-1:0]   unu_x_i6jmr33nz0yitzk, 
  output                         ngyxf4n1cpcgks_s2zmgfb260, 
  output                         c7m50uaw8lmp_iv4ci38q2, 
  output                         m04a1mtbabwezldp1crh4rg6z,
  output                         hwjq1ubtaei44lpk609fm2hb8,
  output                         e28p_fu1k484ncul0p85ko,
  output                         bei3qhdtd0euq2emblogsu_x, 
  output [64-1:0]        bf0_ynb648lqi7s93eieo0ln,
  output [8-1:0]     wf8o7p9_qfthhoxs747wyeuwkky,
  output  [2:0]                  ygro7xue7x7rtdafkj3o4q4,
  output  [1:0]                  drrly3q0ocg8d4pwh3m9o77,
  output                         g654a6a9cesbee7xs6_uu9lu5,
  output                         x7fex0jf9da6a5v1c28upl72t,
  output [1:0]                   ege0_1ufqm8i68zo4il6cwe46d,


  input                          bvg_3t_ujbpur7b_h7f63jse,

  output                         m5l6wu3uz_jfqasz8e3tsvrm,
  input                          g9so28ythfl0q7xnk66p1  ,
  input                          e66wluxk71p2ldu3a1qk994bq  ,
  input  [64-1:0]        ig2roj0y08x8_ntp3knz9rd,


  output                         a0_d_zdz9h9fgk46e8arf,

  output                         twr9y24wxhs3qj2z9f2hzpaig6,

  input                          w8b46r9cof57xvd5zo1u4zh8,
  output [32-1:0]   wn1l4cmih7rwce1rb7wk3f9wy, 
  output                         xo6ciibewn8p8xey97jcsqi5, 
  output                         evz1w_girwszyfnlcg4mwvtjo, 
  output                         ju5f9fb1erjep_bv8gpfn6,
  output                         hadi1_f3quoaotjv5758x8kksot2,
  output                         bdi4gjlb0po4ejcztowoqil7,
  output                         cgnzbuo_1yz6v42seb25duv, 
  output [64-1:0]        zopev7f487spn9mwvuowqo,
  output [8-1:0]     p32jk0lb8g31kqlpvmllo75qim,
  output  [2:0]                  g973rcaou05i456suvk_89dm,
  output  [1:0]                  wflv6rhfdwyxttak111v1l,
  output                         ggsmt4nzx8pwlowehinqvk60f,
  output                         xu8494ii8ectqb91224uuer,
  output [1:0]                   r6rk128ijo839ougen9stbe,


  input                          m7tq_t57mr5bovbb9ghffl4k,

  output                         gpcgdcri3e6_fxrw8wwtysoqqr,
  input                          a6s4kxg1ibr6mntc85jik  ,
  input                          hizzalmpwr8cqkxqi80wvbt65x  ,


  
  output                          p7ah58va5_2njbtv, 
  output [64-1:0]         u981qrwkgi5h0e72b__gg19w,  
  output                          p0i2i3v3j1tclelx51,
  
  output                          mum8f1rtatle7p_55y84,  
  output [6-1:0]  pn5bpwlp5ijfako9m5ao,
  output                          g3s0qe2adsxsx8e6z ,
  output [24-1:0]  a1rl4lmhqp8ydyk07kqkn,          
  input  [24-1:0]  apnns9jlj7y3y5bg8ynz,
   
  output                          pmz7e4mgvbnmimqp0nghk,  
  output [6-1:0]  j61algpxjoycxbswhgsuf, 
  output                          omq1ehm8hp4q9jgp5n5vn ,
  output [24-1:0]  fbv1q6sraswzp91zcn,          
  input  [24-1:0]  jv8kv41vzuir6an4iod,


  
  
  output                          qgl4363n31jx6xjyo05zkn,  
  output [8-1:0] zec78nyllxlfwmpsgncluudf, 
  output [4-1:0] dwvnjl0vxqkgd8t6dtvg5z,
  output [32-1:0] gngmcj5c1jd85csel9ntru,          
  input  [32-1:0] tkt93y5lfluzkia5plvksp,
                                                
  output                          km7co8hqm563od8ga_03_g,  
  output [8-1:0] j4mas6g26o63wvnsdquh8c4p, 
  output [4-1:0] nniah5mh0cunkhyln9,
  output [32-1:0] rcy_v3911lf33nza5j,          
  input  [32-1:0] g4nfgu53_rgc0632w8z97,
                                                
  output                          xzgkclcxsgfuseg87,  
  output [8-1:0] djwlah5bo0r6myit6cal0t, 
  output [4-1:0] qu_ju3lv6nvkdbo8h11uf,
  output [32-1:0] dydwz9i6k80alqfarffop,          
  input  [32-1:0] ql1c7hzoj9kf__7r97krm,
                                                
  output                          kp2j8kv1p1cjcg0lerwm,  
  output [8-1:0] v4a7g1wh3ivw0esp7dye0oiz, 
  output [4-1:0] x9zuk21gpaj58uszvm5,
  output [32-1:0] n_h5oz0c5bo5rpevwjcu8,          
  input  [32-1:0] ryid4_99ns1jc83at_88x,


  input 			              tia1md5dyh6kj4,
  input				              c4ughu0qm5sfai,
  input  			              indfp6mwqdqamez0mex,

  output 			              r5hpbriny8m67sv9e_ylgo1,
  output 			              dyl5g2vgrvy4mb3,
  input                           viuu21jzrv,


  input                          y3iin4ygz2ed73_84l91h73,
  input                          n8mvs5sw2pw48loob7jv6nmjdds,
  input                          dbzz2cu7abqy43de_ky433v,
  input                          gbb0bfnz8wqnjr5sufoh6ojt4pr,
  output                         im70q80i1xh1y_5mo9ndr1,

  input                          mmludd_fnt2yevok8a1a0 ,
  output                         buwj9_8l8bwj80kkinq9p ,

  
  input                                    ysnexkrvlg2s55ajc5g69tm,           
  input  [74-1:0]       p7832rg37bbm7_ssxunhcj7,          
  output                                   t1xtkdoie_8djygqlt1br56pwt,         
  output                                   w33zvryieg8hhgy58581ny437h9,           
  output                                   lv96t6re1w44borcb7do83ndua3vjy,           

  input  gf33atgy,
  input  ru_wi
  );



  wire                         ddl6fq6uyoan19ad7k1e7x6ut;
  wire                         tzjgmrua9xx8r7mtesjlse7ck;
  wire [32-1:0]   k3d3baof2jykxvcnolt; 
  wire                         sndcaz3jnaw0hhh4h34z; 
  wire                         e1ta255hq9y7b1vjvfw39tn9; 
  wire                         ohegnxg1amg08qiwv7ye;
  wire                         bkvescuebx122g6u90z; 
  wire [64-1:0]        ur2ihqhfmkb_slea1h731;
  wire [8-1:0]     r9qbbve4migk8rthusrhs;
  wire                         py08fct30wgf6i2wybxotxxp;
  wire                         yih871wxqwew7vzte1vz;
  wire [1:0]                   ryikyr7mft0ec23vkfx4hc;
  wire                         mtz1ahcj94t_b5n0lwt2np4;
  wire                         g4vv6e5kk3lia0_ykb0v;
  wire                         orf3s90mdtxy8zht0g8;
  wire                         blm6y03yzi8xj45jwfzaz_;
  wire                         ddxbzfgl56dmh0jni2473;
  wire                         yjy7mmnik6nbv0bv7fmw_;
  wire                         xlge7190nk7ecqh4flp7qwsxu;
  wire                         p7fyv9jmvb0qm4ay6qip;
  wire                         cyx_m80vjtb60akb9qxolqxs;
  wire [64-1:0]        si3z5gtgqu6i6mr6lop_s0g1;









  wire                          k5t515v6aa4oilq98cy6lrd8;
  wire                          nbgnnsuqy2oogaz89vmbl1;
  wire                          lkdpdaxvpxpy8w8hpchiph;
  wire  [32-1:0]   c1_3zcfvbhkc9cf7jgm7x; 
  wire                          cki2l53v3p6py9awsecgj; 
  wire                          ddjl2wsfh12b286nsrl3m5z; 
  wire                          y09wfhff_yx31yoe7cxv;
  wire                          zn80vi7_hafilb62kh72jx5d6;
  wire                          e1wmvmyg_x8tobsfzpo;
  wire                          sk43hkjk_z2mer7becad; 
  wire  [64-1:0]        lo0fo8wk5o04f7ezwv474;
  wire  [8-1:0]     zutoko8hik1j9pa64jmpuw;
  wire                          xqdmvgffpmzj6n0l23o;
  wire                          of_yab2i0nf9xv_tek5r;
  wire  [1:0]                   i1pzsd21aml3amhex3sf;


  wire                          ltzq1n1rg2b9lrt8j0bs__wa;
  wire                          qui4zelf64bknwchxnz6;
  wire                          qf_hxpj8b9rdyabqx8q7l  ;
  wire                          pqfnz7dk2f2khe5zxq0081lzv  ;
  wire  [64-1:0]        j3gop6yag94s712e_mipwr484;


  wire r29wk2o3a027n0g, smuejl3ftpm3mb2zgxm3;

  wire bhjn0b8ydp0vfsiy;

  wire [32-1:0] yh9n8rxd7xt9w6cyy9 = 32'h80000000;
  wire [32-1:0] r0bsza4vt3629icr = 32'h90000000;


  upb8yfyhriv8e c7sivq_4mtaa_pgt(
    .dn8riluj40uunvq5         (dn8riluj40uunvq5),
    .w92a5o09fp9dg6        (w92a5o09fp9dg6), 
    .eglor15f7p2ivpny5dc        (eglor15f7p2ivpny5dc), 


    .bhjn0b8ydp0vfsiy       (bhjn0b8ydp0vfsiy),
    .yh9n8rxd7xt9w6cyy9     (yh9n8rxd7xt9w6cyy9),
    .r0bsza4vt3629icr     (r0bsza4vt3629icr),

    .o4qff84vfbn           (o4qff84vfbn ),
    .x74_jhmpouk           (x74_jhmpouk ),
    .z5tnbveujliw633sxlb8       (z5tnbveujliw633sxlb8),
    .l8ng5e_pa1fg07__37       (l8ng5e_pa1fg07__37),
    .erdoc9bbdnq8065yw        (erdoc9bbdnq8065yw  ),
    .ro93aearv5754gz9w      (ro93aearv5754gz9w  ),
    .y9389ymcyh2ia2082yx1_     (y9389ymcyh2ia2082yx1_ ),
    .uiu4_g7j41kz          (uiu4_g7j41kz      ),
    .zqx1cj9lvt0e          (zqx1cj9lvt0e ),
    .zsxgccndqw2suf6          (zsxgccndqw2suf6 ),
    .ytp8_jsqr2sjmu08gdn      (ytp8_jsqr2sjmu08gdn ),

    .qzarx9bid_hex85cnt     (yixt0a_xmh             ),
    .wg5jouh0rdnsnk8kgtlq      (fgnb7mhn1254le9         ),
    .i0o9d6dhf5giw4uln5c      (okt7c24tca9ji6pw         ),
    .o21b8ypt1xiu5ml63d       (o21b8ypt1xiu5ml63d ),

    .badsf4ksbp3k6p_p5hnj2i     (badsf4ksbp3k6p_p5hnj2i ),
    .vrsqde4muadsevgpemk     (vrsqde4muadsevgpemk ),
    .ed4kcy8s9nrisftgx_q     (ed4kcy8s9nrisftgx_q ),
    .bdqo1tgw2_bpi2e8alini      (bdqo1tgw2_bpi2e8alini ),
    .uxlldm0w_h7kicit8gvhqv2    (uxlldm0w_h7kicit8gvhqv2), 
    .yvu98r_7ji4o250r_u      (yvu98r_7ji4o250r_u      ),
    .zdpamqgv7ddf1n3x5t2q     (zdpamqgv7ddf1n3x5t2q), 
    .wpsukhyqhl92dzoam7cm     (wpsukhyqhl92dzoam7cm), 
    .v3oo69y614hgiemyyld     (v3oo69y614hgiemyyld),
    .jp5nha2l14e7kx2jzpke      (jp5nha2l14e7kx2jzpke   ),
    .a4a48egkdkec8d9b_9     (a4a48egkdkec8d9b_9 ),
    .xwfmltfzahuj4qfn4qf2     (xwfmltfzahuj4qfn4qf2 ),
    .za9xg3zsqni_aeqmke      (za9xg3zsqni_aeqmke),
    .c1gmncmorg16sachdas      (c1gmncmorg16sachdas),
    .ggxoqcj7ytp1a4pjf7ee      (ggxoqcj7ytp1a4pjf7ee),
    .szrgf24or2mbt7w_yleh_vt(szrgf24or2mbt7w_yleh_vt),

    .p648zxn2luyxy8mt992a  (p648zxn2luyxy8mt992a ),
    .l3c127qdc9a2mfc13     (l3c127qdc9a2mfc13),
    .oq9b5zfhza9yvdoj      (oq9b5zfhza9yvdoj),
    .sg33s7pt45jp_          (sg33s7pt45jp_),
    .g9i9mf8jq7sc699j         (g9i9mf8jq7sc699j),

    .flcopog5zzpohfautwy     (flcopog5zzpohfautwy ),
    .gtb8f_h0g28itdr8k     (gtb8f_h0g28itdr8k ),
    .wf15djwi2hw25nz_       (wf15djwi2hw25nz_   ),
    .t1q5qmk9jzpf6glng4y   (t1q5qmk9jzpf6glng4y),
    .xsmx4zoewhbt07jxq     (xsmx4zoewhbt07jxq),


    .fkm9up63o1aeauaqhjb      (fkm9up63o1aeauaqhjb),
    .to_1lv9wnb3vmu6tvz5rc      (to_1lv9wnb3vmu6tvz5rc),
    .ju1kbeplcqy314lfj4       (ju1kbeplcqy314lfj4 ), 
    .r985fbe5k7hgzaq9i       (r985fbe5k7hgzaq9i ), 
    .bb04gpwotp2s6c7_p1gqkq      (bb04gpwotp2s6c7_p1gqkq), 
    .sqmey185cu3mtixhl      (sqmey185cu3mtixhl), 
    .rffcsd1o699ytclmx      (rffcsd1o699ytclmx),
    .roa7ljysjukna1_f_rh5l     (smuejl3ftpm3mb2zgxm3),
    .swz29iuutp9bjf_         (r29wk2o3a027n0g),
    .lbr88vbqtg8rht7320frde      (lbr88vbqtg8rht7320frde),
    .g7qq38mx3d58n1b15kcia      (g7qq38mx3d58n1b15kcia),
    .demg_fwfkmaeawq30t       (demg_fwfkmaeawq30t ),
    .grtb6ypa0px2gi1c       (grtb6ypa0px2gi1c ),
    .f128d8ws0seoihu1       (f128d8ws0seoihu1 ),
    .m2r7mfmq3afdd1ine      (m2r7mfmq3afdd1ine),
    .nhafiywg3hg_52kogwh      (nhafiywg3hg_52kogwh),
    .xrqayy6vigrw66z8a        (xrqayy6vigrw66z8a  ),
    .jyy72ywt9nbo10f2jxupacld    (jyy72ywt9nbo10f2jxupacld),
    .drz92qecqx_qtxwro      (drz92qecqx_qtxwro),

    .cxrbvs1hde7j8ziudd4ar      (cxrbvs1hde7j8ziudd4ar),
    .dmzxpdd5dgmp_2ip6h3_6      (dmzxpdd5dgmp_2ip6h3_6),
    .piv1ndd8n8dlaqx9       (piv1ndd8n8dlaqx9 ), 
    .r3rgwuaokuw68zin       (r3rgwuaokuw68zin ), 
    .m2aue5rcrjkbzdwbqvlzvr      (m2aue5rcrjkbzdwbqvlzvr), 
    .u7a8_cbg_zi4w4b4slc08      (u7a8_cbg_zi4w4b4slc08), 
    .fd_1f891ni339pnyzw63mg      (fd_1f891ni339pnyzw63mg),
    .zqnzorh6g9hnwsot5zr     (zqnzorh6g9hnwsot5zr),
    .wic6t212ob4tfa         (wic6t212ob4tfa),
    .p1g5jbgswdsx9v1j01103      (p1g5jbgswdsx9v1j01103),
    .zmrmpw_9vyme3rakn8br8e      (zmrmpw_9vyme3rakn8br8e),
    .sp2wnouu73ujsanhkn0       (sp2wnouu73ujsanhkn0 ),
    .n5w05rcecv47nvnfkkw5       (n5w05rcecv47nvnfkkw5 ),
    .dycy3iz66xw6yj5ea       (dycy3iz66xw6yj5ea ),
    .ro76scx3ggmfi4xp2bjx      (ro76scx3ggmfi4xp2bjx),
    .t9yh0n7ay27ft001vimu6      (t9yh0n7ay27ft001vimu6),
    .gpjxeoxkmf35ldn        (gpjxeoxkmf35ldn  ),
    .owde01ai01h2x5kn3_ng    (owde01ai01h2x5kn3_ng),
    .atur2zwqwk4mnbtz68l2      (atur2zwqwk4mnbtz68l2),



    .k5t515v6aa4oilq98cy6lrd8  (k5t515v6aa4oilq98cy6lrd8),
    .nbgnnsuqy2oogaz89vmbl1  (nbgnnsuqy2oogaz89vmbl1),
    .lkdpdaxvpxpy8w8hpchiph  (lkdpdaxvpxpy8w8hpchiph),
    .c1_3zcfvbhkc9cf7jgm7x   (c1_3zcfvbhkc9cf7jgm7x ),
    .cki2l53v3p6py9awsecgj  (cki2l53v3p6py9awsecgj),
    .ddjl2wsfh12b286nsrl3m5z  (ddjl2wsfh12b286nsrl3m5z),
    .y09wfhff_yx31yoe7cxv  (y09wfhff_yx31yoe7cxv),
    .zn80vi7_hafilb62kh72jx5d6 (zn80vi7_hafilb62kh72jx5d6),
    .e1wmvmyg_x8tobsfzpo     (e1wmvmyg_x8tobsfzpo),
    .sk43hkjk_z2mer7becad   (sk43hkjk_z2mer7becad ),
    .lo0fo8wk5o04f7ezwv474  (lo0fo8wk5o04f7ezwv474),
    .zutoko8hik1j9pa64jmpuw  (zutoko8hik1j9pa64jmpuw),
    .xqdmvgffpmzj6n0l23o   (xqdmvgffpmzj6n0l23o),
    .of_yab2i0nf9xv_tek5r   (of_yab2i0nf9xv_tek5r),
    .i1pzsd21aml3amhex3sf   (i1pzsd21aml3amhex3sf),

    .ltzq1n1rg2b9lrt8j0bs__wa  (ltzq1n1rg2b9lrt8j0bs__wa),
    .qui4zelf64bknwchxnz6  (qui4zelf64bknwchxnz6),
    .qf_hxpj8b9rdyabqx8q7l    (qf_hxpj8b9rdyabqx8q7l  ),
    .pqfnz7dk2f2khe5zxq0081lzv(pqfnz7dk2f2khe5zxq0081lzv  ),
    .j3gop6yag94s712e_mipwr484  (j3gop6yag94s712e_mipwr484),



    .hr7la0400ty0hiwk5d0     (ddl6fq6uyoan19ad7k1e7x6ut),
    .y1ipzdhzcfq282ups6ja     (tzjgmrua9xx8r7mtesjlse7ck),
    .lqv5bv6hq78ov_prb97v5z      (k3d3baof2jykxvcnolt ),
    .o15lm7no18top00l32ra     (sndcaz3jnaw0hhh4h34z),
    .ly1y__c5rzaa9xv_9_m1ppr     (e1ta255hq9y7b1vjvfw39tn9),
    .f1msmreidlchd7rf9w625     (ohegnxg1amg08qiwv7ye),
    .uarhtvlb5te5hc2g3      (bkvescuebx122g6u90z ),
    .g9ayxf51lhjl44vvw62u3     (ur2ihqhfmkb_slea1h731),
    .qfoijjxktg6dht3klxhyw5g     (r9qbbve4migk8rthusrhs),
    .gao2lzva86gawlwp2      (py08fct30wgf6i2wybxotxxp),
    .xpt7vgmhw7tamcpv2l      (yih871wxqwew7vzte1vz),
    .lrh4lctjvrz1rhm6b9oh      (ryikyr7mft0ec23vkfx4hc),
    .krh62hs2scfnb76m67a       (mtz1ahcj94t_b5n0lwt2np4),
    .pyfc_rgr3cwwvo34pf       (g4vv6e5kk3lia0_ykb0v),
    .u6xj18ku9lj1890n7       (orf3s90mdtxy8zht0g8),
    .s3lwpy5def9adgbbvx9ct       (blm6y03yzi8xj45jwfzaz_),
    .q96vjidg4x6ohxl7       (ddxbzfgl56dmh0jni2473),
   
    .b6m1vcd7bmemxnu99_zke     (yjy7mmnik6nbv0bv7fmw_),
    .vqld30a8qt13mzhwoc     (xlge7190nk7ecqh4flp7qwsxu),
    .jpa5gwkjwqz_j0a3cy1       (p7fyv9jmvb0qm4ay6qip  ),
    .kjxe2fpsacp9bx2_0fah36ij   (cyx_m80vjtb60akb9qxolqxs  ),
    .xsw8oz2ni13z6vac1tn61     (si3z5gtgqu6i6mr6lop_s0g1  ),

    .c0x_72w8ddbpt17fn      (c0x_72w8ddbpt17fn    ), 

    .tw0yf9aln_vu06k8l    (tw0yf9aln_vu06k8l  ), 
    .q84eo09gg53r2jj5a5xn    (q84eo09gg53r2jj5a5xn  ),
    .ss4cm882613f24kdjqsyl     (ss4cm882613f24kdjqsyl   ),
    .zm9uosdggg7ntkh97elw    (zm9uosdggg7ntkh97elw  ),
    .g_ahl2zik6mj75atnp_hej    (g_ahl2zik6mj75atnp_hej  ),
    .bjl40q8m35dwdn_mn9    (bjl40q8m35dwdn_mn9  ),
    .oefdpb9h9kx627r_0y5     (oefdpb9h9kx627r_0y5   ),
    .fh1jm1za5zvqmvdloi    (fh1jm1za5zvqmvdloi  ),
    .sp_0hv_ae5rrl9vagusi    (sp_0hv_ae5rrl9vagusi  ),
    .b4oh48a9a0g269ybrm     (b4oh48a9a0g269ybrm   ),
    .r5s3ykb7_xkl6t12oucf     (r5s3ykb7_xkl6t12oucf   ),
    .ssswxj_bpfx_ebsbj     (ssswxj_bpfx_ebsbj   ),
                           
    .fsj22rallxmhdrvuwenpq    (fsj22rallxmhdrvuwenpq  ),
    .yign8d_dhrow0i5wjts4bd    (yign8d_dhrow0i5wjts4bd  ),
    .hhlfu4md9k5v7naf1qt      (hhlfu4md9k5v7naf1qt    ),
    .j8m9s_du9fk99idlbh80  (j8m9s_du9fk99idlbh80), 
    .aapsfpke41r7dyya4ah    (aapsfpke41r7dyya4ah  ),

    .y1rlahaedj99shvl6uc      (y1rlahaedj99shvl6uc    ), 

    .rqf8b5xxbw0n1_qaw    (rqf8b5xxbw0n1_qaw  ), 
    .ocwcf75wgxfb1bawe    (ocwcf75wgxfb1bawe  ),
    .holgl43_yucp7f7l     (holgl43_yucp7f7l   ),
    .oyev1ipmdflkvxygwr    (oyev1ipmdflkvxygwr  ),
    .ihknw7_lm_572tv6s    (ihknw7_lm_572tv6s  ),
    .o31l03k34sdhwt4lkazfa5    (o31l03k34sdhwt4lkazfa5  ),
    .gy2sgn_1bpkac7msq3     (gy2sgn_1bpkac7msq3   ),
    .r_1u6q2lzkfus3o9nfl    (r_1u6q2lzkfus3o9nfl  ),
    .yff7wf8wth2vjkdjpr    (yff7wf8wth2vjkdjpr  ),
    .lppjhpov_5lgvx7n7fm4g     (lppjhpov_5lgvx7n7fm4g   ),
    .sdfg9zykj79rz_7thf9k     (sdfg9zykj79rz_7thf9k   ),
    .wt4e4tlh0u_4cljr2j5f9     (wt4e4tlh0u_4cljr2j5f9   ),
     
    .o4wuryrcvw13y2v5m6b6u    (o4wuryrcvw13y2v5m6b6u  ),
    .bt4howrm5xnf6u4fuwrum6    (bt4howrm5xnf6u4fuwrum6  ),
    .vnqegbzme0jutvf      (vnqegbzme0jutvf    ),
    .jdj122rbumyogtin6xpg97  (jdj122rbumyogtin6xpg97), 
    .p9mcc6npaw32uigcp6    (p9mcc6npaw32uigcp6  ),

    .gf33atgy                   (gf33atgy),
    .ru_wi                 (ru_wi)
  );

  ktpcxlh_26k125r eqvz5ukgpywwbk3v(
                           .rm1dxjejhq7dh3q5m (rm1dxjejhq7dh3q5m ),
                           .sxvvsxtbhyvt   (sxvvsxtbhyvt   ),

                           .pcr4upio7_tx37    (pcr4upio7_tx37    ), 
                           .uzklqlncpqqm1rav (uzklqlncpqqm1rav ),
                           .ortueunvnkx_l5m_j (ortueunvnkx_l5m_j ),
                           .hwuhtb7ucto_utk56 (hwuhtb7ucto_utk56 ),
                           .i1env2kmns7qvvuuc (i1env2kmns7qvvuuc ),
                           .g3s3vpafvy3i (g3s3vpafvy3i ),


                           .tia1md5dyh6kj4     (tia1md5dyh6kj4),
                           .c4ughu0qm5sfai (c4ughu0qm5sfai),
                           .indfp6mwqdqamez0mex (indfp6mwqdqamez0mex),

                           .p7ah58va5_2njbtv      (p7ah58va5_2njbtv), 
                           .u981qrwkgi5h0e72b__gg19w (u981qrwkgi5h0e72b__gg19w),  
                           .p0i2i3v3j1tclelx51     (p0i2i3v3j1tclelx51),
                       
                           .mum8f1rtatle7p_55y84     (mum8f1rtatle7p_55y84  ),   
                           .pn5bpwlp5ijfako9m5ao   (pn5bpwlp5ijfako9m5ao),
                           .g3s0qe2adsxsx8e6z     (g3s0qe2adsxsx8e6z  ),
                           .a1rl4lmhqp8ydyk07kqkn    (a1rl4lmhqp8ydyk07kqkn ),       
                           .apnns9jlj7y3y5bg8ynz   (apnns9jlj7y3y5bg8ynz),
                                                                      
                           .pmz7e4mgvbnmimqp0nghk     (pmz7e4mgvbnmimqp0nghk  ),
                           .j61algpxjoycxbswhgsuf   (j61algpxjoycxbswhgsuf),
                           .omq1ehm8hp4q9jgp5n5vn     (omq1ehm8hp4q9jgp5n5vn  ),
                           .fbv1q6sraswzp91zcn    (fbv1q6sraswzp91zcn ),       
                           .jv8kv41vzuir6an4iod   (jv8kv41vzuir6an4iod),
                                                                      
                                                                      
                           .qgl4363n31jx6xjyo05zkn     (qgl4363n31jx6xjyo05zkn  ),
                           .zec78nyllxlfwmpsgncluudf   (zec78nyllxlfwmpsgncluudf),
                           .dwvnjl0vxqkgd8t6dtvg5z    (dwvnjl0vxqkgd8t6dtvg5z ),
                           .gngmcj5c1jd85csel9ntru    (gngmcj5c1jd85csel9ntru ),       
                           .tkt93y5lfluzkia5plvksp   (tkt93y5lfluzkia5plvksp),
                                                                      
                           .km7co8hqm563od8ga_03_g     (km7co8hqm563od8ga_03_g  ),
                           .j4mas6g26o63wvnsdquh8c4p   (j4mas6g26o63wvnsdquh8c4p),
                           .nniah5mh0cunkhyln9    (nniah5mh0cunkhyln9 ),
                           .rcy_v3911lf33nza5j    (rcy_v3911lf33nza5j ),       
                           .g4nfgu53_rgc0632w8z97   (g4nfgu53_rgc0632w8z97),
                                                                      
                           .xzgkclcxsgfuseg87     (xzgkclcxsgfuseg87  ),
                           .djwlah5bo0r6myit6cal0t   (djwlah5bo0r6myit6cal0t),
                           .qu_ju3lv6nvkdbo8h11uf    (qu_ju3lv6nvkdbo8h11uf ),
                           .dydwz9i6k80alqfarffop    (dydwz9i6k80alqfarffop ),       
                           .ql1c7hzoj9kf__7r97krm   (ql1c7hzoj9kf__7r97krm),
                                                                      
                           .kp2j8kv1p1cjcg0lerwm     (kp2j8kv1p1cjcg0lerwm  ),
                           .v4a7g1wh3ivw0esp7dye0oiz   (v4a7g1wh3ivw0esp7dye0oiz),
                           .x9zuk21gpaj58uszvm5    (x9zuk21gpaj58uszvm5 ),
                           .n_h5oz0c5bo5rpevwjcu8    (n_h5oz0c5bo5rpevwjcu8 ),       
                           .ryid4_99ns1jc83at_88x   (ryid4_99ns1jc83at_88x),

                           .ysnexkrvlg2s55ajc5g69tm      (ysnexkrvlg2s55ajc5g69tm     ),           
                           .p7832rg37bbm7_ssxunhcj7     (p7832rg37bbm7_ssxunhcj7    ),          
                           .t1xtkdoie_8djygqlt1br56pwt    (t1xtkdoie_8djygqlt1br56pwt   ),         
                           .w33zvryieg8hhgy58581ny437h9 (w33zvryieg8hhgy58581ny437h9),           
                           .lv96t6re1w44borcb7do83ndua3vjy (lv96t6re1w44borcb7do83ndua3vjy),      


                           .dyl5g2vgrvy4mb3 (dyl5g2vgrvy4mb3),
                           .r5hpbriny8m67sv9e_ylgo1 (r5hpbriny8m67sv9e_ylgo1),


                           .q7ru87fmzxczveihcxcwh(y3iin4ygz2ed73_84l91h73),
                           .umc_2tn6um_9xaiy7_ksg0w(n8mvs5sw2pw48loob7jv6nmjdds),
                           .uiyh4da4134sjv7gnmc(dbzz2cu7abqy43de_ky433v),
                           .j8cjhcuf0m6xjvemdaz (gbb0bfnz8wqnjr5sufoh6ojt4pr),
                           .s_eowfyzlvx7gjv542upo (im70q80i1xh1y_5mo9ndr1),


                           .th06du2c8e2_b7k (k5t515v6aa4oilq98cy6lrd8),
                           .irjoi8wvo25u209f_5 (lkdpdaxvpxpy8w8hpchiph),

                           .zvk11dhgg2s67mkq (c1_3zcfvbhkc9cf7jgm7x), 
                           .fbzs0o4ysyuzeg_qdj (cki2l53v3p6py9awsecgj), 
                           .me1n4pvwxa7n3u8l05 (ddjl2wsfh12b286nsrl3m5z), 
                           .qaidts35dk5jcji0n (y09wfhff_yx31yoe7cxv), 
                           .uo0ftugxv_yuoh (zn80vi7_hafilb62kh72jx5d6), 
                           .dcj485cah5 (e1wmvmyg_x8tobsfzpo), 
                           .zxe59xihintdqfy9d (sk43hkjk_z2mer7becad), 
                           .u4r4b_6kp09q767q (lo0fo8wk5o04f7ezwv474),
                           .lhibcc3xwm6cy (zutoko8hik1j9pa64jmpuw),
                           .hc2ava5u3xa_bw0 (1'b0),
                           .erz5xg5fnrald (of_yab2i0nf9xv_tek5r),
                           .r19ik0uppwcr (i1pzsd21aml3amhex3sf),

                           .klkflmsyyf5w7ar (ltzq1n1rg2b9lrt8j0bs__wa),
                           .wy36iirxspfw56864 (qui4zelf64bknwchxnz6),
                           .lkjqs6kiuyj (qf_hxpj8b9rdyabqx8q7l),
                           .u245it8jnyhc3eqcy0 (pqfnz7dk2f2khe5zxq0081lzv),
                           .h7f6k_ims_9p3 (j3gop6yag94s712e_mipwr484), 

                           .cv0k9k_ijjnnylw1s7b_0d (cv0k9k_ijjnnylw1s7b_0d),
                           .swpk4h0gei3t_34xogbqncbo4 (swpk4h0gei3t_34xogbqncbo4),
                           .u9qmfl3rwx0dhr92z875vx7q (u9qmfl3rwx0dhr92z875vx7q),
                           .unu_x_i6jmr33nz0yitzk (unu_x_i6jmr33nz0yitzk), 
                           .bei3qhdtd0euq2emblogsu_x (bei3qhdtd0euq2emblogsu_x), 
                           .bf0_ynb648lqi7s93eieo0ln (bf0_ynb648lqi7s93eieo0ln),
                           .wf8o7p9_qfthhoxs747wyeuwkky (wf8o7p9_qfthhoxs747wyeuwkky),
                           .ygro7xue7x7rtdafkj3o4q4 (ygro7xue7x7rtdafkj3o4q4),
                           .drrly3q0ocg8d4pwh3m9o77 (drrly3q0ocg8d4pwh3m9o77),
                           .g654a6a9cesbee7xs6_uu9lu5 (g654a6a9cesbee7xs6_uu9lu5),
                           .x7fex0jf9da6a5v1c28upl72t (x7fex0jf9da6a5v1c28upl72t),
                           .ege0_1ufqm8i68zo4il6cwe46d (ege0_1ufqm8i68zo4il6cwe46d),
                           .ngyxf4n1cpcgks_s2zmgfb260 (ngyxf4n1cpcgks_s2zmgfb260), 
                           .c7m50uaw8lmp_iv4ci38q2 (c7m50uaw8lmp_iv4ci38q2), 
                           .m04a1mtbabwezldp1crh4rg6z (m04a1mtbabwezldp1crh4rg6z), 
                           .hwjq1ubtaei44lpk609fm2hb8 (hwjq1ubtaei44lpk609fm2hb8), 
                           .e28p_fu1k484ncul0p85ko (e28p_fu1k484ncul0p85ko), 

                           .a0_d_zdz9h9fgk46e8arf (a0_d_zdz9h9fgk46e8arf),
                           .twr9y24wxhs3qj2z9f2hzpaig6 (twr9y24wxhs3qj2z9f2hzpaig6),
                           .w8b46r9cof57xvd5zo1u4zh8 (w8b46r9cof57xvd5zo1u4zh8),
                           .wn1l4cmih7rwce1rb7wk3f9wy (wn1l4cmih7rwce1rb7wk3f9wy), 
                           .cgnzbuo_1yz6v42seb25duv (cgnzbuo_1yz6v42seb25duv), 
                           .zopev7f487spn9mwvuowqo (zopev7f487spn9mwvuowqo),
                           .p32jk0lb8g31kqlpvmllo75qim (p32jk0lb8g31kqlpvmllo75qim),
                           .g973rcaou05i456suvk_89dm (g973rcaou05i456suvk_89dm),
                           .wflv6rhfdwyxttak111v1l (wflv6rhfdwyxttak111v1l),
                           .ggsmt4nzx8pwlowehinqvk60f (ggsmt4nzx8pwlowehinqvk60f),
                           .xu8494ii8ectqb91224uuer (xu8494ii8ectqb91224uuer),
                           .r6rk128ijo839ougen9stbe (r6rk128ijo839ougen9stbe),
                           .xo6ciibewn8p8xey97jcsqi5 (xo6ciibewn8p8xey97jcsqi5), 
                           .evz1w_girwszyfnlcg4mwvtjo (evz1w_girwszyfnlcg4mwvtjo), 
                           .ju5f9fb1erjep_bv8gpfn6 (ju5f9fb1erjep_bv8gpfn6), 
                           .hadi1_f3quoaotjv5758x8kksot2 (hadi1_f3quoaotjv5758x8kksot2), 
                           .bdi4gjlb0po4ejcztowoqil7 (bdi4gjlb0po4ejcztowoqil7), 

                           .bvg_3t_ujbpur7b_h7f63jse (bvg_3t_ujbpur7b_h7f63jse),

                           .m5l6wu3uz_jfqasz8e3tsvrm (m5l6wu3uz_jfqasz8e3tsvrm),
                           .g9so28ythfl0q7xnk66p1   (g9so28ythfl0q7xnk66p1  ),
                           .e66wluxk71p2ldu3a1qk994bq (e66wluxk71p2ldu3a1qk994bq),
                           .ig2roj0y08x8_ntp3knz9rd (ig2roj0y08x8_ntp3knz9rd), 
                           .m7tq_t57mr5bovbb9ghffl4k (m7tq_t57mr5bovbb9ghffl4k),

                           .gpcgdcri3e6_fxrw8wwtysoqqr (gpcgdcri3e6_fxrw8wwtysoqqr),
                           .a6s4kxg1ibr6mntc85jik   (a6s4kxg1ibr6mntc85jik  ),
                           .hizzalmpwr8cqkxqi80wvbt65x (hizzalmpwr8cqkxqi80wvbt65x),

                           .gf33atgy (viuu21jzrv),
                           .ru_wi (ru_wi)
		  );

  assign rqy9v1_k_o74etonfc  = 1'b0;


  assign umnrzb6pv8dzc = (bhjn0b8ydp0vfsiy 
                      | dyl5g2vgrvy4mb3
                      | gbb0bfnz8wqnjr5sufoh6ojt4pr
                    )  



                  ;





  
  localparam es8lgh7odkstv = 7
                         +1 
                         ; 
  wire [es8lgh7odkstv-1:0] i9cfirek_4134tufh9mm;
  wire [es8lgh7odkstv-1:0] raqdtyu5e0petsz3set9f;
  assign raqdtyu5e0petsz3set9f = {
                               sndcaz3jnaw0hhh4h34z, 
                               e1ta255hq9y7b1vjvfw39tn9, 
                               ohegnxg1amg08qiwv7ye,
                               mtz1ahcj94t_b5n0lwt2np4,
                               g4vv6e5kk3lia0_ykb0v,
                               orf3s90mdtxy8zht0g8,
                               blm6y03yzi8xj45jwfzaz_,
                               ddxbzfgl56dmh0jni2473
                              };
  assign{
          o15lm7no18top00l32ra, 
          ly1y__c5rzaa9xv_9_m1ppr, 
          f1msmreidlchd7rf9w625,
          krh62hs2scfnb76m67a,
          pyfc_rgr3cwwvo34pf,
          u6xj18ku9lj1890n7,
          s3lwpy5def9adgbbvx9ct,
          q96vjidg4x6ohxl7
         } = i9cfirek_4134tufh9mm;

     ux607_gnrl_icb_w2n # (
       .LATE_READY (0),
       .AW (32),
       .USR_W (es8lgh7odkstv),
       .FIFO_OUTS_NUM (2),
       .FIFO_CUT_READY (1),
       .X_W (64),
       .Y_W (32)
     ) f5cdre_p3whzmfan7h(
       .i_icb_cmd_valid (ddl6fq6uyoan19ad7k1e7x6ut), 
       .i_icb_cmd_ready (tzjgmrua9xx8r7mtesjlse7ck), 
       .i_icb_cmd_read  (bkvescuebx122g6u90z), 
       .i_icb_cmd_addr  (k3d3baof2jykxvcnolt ), 
       .i_icb_cmd_wdata (ur2ihqhfmkb_slea1h731), 
       .i_icb_cmd_wmask (r9qbbve4migk8rthusrhs),
       .i_icb_cmd_lock  (py08fct30wgf6i2wybxotxxp ),
       .i_icb_cmd_excl  (yih871wxqwew7vzte1vz ),
       .i_icb_cmd_size  (ryikyr7mft0ec23vkfx4hc ),
       .i_icb_cmd_burst (3'b0),
       .i_icb_cmd_beat  (2'b0),
       .i_icb_cmd_usr   (raqdtyu5e0petsz3set9f),
   
       .i_icb_rsp_valid    (yjy7mmnik6nbv0bv7fmw_), 
       .i_icb_rsp_ready    (xlge7190nk7ecqh4flp7qwsxu), 
       .i_icb_rsp_err      (p7fyv9jmvb0qm4ay6qip ),
       .i_icb_rsp_excl_ok  (cyx_m80vjtb60akb9qxolqxs),
       .i_icb_rsp_rdata    (si3z5gtgqu6i6mr6lop_s0g1), 
       .i_icb_rsp_usr      (),
       
       .o_icb_cmd_valid  (hr7la0400ty0hiwk5d0),  
       .o_icb_cmd_ready  (y1ipzdhzcfq282ups6ja),  
       .o_icb_cmd_read   (uarhtvlb5te5hc2g3), 
       .o_icb_cmd_addr   (lqv5bv6hq78ov_prb97v5z), 
       .o_icb_cmd_wdata  (g9ayxf51lhjl44vvw62u3),  
       .o_icb_cmd_wmask  (qfoijjxktg6dht3klxhyw5g),
       .o_icb_cmd_lock   (gao2lzva86gawlwp2),
       .o_icb_cmd_excl   (xpt7vgmhw7tamcpv2l),
       .o_icb_cmd_size   (lrh4lctjvrz1rhm6b9oh),
       .o_icb_cmd_burst  (),
       .o_icb_cmd_beat   (),
       .o_icb_cmd_usr    (i9cfirek_4134tufh9mm),
   
       .o_icb_rsp_valid    (b6m1vcd7bmemxnu99_zke),
       .o_icb_rsp_ready    (vqld30a8qt13mzhwoc),
       .o_icb_rsp_err      (jpa5gwkjwqz_j0a3cy1 ),
       .o_icb_rsp_excl_ok  (kjxe2fpsacp9bx2_0fah36ij),
       .o_icb_rsp_rdata    (xsw8oz2ni13z6vac1tn61),
       .o_icb_rsp_usr      ({es8lgh7odkstv{1'b0}}),
   
       .clk (gf33atgy),  
       .rst_n (ru_wi)
    );




  wc2lipjaiimwuy7fx9zp32mr  gq_vyaa01iv9ga3b7blcdk5to5f8i(
     .e98zc_xde8d   (ju1kbeplcqy314lfj4),
     .lms849k     (r29wk2o3a027n0g),
     .dhzk00cwbk (smuejl3ftpm3mb2zgxm3)
  );


  assign buwj9_8l8bwj80kkinq9p = ~umnrzb6pv8dzc;

endmodule




























































module i6_4g5fspqlv1svn # (
  parameter onr7l = 32
) (
  input  [onr7l-1:0] qbjvs30wtb,
  output [onr7l-1:0] dqgck5s
);

  genvar i;
  generate 

  for(i=0;i<onr7l;i=i+1) begin: xiki82evp7g
    assign dqgck5s[i] = qbjvs30wtb[onr7l-1-i];
  end
  endgenerate


endmodule 



















module wc2lipjaiimwuy7fx9zp32mr (
  input  [32-1:0]   e98zc_xde8d,
  output lms849k,
  output dhzk00cwbk
  );







  wire [32-1:0] rqbq0wq0_ojyw61v5 = 32'h02000000;
  wire gay5seknj4v = (e98zc_xde8d[32-1:16] ==  rqbq0wq0_ojyw61v5[32-1:16]);

  wire [32-1:0] zys87dxafg7t5ll4o9 = 32'h0c000000;
  wire vbw11p9a6c6v = (e98zc_xde8d[32-1:16] ==  zys87dxafg7t5ll4o9[32-1:16]);

  wire [32-1:0] o4f5s69ex_fk0k7q13x = 32'h08000000;
  wire x68nff2f2n = (e98zc_xde8d[32-1:26] ==  o4f5s69ex_fk0k7q13x[32-1:26]);


  wire [32-1:0] dak283_f21dou11_grfkt = 32'h10000000;
  wire mpmtuxv2k_7aj0 = (e98zc_xde8d[32-1:20] ==  dak283_f21dou11_grfkt[32-1:20]);

  wire [32-1:0] r480zryu00zrqkrbk = 32'h00000000;
  wire g0tm56qj3_ = (e98zc_xde8d[32-1:12] ==  r480zryu00zrqkrbk[32-1:12]);

  wire lag657ufi590q = (1 > 0) & ((e98zc_xde8d & 32'hffff0000) ==  (32'h10010000 & 32'hffff0000));
  wire a_pyg8cnnivox4q = (1 > 1) & ((e98zc_xde8d & 32'b0) ==  (32'b0 & 32'b0));
  wire vjakd9g0uqfmj = (1 > 2) & ((e98zc_xde8d & 32'b0) ==  (32'b0 & 32'b0));
  wire rfva66olxq4g0jv = (1 > 3) & ((e98zc_xde8d & 32'b0) ==  (32'b0 & 32'b0));
  wire iywkhh6zq93vmewq = (1 > 4) & ((e98zc_xde8d & 32'b0) ==  (32'b0 & 32'b0));
  wire qcuu4wnp0nzvpfi = (1 > 5) & ((e98zc_xde8d & 32'b0) ==  (32'b0 & 32'b0));
  wire cbe5bswmcp52st9g = (1 > 6) & ((e98zc_xde8d & 32'b0) ==  (32'b0 & 32'b0));
  wire l8cs8556lz0hi_ = (1 > 7) & ((e98zc_xde8d & 32'b0) ==  (32'b0 & 32'b0));

  wire iyv1vya7vnywj5 = (1 > 0) & ((e98zc_xde8d & 32'hffffffff) ==  (32'h00000000 & 32'hffffffff));
  wire kiaw5590qrocm = (1 > 1) & ((e98zc_xde8d & 32'b0) ==  (32'b0 & 32'b0));
  wire z2ml5unafnd9 = (1 > 2) & ((e98zc_xde8d & 32'b0) ==  (32'b0 & 32'b0));
  wire pxvput9ybilro = (1 > 3) & ((e98zc_xde8d & 32'b0) ==  (32'b0 & 32'b0));
  wire lvspe8ctauaf = (1 > 4) & ((e98zc_xde8d & 32'b0) ==  (32'b0 & 32'b0));
  wire d7lmg6o1aplfg = (1 > 5) & ((e98zc_xde8d & 32'b0) ==  (32'b0 & 32'b0));
  wire wb0e5yne8mn = (1 > 6) & ((e98zc_xde8d & 32'b0) ==  (32'b0 & 32'b0));
  wire na3to0h77ey = (1 > 7) & ((e98zc_xde8d & 32'b0) ==  (32'b0 & 32'b0));



  assign dhzk00cwbk = ( 1'b0
                          | gay5seknj4v 
                          | vbw11p9a6c6v
                          | x68nff2f2n
                          | mpmtuxv2k_7aj0 
                          | lag657ufi590q
                          | a_pyg8cnnivox4q
                          | vjakd9g0uqfmj
                          | rfva66olxq4g0jv
                          | iywkhh6zq93vmewq
                          | qcuu4wnp0nzvpfi
                          | cbe5bswmcp52st9g
                          | l8cs8556lz0hi_
                          );
  assign lms849k	 = ( 1'b0
                          | iyv1vya7vnywj5
                          | kiaw5590qrocm
                          | z2ml5unafnd9
                          | pxvput9ybilro
                          | lvspe8ctauaf
                          | d7lmg6o1aplfg
                          | wb0e5yne8mn
                          | na3to0h77ey
                          | g0tm56qj3_
                          );

endmodule








































module k6pp01__lz7owqwu (
  input  dk2xhkj77a,
  input  zh6e0v0mmz,
  input  ru_wi,   



  input  avs1_7j,



  input  wxmxi1zq5,
  input  g0sg4nb6l3f,
  input  aey60u5dsgv,
  input  gf9zfb8tq9sv,
  input  iqg2bp31t,

  output uc5qxb4d2b28ye5,
  input  o2qkf90r783,

  input  z1l80uwh6vyyg34,

  output rn1o3sl83, 
  output zz5wo47gw146x4,
  output fgr486jx5kevbua,
  output pvfk1_6o89lmby,
  output xx87vzbpchg 
);

ux607_gnrl_dffr #(1) yebufj559oxyr(g0sg4nb6l3f, zz5wo47gw146x4, dk2xhkj77a, ru_wi);
ux607_gnrl_dffr #(1) iok8kkslh1d8_xzk0(aey60u5dsgv, fgr486jx5kevbua, dk2xhkj77a, ru_wi);
ux607_gnrl_dffr #(1) lwnytug2gf_nl5g9(gf9zfb8tq9sv, pvfk1_6o89lmby, dk2xhkj77a, ru_wi);
ux607_gnrl_dffr #(1) if7sx0g25tp7(iqg2bp31t, xx87vzbpchg, dk2xhkj77a, ru_wi);

wire ynmoengvzeeacdv;
wire j2doaov3294k;
ux607_gnrl_dffr #(1) b7csg1flnercwspofl7h7nd08_s0x(z1l80uwh6vyyg34, ynmoengvzeeacdv, zh6e0v0mmz, ru_wi);
ux607_gnrl_dffr #(1) l1gr8m0opa8_bcasz2vdbr4(o2qkf90r783, j2doaov3294k, zh6e0v0mmz, ru_wi);


wire zpfenxx7xnj;
wire zfte3vi0pfm7r3 = avs1_7j;
wire i8d70y0tuh1 = j2doaov3294k;
wire okwz17fsn22rg = zfte3vi0pfm7r3 | i8d70y0tuh1;
wire sznj6g2prhw57 = zfte3vi0pfm7r3 | (~i8d70y0tuh1);
ux607_gnrl_dfflr #(1) x9reesbi6nrw8 (okwz17fsn22rg, sznj6g2prhw57 , zpfenxx7xnj,  dk2xhkj77a, ru_wi);

assign uc5qxb4d2b28ye5 = zpfenxx7xnj;

wire egp2wyj39hah7;
ux607_gnrl_dffr #(1) aeijgq9e0xtivwsdbb(wxmxi1zq5, egp2wyj39hah7, dk2xhkj77a, ru_wi);

wire aobrltq_4foo4ih = wxmxi1zq5 & (~egp2wyj39hah7);
wire uctxe44ox7fjkgy = ynmoengvzeeacdv;
wire bdyay6mvy2t = aobrltq_4foo4ih | uctxe44ox7fjkgy; 
wire g3ukeq6cfbyz = aobrltq_4foo4ih | (~uctxe44ox7fjkgy); 
ux607_gnrl_dfflr #(1) en69d09blq0_emt9(bdyay6mvy2t, g3ukeq6cfbyz, rn1o3sl83, dk2xhkj77a, ru_wi);

endmodule




















module z_b0afg39m33f0qw0xb(
  input xoauecm4__2ehfjw,
  input by9h8n_pa6tbzsr5m,
  input [64-1:0] vf5xcr67bqhzlo43_,

  input [5-1:0] nra91e61s7u,
  input [64-1:0] yd6gywn1pn,
  input atqel3v0fzjjsz,
  output [64-1:0] wuke41p8s ,
  output [64-1:0] dez6c7e0g2w,
  output hk9dhg3ue,

  input  dk2xhkj77a,
  input  gf33atgy,
  input  ru_wi

  );


  wire ing9xff_u89x = yd6gywn1pn[nra91e61s7u[4:0]]; 

  wire [64-1:0] s6er21uf;
  wire l4ylal_gzpjxcqxv = ((s6er21uf == (~(64'b0))));
  wire t_fdz268gdu4    = xoauecm4__2ehfjw    |
                       ((~atqel3v0fzjjsz) & ing9xff_u89x);
  
  wire [64-1:0] qd_0tqy7a    = xoauecm4__2ehfjw  ? vf5xcr67bqhzlo43_ : (s6er21uf  + {{64-1{1'b0}},1'b1});
  
  ux607_gnrl_dfflr #(64) pyjjf7_txbyb (t_fdz268gdu4, qd_0tqy7a, s6er21uf   , dk2xhkj77a, ru_wi);
  assign wuke41p8s    = s6er21uf;
  
  

  assign hk9dhg3ue = 1'b1
                     & l4ylal_gzpjxcqxv 
                     & (~xoauecm4__2ehfjw) 
                     & ((~atqel3v0fzjjsz) & ing9xff_u89x);


  wire lr_3gt3i_ = by9h8n_pa6tbzsr5m;
  wire [64-1:0] md9mnc1f2lf;
  wire [64-1:0] xjj3qdbat = {{(64-9){1'b0}},vf5xcr67bqhzlo43_[8:4],4'b0};
  ux607_gnrl_dfflr #(64) q5hhls_dc9ewbi_ (lr_3gt3i_, xjj3qdbat, md9mnc1f2lf, gf33atgy, ru_wi);
  assign dez6c7e0g2w = md9mnc1f2lf;



endmodule




















module pcw8e2c5o1b_8(

  input aw82i964do,
  input y8_gkxsfle,

  input pydatzxqqi,
  input zmwq3e9oijvo7d7,
  input btwmhh91h50d5flgwx4o6pwu,

  input rb050tnl,
  input a94vd35etec4,
  input el7_p8jit09,
  input [12-1:0] e1go3iu,
  input izhvh9xxvwe2,
  input  [64-1:0] vf5xcr67bqhzlo43_,
  output [64-1:0] l9erxxpnphqd26vg9,

  output u2dvoyt5e7o_03z9z5,

  output um1_bmln_sf2i4vzbya_,

  output chjt9v0na3idosi9_0j5fe,
  output i72_qcuo70vljgkcb0fbj,

  output gjyhd0u2t3wy11drm07,
  output an0s8c6hcabd901wob_8zo,
  output e280ym1w614qoep160njy,

  input  ftp0juzjm2b587cyw5,
  input [31:0] fw4r5i27mgu0_,

  input [31:0] ij_sgq3rtvw2,
  input [31:0] k9jntnqwqp,


  output l0hrd_ubxbkay3zy8yz,

  input  gf33atgy,
  input  dk2xhkj77a,
  input  ru_wi

  );


  wire n8wchbzg_bh0842ixfy   ;
  wire w1cxh8pavpq2q547w7s   ;
  wire s7n9pzp2_lkcxidvvlx3 ;
  wire nr49mmvj0b7u6pwigbs_c ;
  wire ld5yq_b89a6sygy4db ;
  wire r4xqox_3f9vnymda3s ;

  wire kqlt5dn5j_9ssgd4c_6r   ;
  wire gjuz0xoojxqebmufd   ;
  wire g6pqxgmhk51jqwlulfg_8s ;
  wire gxdw47lxivtnooi_lskx ;
  wire btvvfzv564gvdraohzba0 ;
  wire w3e2huzmkc56w0h7beu0qb ;

  wire pt59ki6znxmbz3ghc6w   ;
  wire rtydd5c8x9iyr93kh   ;
  wire hptxny5nc0vmhpggj2c ;
  wire rsifu2upb5ml53lssvgzbe ;
  wire qhyfb11m9idvddngwcmhlg ;
  wire sbkvckx34gx323tsogkphx ;



  wire [31:0] zo6ft__dlnzl7dkr5qugp;
  wire [31:0] zwyd7w908csrxdqcda;
  wire [31:0] zh5di64w3lxurvyr3b    ;
  wire [31:0] skdz4fjkpq7ac0zq    ;
  wire [31:0] ow9fve_mr7bvw_wtmgl7   ;

  wire f3nolyi4jv6dte       = (e1go3iu == 12'hc00);
  wire e_kz098g        = (e1go3iu == 12'hc01);
  wire h0m0j6wupakd3zh     = (e1go3iu == 12'hc02);
  wire h8cnpp9r96r5jt3s  = (e1go3iu == 12'h306);
  wire yryyg8udb_4akvy  = (e1go3iu == 12'h106);
  wire tovyzk79in_cu3xt2fy = (e1go3iu == 12'h7ce);
  wire w4w2ra2eqzikjlg   = (e1go3iu == 12'hc03);
  wire ek78h0rdvr2jbnet5d   = (e1go3iu == 12'hc04);
  wire u62i7sw55i0ixtfn   = (e1go3iu == 12'hc05);
  wire b1u7q1bl0kcxqkk9lh   = (e1go3iu == 12'hc06);
  wire atqs6e48ujtlb69kq   = (e1go3iu == 12'hc07);
  wire m3s9phawcb5x9ggpi   = (e1go3iu == 12'hc08);
  wire bbupfe_9mnq91m2i5a2   = (e1go3iu == 12'hc09);
  wire msnj2ra1no6ygsuqoqp  = (e1go3iu == 12'hc0a);
  wire b9miqns7863wkebj4mx  = (e1go3iu == 12'hc0b);
  wire qwiayg271y7oeoc489  = (e1go3iu == 12'hc0c);
  wire x15dpsgnj3pv30wcv29s3  = (e1go3iu == 12'hc0d);
  wire cward2fs662rfpiht  = (e1go3iu == 12'hc0e);
  wire gqsc7i4m_9qz5uj9y3  = (e1go3iu == 12'hc0f);
  wire d3j6m80dne1gc9mm1  = (e1go3iu == 12'hc10);
  wire o7105xr36ce4gs38vq85  = (e1go3iu == 12'hc11);
  wire w8cnmp_jfu0jegjev  = (e1go3iu == 12'hc12);
  wire zd_u7f6fwo9yzoh1lvgpz  = (e1go3iu == 12'hc13);
  wire ppoyy50dz_tg4_hb2w1h  = (e1go3iu == 12'hc14);
  wire f4ojjkposvudt33guq  = (e1go3iu == 12'hc15);
  wire px4sutw16ys1h1dzhy90  = (e1go3iu == 12'hc16);
  wire uf6yc2ray6umf1z9y7ef  = (e1go3iu == 12'hc17);
  wire xpxi0rp39arefykelf4  = (e1go3iu == 12'hc18);
  wire ia3bm9atiopwvx52n7fux  = (e1go3iu == 12'hc19);
  wire kyby313yb5ca9djkzan  = (e1go3iu == 12'hc1a);
  wire firzx78r_e7t287kr  = (e1go3iu == 12'hc1b);
  wire nje80kd1i1pqhczz04  = (e1go3iu == 12'hc1c);
  wire om2footjljs7rqp3  = (e1go3iu == 12'hc1d);
  wire gwxoxa0q52lbsnv7  = (e1go3iu == 12'hc1e);
  wire iip0_by0868bv1qtl71qa  = (e1go3iu == 12'hc1f);

  
  wire exvzt_vf1mmht        = 1'b0;
  wire n0hf68fqn6tl         = 1'b0;
  wire di0_fvfp1wszdubcc      = 1'b0;
  wire ibihcuxenb1h85msj  = 1'b0;
  wire xiv4a67_96psl3rnqmp  = 1'b0;
  wire wrwhm830pc1woxrw  = 1'b0;
  wire cdtdn0g9ejv3kd5b  = 1'b0;
  wire ifxpvbmuyc_pwaz1l11  = 1'b0;
  wire da6ktvhw9k3es2c2d6ny  = 1'b0;
  wire szl7vw62u60k8_ec  = 1'b0;
  wire q6eajkfxmvgr7zezw = 1'b0;
  wire mt0yfe5jvmj3qq22q4gqv0 = 1'b0;
  wire k2iy3iepnrq2p0jbdy7 = 1'b0;
  wire vb68g5becvacfb5vw = 1'b0;
  wire cgsldj0fn4rv0jq9hgi3v = 1'b0;
  wire s7hwf0hvylsgsr_j6mxkj = 1'b0;
  wire ztgid5grbo8ocvbyx8ci = 1'b0;
  wire dxm9cwgp22i0alrice2k = 1'b0;
  wire cs6dm4hhsohstk8nrq = 1'b0;
  wire dkuckj4op4kdhw_5_t9j = 1'b0;
  wire zc_cweb5hhx8lixq4v = 1'b0;
  wire hkyq2ytin5akeb3ska = 1'b0;
  wire cfvznyjjj_o6wjz5u = 1'b0;
  wire iy71b9ln5s4dil291qeif = 1'b0;
  wire s1l4lgtbnqtz70zkucinz9 = 1'b0;
  wire vzlk0jh0n7gqlk3btw0 = 1'b0;
  wire e5uiim0onnmny13k15sm = 1'b0;
  wire snxumt7xwllnqlz3z = 1'b0;
  wire bxrvg7zifn8rg8_9pcb6 = 1'b0;
  wire vkf55sffofrevohin4uc = 1'b0;
  wire o55a67_plzpw6ma0_ = 1'b0;
  wire he4pomdstab68w18rn43_a = 1'b0;

  wire epn62p5usa2lzg6jq5l8l = (e1go3iu == 12'h7d1);
  wire xxhjtammdaysxdrgu_zq3 = (e1go3iu == 12'h7d3);
  
  wire etxyt17c       = el7_p8jit09 & f3nolyi4jv6dte   ;
  wire el4g39jr8hkit      = el7_p8jit09 & exvzt_vf1mmht  ;
  wire z2euvwgdf        = el7_p8jit09 & e_kz098g    ;
  wire ho_dmarc00       = el7_p8jit09 & n0hf68fqn6tl   ;
  wire vfr_4vmmkzbo6sp     = el7_p8jit09 & h0m0j6wupakd3zh ;
  wire s1qp0h9wv806    = el7_p8jit09 & di0_fvfp1wszdubcc;
  wire t6itxdn9xduvsw  = el7_p8jit09 & h8cnpp9r96r5jt3s;
  wire v9_rfvit5ecg18vn  = el7_p8jit09 & yryyg8udb_4akvy;
  wire xmfckyvtj9tkavm05cl = el7_p8jit09 & tovyzk79in_cu3xt2fy;
  wire saua96jt58f2vheh6d   = w4w2ra2eqzikjlg   & el7_p8jit09;
  wire vl3_0uq9ljyel49qm   = ek78h0rdvr2jbnet5d   & el7_p8jit09;
  wire e1ggq2ytz6l382l3jg   = u62i7sw55i0ixtfn   & el7_p8jit09;
  wire amzf3dktfg71xul98hi   = b1u7q1bl0kcxqkk9lh   & el7_p8jit09;
  wire lrpcc6xutnlegsrctfe   = atqs6e48ujtlb69kq   & el7_p8jit09; 
  wire b7zcd2bw3av_my   = m3s9phawcb5x9ggpi   & el7_p8jit09;
  wire xaw7ey1s6xx5rnkr   = bbupfe_9mnq91m2i5a2   & el7_p8jit09;
  wire o22k49cqoesn2oo2  = msnj2ra1no6ygsuqoqp  & el7_p8jit09;
  wire oska8h434cjp6zu6tiaq  = b9miqns7863wkebj4mx  & el7_p8jit09;
  wire ps7w4purbzr_i10x5i  = qwiayg271y7oeoc489  & el7_p8jit09;
  wire jjq1dceyzrzyes968  = x15dpsgnj3pv30wcv29s3  & el7_p8jit09;
  wire u8l2wf2m78gyp4j  = cward2fs662rfpiht  & el7_p8jit09;
  wire ux1k115isiuamx1e  = gqsc7i4m_9qz5uj9y3  & el7_p8jit09;
  wire up6ar789i17u5ra3fgor  = d3j6m80dne1gc9mm1  & el7_p8jit09;
  wire s8579tu61aj_f44  = o7105xr36ce4gs38vq85  & el7_p8jit09;
  wire hzabo0zo11yc4k37lqv  = w8cnmp_jfu0jegjev  & el7_p8jit09;
  wire ez47ti1d8gb0d93aro  = zd_u7f6fwo9yzoh1lvgpz  & el7_p8jit09;
  wire a3lqz8zf8izszn165yle  = ppoyy50dz_tg4_hb2w1h  & el7_p8jit09;
  wire e5s0u0c3jx64fvp0  = f4ojjkposvudt33guq  & el7_p8jit09;
  wire d3_m9cfog_c1tln5  = px4sutw16ys1h1dzhy90  & el7_p8jit09;
  wire wn9mt7zk595vn8p4mtxi  = uf6yc2ray6umf1z9y7ef  & el7_p8jit09;
  wire bobarmb1ci8jsesfgm  = xpxi0rp39arefykelf4  & el7_p8jit09;
  wire ue1jhuvuqi2ezv9vkr0  = ia3bm9atiopwvx52n7fux  & el7_p8jit09;
  wire ipcfszc_db2ggflm28l  = kyby313yb5ca9djkzan  & el7_p8jit09;
  wire rvc03sew724c0hn9  = firzx78r_e7t287kr  & el7_p8jit09;
  wire slbxk7eoe968is4m8  = nje80kd1i1pqhczz04  & el7_p8jit09;
  wire aqn143sj8jq7a8ved  = om2footjljs7rqp3  & el7_p8jit09;
  wire gbexxxkryjwqywc  = gwxoxa0q52lbsnv7  & el7_p8jit09;
  wire e0pc4vcinzwwn1jzcne  = iip0_by0868bv1qtl71qa  & el7_p8jit09;

  wire m938n32g7ii_hd0xc6  = ibihcuxenb1h85msj  & el7_p8jit09;
  wire fkut7_7ntf82jklyk  = xiv4a67_96psl3rnqmp  & el7_p8jit09;
  wire dy7yna1cgh95r_h  = wrwhm830pc1woxrw  & el7_p8jit09;
  wire cnpslhb184w6eseyj  = cdtdn0g9ejv3kd5b  & el7_p8jit09;
  wire anftxlsrefgv_3eqde5 = ifxpvbmuyc_pwaz1l11  & el7_p8jit09; 
  wire siyau38verruc640hm = da6ktvhw9k3es2c2d6ny  & el7_p8jit09;
  wire v7c7cqsl3pnqrtcl = szl7vw62u60k8_ec  & el7_p8jit09;
  wire k5p4vm2nwlnln4zhb= q6eajkfxmvgr7zezw & el7_p8jit09;
  wire knjj4hx9j_i8gnp_6s= mt0yfe5jvmj3qq22q4gqv0 & el7_p8jit09;
  wire cv_j2aqjiabk8f1jq= k2iy3iepnrq2p0jbdy7 & el7_p8jit09;
  wire ypy2mxdxutdtq4oq1e= vb68g5becvacfb5vw & el7_p8jit09;
  wire ulsb07fx57abjmdpn= cgsldj0fn4rv0jq9hgi3v & el7_p8jit09;
  wire sz4jk9vbnxc2616i= s7hwf0hvylsgsr_j6mxkj & el7_p8jit09;
  wire wn79nudil4f0lh9l4_t= ztgid5grbo8ocvbyx8ci & el7_p8jit09;
  wire vzl3dx5c5bzl5jxfx= dxm9cwgp22i0alrice2k & el7_p8jit09;
  wire hf_quo0pwq1ozp9d= cs6dm4hhsohstk8nrq & el7_p8jit09;
  wire fm56xxqzxuj614e6e4_ya= dkuckj4op4kdhw_5_t9j & el7_p8jit09;
  wire ldn075ya9eqsh88flm= zc_cweb5hhx8lixq4v & el7_p8jit09;
  wire ix8orbld9wpp9jpvaqq= hkyq2ytin5akeb3ska & el7_p8jit09;
  wire xrpb7eq89xqww5exjd3= cfvznyjjj_o6wjz5u & el7_p8jit09;
  wire gp36zq9cuerz4xycg= iy71b9ln5s4dil291qeif & el7_p8jit09;
  wire l079h3jnhz1d01_m60b= s1l4lgtbnqtz70zkucinz9 & el7_p8jit09;
  wire hkcs1nwvb3_53sa2nekga= vzlk0jh0n7gqlk3btw0 & el7_p8jit09;
  wire orkdamsky5y7oop2h549x= e5uiim0onnmny13k15sm & el7_p8jit09;
  wire ezbjbo9sr98uecjc= snxumt7xwllnqlz3z & el7_p8jit09;
  wire yhe9g6ovhg_zvw173= bxrvg7zifn8rg8_9pcb6 & el7_p8jit09;
  wire r9ioxzwla4_gvskfx61nj= vkf55sffofrevohin4uc & el7_p8jit09;
  wire jaw5sg6l42tk92f_u0ims= o55a67_plzpw6ma0_ & el7_p8jit09;
  wire vr_23ujl4y5nf7tmp= he4pomdstab68w18rn43_a & el7_p8jit09;

  wire x5oxp_rctueob44spc = epn62p5usa2lzg6jq5l8l & el7_p8jit09;
  wire ggkpi6kuym4_clvns8y41 = xxhjtammdaysxdrgu_zq3 & el7_p8jit09;

  wire zr77t9jqqfl       = f3nolyi4jv6dte       & izhvh9xxvwe2;
  wire ln2gmaay5u      = exvzt_vf1mmht      & izhvh9xxvwe2;
  wire nlw0hy8wyo7p9b4     = h0m0j6wupakd3zh     & izhvh9xxvwe2;
  wire aqlm13cyxzsa0    = di0_fvfp1wszdubcc    & izhvh9xxvwe2;
  wire ezm_pxkn5ocw0gh3a  = h8cnpp9r96r5jt3s  & izhvh9xxvwe2;
  wire duvtv2rabgkvc6sr  = yryyg8udb_4akvy  & izhvh9xxvwe2;
  wire a6zawvzasoonc9m = tovyzk79in_cu3xt2fy & izhvh9xxvwe2;
  wire u0ih2071ozg8hber   = w4w2ra2eqzikjlg   & izhvh9xxvwe2;
  wire pi8d3kvjvmzksr3l4   = ek78h0rdvr2jbnet5d   & izhvh9xxvwe2;
  wire mdeozybxpw0xhbo   = u62i7sw55i0ixtfn   & izhvh9xxvwe2;
  wire nbk22l2dcyhr_1oy   = b1u7q1bl0kcxqkk9lh   & izhvh9xxvwe2;
  wire o5jhzh7_ij66v0i0  = ibihcuxenb1h85msj  & izhvh9xxvwe2;
  wire okvdsshdlar77zxnf  = xiv4a67_96psl3rnqmp  & izhvh9xxvwe2;
  wire l4sxspwy35191q14ehw  = wrwhm830pc1woxrw  & izhvh9xxvwe2;
  wire esrovb5lx010_xdv52  = cdtdn0g9ejv3kd5b  & izhvh9xxvwe2;
  wire owkf2vvzq562oym6txue = epn62p5usa2lzg6jq5l8l & izhvh9xxvwe2;
  wire d42is86eedn26d0canw05y = xxhjtammdaysxdrgu_zq3 & izhvh9xxvwe2;



  wire rj6z05qy7n1gn3         = (e1go3iu == 12'hB00);
  wire z9dm6e6fby2aqjhy       = (e1go3iu == 12'hB02);
  wire f_es_90qk00g6opdh6x   = (e1go3iu == 12'hb03);
  wire fgzgnxejjal7h9rd   = (e1go3iu == 12'hb04);
  wire pcy6ei4r14x6ov28ryj   = (e1go3iu == 12'hb05);
  wire ocm0al346_oq8r_rk4saq   = (e1go3iu == 12'hb06);
  wire vsh2md0k8btsgo0fi   = (e1go3iu == 12'hb07);
  wire dy_4z613pc3tkdexyr2h7   = (e1go3iu == 12'hb08);
  wire xvlicu0ext8wdgxaxe   = (e1go3iu == 12'hb09);
  wire jsopbsj58ttr78ayz  = (e1go3iu == 12'hb0a);
  wire nk5xjy4ed8_rbp4pzyoxd  = (e1go3iu == 12'hb0b);
  wire e5g_pgu_jge9y177bzkk  = (e1go3iu == 12'hb0c);
  wire e2nua7o2jtyu0_g2gd  = (e1go3iu == 12'hb0d);
  wire it_k1w7q01tsk7pbr  = (e1go3iu == 12'hb0e);
  wire nzb9xw_eqn8iwu97rh1peh  = (e1go3iu == 12'hb0f);
  wire cw_4mgv8ahyjnni2ve  = (e1go3iu == 12'hb10);
  wire sdm457413c0japs5y1a5g  = (e1go3iu == 12'hb11);
  wire m4adp9ivz13luoy3p6n0  = (e1go3iu == 12'hb12);
  wire ako6g9a473i_du0c3c  = (e1go3iu == 12'hb13);
  wire i8k45cm1_hu1vr0yw  = (e1go3iu == 12'hb14);
  wire gnn1m6xd1mfmldxgvkpcm  = (e1go3iu == 12'hb15);
  wire pig91ircgpxokm21b0  = (e1go3iu == 12'hb16);
  wire zqi9hs4u7wi2xyenc  = (e1go3iu == 12'hb17);
  wire rjhbpotkkuqex6ngypg4  = (e1go3iu == 12'hb18);
  wire sujv8mssps3r3c0yvsk  = (e1go3iu == 12'hb19);
  wire x5z48ok_9ybuzzdqi  = (e1go3iu == 12'hb1a);
  wire dwcebcicgji91syba9vx35  = (e1go3iu == 12'hb1b);
  wire znodfh_5p8v6vy6i_29  = (e1go3iu == 12'hb1c);
  wire d0vcl63fuxsrv3a17eu  = (e1go3iu == 12'hb1d);
  wire bfix2k7kj4_cymu49h  = (e1go3iu == 12'hb1e);
  wire wh_whkedg1heijxqwe7ow  = (e1go3iu == 12'hb1f);



  wire iau25a3bde_t570        = 1'b0;
  wire ev00xx_m_ygc1f      = 1'b0;
  wire jywy59gh6tun9agkx  = 1'b0;
  wire c344aeyvo7fl8b4u5  = 1'b0;
  wire w54nli2z1nf5lhjabnv  = 1'b0;
  wire ql650jaoazwu2ppy27a  = 1'b0;
  wire bl3ql8yhyvm0j1hzey2  = 1'b0;
  wire szx_494r91n7lfktb50  = 1'b0;
  wire t8tz8_pdbmsiwmybl_6o  = 1'b0;
  wire ytbi6ubqw5j5__377nqb1 = 1'b0;
  wire tw_epfx1m93ilyi1be2m2 = 1'b0;
  wire n5fuwx4idtuxc7tct809c = 1'b0;
  wire fjx4uyep1wc4g3eu_vool = 1'b0;
  wire sjxk0a2xndebcgiml86 = 1'b0;
  wire g7iiqrs687lvtkb1ka = 1'b0;
  wire gzsdi4bs7ub5271rfqw = 1'b0;
  wire aeslm2tbru5a7_rixxj5m = 1'b0;
  wire p955_g_2i3jzj7cku4m = 1'b0;
  wire od0n9fap1dx46bxku_vuyuw = 1'b0;
  wire bpa8bumb36cks50x9nd = 1'b0;
  wire q_iz_w47hygrauver7g68 = 1'b0;
  wire tmj8i01xw0hzor8gu7 = 1'b0;
  wire pn_h7mrr0xdv0pe7dbs = 1'b0;
  wire mjbtpsfluunazpwqxsc5s7 = 1'b0;
  wire rmszohduwkl67ku12apqau = 1'b0;
  wire sx4gfxks7j_rndgzy65e = 1'b0;
  wire lqicd_93ufdrb29kpr15ee = 1'b0;
  wire gy7c8c0rxd6piv9j9e = 1'b0;
  wire uvornd3dvu5bss_cr_ = 1'b0;
  wire s_n6oz67gwnrvmq7tog5i_g = 1'b0;
  wire b2fdgj9jx0wm3vc1_z = 1'b0;


  wire b6gm4ouemqaev197d     = (e1go3iu == 12'h323);
  wire pay_6h44hjxz6wk     = (e1go3iu == 12'h324);
  wire qq2d9lmnwyq7st0_ek     = (e1go3iu == 12'h325);
  wire glodf0ee6jv3epkx     = (e1go3iu == 12'h326);
  wire e2mqz0x2e98z37fkk  = (e1go3iu == 12'h7cf);
  wire bcel2b05bj4rashyehe  = (e1go3iu == 12'h320);
  wire udpcqw7wqq89_qt    = (e1go3iu == 12'h7d4);

  wire a2152sbihdib         = rj6z05qy7n1gn3         & el7_p8jit09;
  wire j4haav4vmkkbvu        = iau25a3bde_t570        & el7_p8jit09;
  wire ayvfv16uem7g44db       = z9dm6e6fby2aqjhy       & el7_p8jit09;
  wire izi3g9mv6309mk      = ev00xx_m_ygc1f      & el7_p8jit09;
  wire ugg4ygya0e7093647   = f_es_90qk00g6opdh6x   & el7_p8jit09;
  wire f__p9_za313d8e0r   = fgzgnxejjal7h9rd   & el7_p8jit09;
  wire mhhil04nqg19efvv0_   = pcy6ei4r14x6ov28ryj   & el7_p8jit09;
  wire v9wd7zoiw_v9hv35ol   = ocm0al346_oq8r_rk4saq   & el7_p8jit09;
  wire lnt9d0tt4t2a3db   = vsh2md0k8btsgo0fi   & el7_p8jit09;
  wire fac3zsi4lyeiytxhn7kf   = dy_4z613pc3tkdexyr2h7   & el7_p8jit09;
  wire t__8hl9hyxi3xvs4ny9b   = xvlicu0ext8wdgxaxe   & el7_p8jit09;
  wire iqgwv1j2_ep8qmzp5  = jsopbsj58ttr78ayz  & el7_p8jit09;
  wire zxu8tncgm17k4ad6s6zht  = nk5xjy4ed8_rbp4pzyoxd  & el7_p8jit09;
  wire knzxmbncn5juz_ce  = e5g_pgu_jge9y177bzkk  & el7_p8jit09;
  wire tvij21_pu4txsd0y1cx  = e2nua7o2jtyu0_g2gd  & el7_p8jit09;
  wire qxuijdu07rcenvnwbyv  = it_k1w7q01tsk7pbr  & el7_p8jit09;
  wire wnbxn_fxj6b_act11jh  = nzb9xw_eqn8iwu97rh1peh  & el7_p8jit09;
  wire bxs3fd5gqwpta8nzaokh3  = cw_4mgv8ahyjnni2ve  & el7_p8jit09;
  wire u_psvzndlof4onsd  = sdm457413c0japs5y1a5g  & el7_p8jit09;
  wire x8jw220su9rl0jq_  = m4adp9ivz13luoy3p6n0  & el7_p8jit09;
  wire a9ck7mbx5squ3a1lvhz2k  = ako6g9a473i_du0c3c  & el7_p8jit09;
  wire ehvqob6usue9ira7hi0  = i8k45cm1_hu1vr0yw  & el7_p8jit09;
  wire k1pxlj3pkwavmz1ud  = gnn1m6xd1mfmldxgvkpcm  & el7_p8jit09;
  wire vyynogzp0y8paocqysgw6  = pig91ircgpxokm21b0  & el7_p8jit09;
  wire xhdifl547wtmxewr  = zqi9hs4u7wi2xyenc  & el7_p8jit09;
  wire lz0bdiv1w155ykfxore  = rjhbpotkkuqex6ngypg4  & el7_p8jit09;
  wire nkc01_m88jm8yvuk  = sujv8mssps3r3c0yvsk  & el7_p8jit09;
  wire ki3u2svcdfr7rqkq0t  = x5z48ok_9ybuzzdqi  & el7_p8jit09;
  wire ya_yx_os934avdybczhms  = dwcebcicgji91syba9vx35  & el7_p8jit09;
  wire z_oq7d2y6t47iv3mfg  = znodfh_5p8v6vy6i_29  & el7_p8jit09;
  wire g0eccm7oezzx707vxnpm  = d0vcl63fuxsrv3a17eu  & el7_p8jit09;
  wire zfid8vodcdo8565p7si  = bfix2k7kj4_cymu49h  & el7_p8jit09;
  wire oz7ge_4d2ujfqev27lrw  = wh_whkedg1heijxqwe7ow  & el7_p8jit09;

  wire cm95vygayrjauzd77y9_5  = jywy59gh6tun9agkx  & el7_p8jit09;
  wire mdd293u4cc_z55rhpw3r  = c344aeyvo7fl8b4u5  & el7_p8jit09;
  wire kdfqf15_615c_n1hqp240  = w54nli2z1nf5lhjabnv  & el7_p8jit09;
  wire n2tlae_r_pwl7wdmxlnj  = ql650jaoazwu2ppy27a  & el7_p8jit09;
  wire q5ytndij3ua9ib1m  = bl3ql8yhyvm0j1hzey2  & el7_p8jit09;
  wire xk45vrbmnrwmmfot  = szx_494r91n7lfktb50  & el7_p8jit09;
  wire cbv9gawz0e6r7q2l9knak  = t8tz8_pdbmsiwmybl_6o  & el7_p8jit09;
  wire zg1gmduc61biexqyjzo = ytbi6ubqw5j5__377nqb1 & el7_p8jit09;
  wire i4z3t0xqrj4n0k2r6yk_cx = tw_epfx1m93ilyi1be2m2 & el7_p8jit09;
  wire h6hkxd_ea12aa8c8sly = n5fuwx4idtuxc7tct809c & el7_p8jit09;
  wire b_1_5ck6n6yueyl_2v9z5u = fjx4uyep1wc4g3eu_vool & el7_p8jit09;
  wire bmp_xtvz_jvv62qvbj = sjxk0a2xndebcgiml86 & el7_p8jit09;
  wire ntd7kr9mt1ebjpvfu4c = g7iiqrs687lvtkb1ka & el7_p8jit09;
  wire z9muwxuqsv_ewu2r743d = gzsdi4bs7ub5271rfqw & el7_p8jit09;
  wire nle9soi2avivz7gudyq = aeslm2tbru5a7_rixxj5m & el7_p8jit09;
  wire acziqc95enp6s8nr3cc = p955_g_2i3jzj7cku4m & el7_p8jit09;
  wire mfm9kpan00kyxwlle48 = od0n9fap1dx46bxku_vuyuw & el7_p8jit09;
  wire l6tdd8ye847wqwafh = bpa8bumb36cks50x9nd & el7_p8jit09;
  wire vocnzx4d181giogclkir = q_iz_w47hygrauver7g68 & el7_p8jit09;
  wire x2x6qypmfdxybe0j_eg_cw = tmj8i01xw0hzor8gu7 & el7_p8jit09;
  wire cr_vfwpe75_b5prq2vv = pn_h7mrr0xdv0pe7dbs & el7_p8jit09;
  wire gld2hxb2y9qay27v7nh40w = mjbtpsfluunazpwqxsc5s7 & el7_p8jit09;
  wire xuogz8gc9n6zxgpcw = rmszohduwkl67ku12apqau & el7_p8jit09;
  wire qm00ottp0gobf61ju_a = sx4gfxks7j_rndgzy65e & el7_p8jit09;
  wire ubvjvn39xfkm6qq6o2cht = lqicd_93ufdrb29kpr15ee & el7_p8jit09;
  wire dgtul488nhno8epbk5 = gy7c8c0rxd6piv9j9e & el7_p8jit09;
  wire s44cgwshmsan_5igy = uvornd3dvu5bss_cr_ & el7_p8jit09;
  wire jy8uqowvshcdph_djto2 = s_n6oz67gwnrvmq7tog5i_g & el7_p8jit09;
  wire tt9wfj72e6ctzc9t08x = b2fdgj9jx0wm3vc1_z & el7_p8jit09;


  wire ql_5l6uckqbw5hfi     = b6gm4ouemqaev197d     & el7_p8jit09;
  wire ej22x93t1j2q09tv     = pay_6h44hjxz6wk     & el7_p8jit09;
  wire q19nl4ih99yhzfuh9y     = qq2d9lmnwyq7st0_ek     & el7_p8jit09;
  wire er98dls51_yfu8x     = glodf0ee6jv3epkx     & el7_p8jit09;
  wire z1goz2htj2xk6qeor  = e2mqz0x2e98z37fkk  & el7_p8jit09;
  wire wtv9m96nm63mgnzs  = bcel2b05bj4rashyehe  & el7_p8jit09;
  wire iaemsrwgo8mr8jg    = udpcqw7wqq89_qt    & el7_p8jit09;

  wire q42bebf3t5         = (rj6z05qy7n1gn3        | (f3nolyi4jv6dte        & n8wchbzg_bh0842ixfy  )) & izhvh9xxvwe2;
  wire f3kwcwki3be1        = (iau25a3bde_t570       | (exvzt_vf1mmht       & n8wchbzg_bh0842ixfy  )) & izhvh9xxvwe2;
  wire jbzubn1704nr       = (z9dm6e6fby2aqjhy      | (h0m0j6wupakd3zh      & w1cxh8pavpq2q547w7s  )) & izhvh9xxvwe2;
  wire s1oe4i7a9vc21i7aq      = (ev00xx_m_ygc1f     | (di0_fvfp1wszdubcc     & w1cxh8pavpq2q547w7s  )) & izhvh9xxvwe2;
  wire y8u5kzbhdn8_p5ow8   = (f_es_90qk00g6opdh6x  | (w4w2ra2eqzikjlg  & s7n9pzp2_lkcxidvvlx3)) & izhvh9xxvwe2;
  wire q1o7ht52byrd3lfjp4z   = (fgzgnxejjal7h9rd  | (ek78h0rdvr2jbnet5d  & nr49mmvj0b7u6pwigbs_c)) & izhvh9xxvwe2;
  wire uc0vudn7ey_lgwz4qvbd   = (pcy6ei4r14x6ov28ryj  | (u62i7sw55i0ixtfn  & ld5yq_b89a6sygy4db)) & izhvh9xxvwe2;
  wire mpq2ea0dzye6n2_   = (ocm0al346_oq8r_rk4saq  | (b1u7q1bl0kcxqkk9lh  & r4xqox_3f9vnymda3s)) & izhvh9xxvwe2;
  wire x5m4eoddc_s70vpwft3i  = (jywy59gh6tun9agkx | (ibihcuxenb1h85msj & s7n9pzp2_lkcxidvvlx3)) & izhvh9xxvwe2;
  wire q83ghpecvss6zodufz  = (c344aeyvo7fl8b4u5 | (xiv4a67_96psl3rnqmp & nr49mmvj0b7u6pwigbs_c)) & izhvh9xxvwe2;
  wire ia9e3_3rxhy9oryld  = (w54nli2z1nf5lhjabnv | (wrwhm830pc1woxrw & ld5yq_b89a6sygy4db)) & izhvh9xxvwe2;
  wire ib66r5rh9bioma8g2  = (ql650jaoazwu2ppy27a | (cdtdn0g9ejv3kd5b & r4xqox_3f9vnymda3s)) & izhvh9xxvwe2;

  wire d_05rkl4v555gcy     = b6gm4ouemqaev197d     & izhvh9xxvwe2;
  wire u4fpeyh2zr48j3     = pay_6h44hjxz6wk     & izhvh9xxvwe2;
  wire u_3xprdo9le2u     = qq2d9lmnwyq7st0_ek     & izhvh9xxvwe2;
  wire rd0tnkzv4tddj5ptx     = glodf0ee6jv3epkx     & izhvh9xxvwe2;
  wire zav0eknbhw3hwm0p33q  = e2mqz0x2e98z37fkk  & izhvh9xxvwe2;
  wire kutmbpkocduuslmby3m  = bcel2b05bj4rashyehe  & izhvh9xxvwe2;
  wire d3zb3re2q1lc9oe    = udpcqw7wqq89_qt    & izhvh9xxvwe2;


  wire s36z1abpqp = (~aw82i964do) & (~pydatzxqqi) & (~y8_gkxsfle);


  wire [64-1:0] bf27qv9x0e066       ;
  wire [64-1:0] h6t4j73gprqefaq03     ;
  wire [64-1:0] pswr19y981daoeip06 ;
  wire [64-1:0] ztnj98izh201_rom5xq8 ;
  wire [64-1:0] l4s95jgdzel2lkmw94oc ;
  wire [64-1:0] mx972bswiveneg0m3 ;
  wire [64-1:0] vmfc_5svhx5rgxdu ;
  wire [64-1:0] cuq97nfp4o3ljhlf ;
  wire [64-1:0] f_9h0p2ph4yezeyzc ;
  wire [64-1:0] fyzwg36odf2yct ;
  wire [31:0]           fu0bzqm3dpnn7r42aqz ;
  wire [31:0]           yide5ljyfkky_y2g6ek ;
  wire [31:0]           x1yjx1ygbxz3itn4unk;
  wire [31:0]           sv83e3r3rq0uml1xp2ye7lra;



  

  wire tfll_0gaqxiicaadd1zt  ;
  wire znk2n_ixp279qpzl9bd1h  ;
  wire t6z4oat4ia__jrbb1fwo;
  wire vf2yyykxidp14wtiif8t;
  wire y7knzb9echk4xuxrron9;
  wire si3w7ajsm0ju0o11tq5ly;

  wire o62cauzc87ljo = pydatzxqqi ? (zmwq3e9oijvo7d7 | btwmhh91h50d5flgwx4o6pwu): 1'b0;  

  wire clsdv9ql7   = o62cauzc87ljo | tfll_0gaqxiicaadd1zt   | ((~s36z1abpqp) & kqlt5dn5j_9ssgd4c_6r  ) | (s36z1abpqp & pt59ki6znxmbz3ghc6w  );  
  wire rr8nu2j9   = o62cauzc87ljo | znk2n_ixp279qpzl9bd1h   | ((~s36z1abpqp) & gjuz0xoojxqebmufd  ) | (s36z1abpqp & rtydd5c8x9iyr93kh  );
  wire x_mbnzybftw3x = o62cauzc87ljo | t6z4oat4ia__jrbb1fwo | ((~s36z1abpqp) & g6pqxgmhk51jqwlulfg_8s) | (s36z1abpqp & hptxny5nc0vmhpggj2c);
  wire rvfce__eg = o62cauzc87ljo | vf2yyykxidp14wtiif8t | ((~s36z1abpqp) & gxdw47lxivtnooi_lskx) | (s36z1abpqp & rsifu2upb5ml53lssvgzbe);
  wire t0t77x63g = o62cauzc87ljo | y7knzb9echk4xuxrron9 | ((~s36z1abpqp) & btvvfzv564gvdraohzba0) | (s36z1abpqp & qhyfb11m9idvddngwcmhlg);
  wire ddz3c_885r = o62cauzc87ljo | si3w7ajsm0ju0o11tq5ly | ((~s36z1abpqp) & w3e2huzmkc56w0h7beu0qb) | (s36z1abpqp & sbkvckx34gx323tsogkphx);
  
  wire gpbhuvuyoc812d;
  wire epcc1cvm2vllui4l;

  ihs34rgb4pudd03 n6b1yp267d4pby5srvff_1(
    .xoauecm4__2ehfjw   (q42bebf3t5), 


    .vf5xcr67bqhzlo43_   (vf5xcr67bqhzlo43_),
          
    .atqel3v0fzjjsz     (clsdv9ql7),
    .wuke41p8s      (bf27qv9x0e066),


    .hk9dhg3ue      (gpbhuvuyoc812d),
         
    .dk2xhkj77a        (dk2xhkj77a ),
    .ru_wi          (ru_wi) 
    );
  
  z_b0afg39m33f0qw0xb dtri55tmn9ffizi_469m(
    .xoauecm4__2ehfjw   (jbzubn1704nr),
    .by9h8n_pa6tbzsr5m   (1'b0),
    .vf5xcr67bqhzlo43_   (vf5xcr67bqhzlo43_),
          
    .nra91e61s7u        (5'b0),
    .yd6gywn1pn        ({{(64-1){1'b0}},ftp0juzjm2b587cyw5}),
    .atqel3v0fzjjsz     (rr8nu2j9),
    .wuke41p8s      (h6t4j73gprqefaq03),
    .dez6c7e0g2w      (),
  
    .hk9dhg3ue      (epcc1cvm2vllui4l),
         
    .dk2xhkj77a        (gf33atgy    ),
    .gf33atgy            (gf33atgy    ),
    .ru_wi          (ru_wi) 
    );
  
  wire [4:0] n3mubpr90bqtfvw5p533wvz9 = vmfc_5svhx5rgxdu[8:4];
  wire [4:0] awv46hulkygxrgy10h838iq_ = cuq97nfp4o3ljhlf[8:4];
  wire [4:0] qcghkdviru0w7xe2qoc5n84 = f_9h0p2ph4yezeyzc[8:4];
  wire [4:0] hmfouyhbmo7lz7yqpzfbhz = fyzwg36odf2yct[8:4];

  wire n5_szpwk_qwn65mqad;
  wire m0zd4aiaewfuvxrmvnw;
  wire m09xs6jue5l4cm6v0;
  wire u737k7dgs499utqiks;

      
   assign pswr19y981daoeip06   = 64'b0; 
   assign vmfc_5svhx5rgxdu     = 64'b0;  
   assign n5_szpwk_qwn65mqad   = 1'b0; 

   assign ztnj98izh201_rom5xq8   = 64'b0; 
   assign cuq97nfp4o3ljhlf     = 64'b0;  
   assign m0zd4aiaewfuvxrmvnw   = 1'b0; 

   assign l4s95jgdzel2lkmw94oc   = 64'b0; 
   assign f_9h0p2ph4yezeyzc     = 64'b0;  
   assign m09xs6jue5l4cm6v0   = 1'b0; 

   assign mx972bswiveneg0m3   = 64'b0; 
   assign fyzwg36odf2yct     = 64'b0;  
   assign u737k7dgs499utqiks   = 1'b0; 


  wire vtw_ipcez6h72qdp3fsmh = zav0eknbhw3hwm0p33q;
  wire [31:0] vus80e40sfur8oorvvfq;
  wire [31:0] zuek2ajp0_oih2cz0a = 32'b0;
  ux607_gnrl_dfflr #(32) s3tnb2k80ef9stf4cyyepq (vtw_ipcez6h72qdp3fsmh, zuek2ajp0_oih2cz0a, vus80e40sfur8oorvvfq, gf33atgy, ru_wi);
  assign fu0bzqm3dpnn7r42aqz = vus80e40sfur8oorvvfq;
  
  wire pewhcacpe3y_wbblo2x = kutmbpkocduuslmby3m;
  wire [31:0] kl25_6ll_hp6ez6d53l;
  wire [31:0] z626nm66qq0gyu7j7r = {29'b0,vf5xcr67bqhzlo43_[2],1'b0,vf5xcr67bqhzlo43_[0]};
  ux607_gnrl_dfflr #(32) or2bo8an2jxhfat6jbnyz9p (pewhcacpe3y_wbblo2x, z626nm66qq0gyu7j7r, kl25_6ll_hp6ez6d53l, gf33atgy, ru_wi);
  assign yide5ljyfkky_y2g6ek = kl25_6ll_hp6ez6d53l;
  
  assign tfll_0gaqxiicaadd1zt   = kl25_6ll_hp6ez6d53l[0];
  assign znk2n_ixp279qpzl9bd1h   = kl25_6ll_hp6ez6d53l[2];
  assign t6z4oat4ia__jrbb1fwo = kl25_6ll_hp6ez6d53l[3];
  assign vf2yyykxidp14wtiif8t = kl25_6ll_hp6ez6d53l[4];
  assign y7knzb9echk4xuxrron9 = kl25_6ll_hp6ez6d53l[5];
  assign si3w7ajsm0ju0o11tq5ly = kl25_6ll_hp6ez6d53l[6];
  
  wire zww3b0gwrn6iip24wf;
  wire p94xhwg2mjjdi16g_fd4h = u737k7dgs499utqiks;
  wire rceg531ybqbakabxtqud = d3zb3re2q1lc9oe & vf5xcr67bqhzlo43_[6];
  wire gm1n62_je4cf42hsns8pl7g = p94xhwg2mjjdi16g_fd4h | rceg531ybqbakabxtqud;
  wire tlp61m5adc8aualkwdmy9 = p94xhwg2mjjdi16g_fd4h & (~rceg531ybqbakabxtqud);
  ux607_gnrl_dfflr #(1) sssgnpzgau8sb9qn7z62f1flb0 (gm1n62_je4cf42hsns8pl7g, tlp61m5adc8aualkwdmy9, zww3b0gwrn6iip24wf, dk2xhkj77a, ru_wi);
  assign x1yjx1ygbxz3itn4unk[6] = zww3b0gwrn6iip24wf;
  assign sv83e3r3rq0uml1xp2ye7lra[6] = p94xhwg2mjjdi16g_fd4h;
  
  wire k6e0_yza67v2jxtpu04dj6;
  wire x2njxm7h7_nd6g2d_a00mvhzw = m09xs6jue5l4cm6v0;
  wire lp39nilru07s1jngqcio = d3zb3re2q1lc9oe & vf5xcr67bqhzlo43_[5];
  wire mzutqssu7gcaeozw3qql8 = x2njxm7h7_nd6g2d_a00mvhzw | lp39nilru07s1jngqcio;
  wire edd33o_1p3_lkuvewfqq81n3 = x2njxm7h7_nd6g2d_a00mvhzw & (~lp39nilru07s1jngqcio);
  ux607_gnrl_dfflr #(1) hl7szhqxucok67s4qoj4tmxyqo (mzutqssu7gcaeozw3qql8, edd33o_1p3_lkuvewfqq81n3, k6e0_yza67v2jxtpu04dj6, dk2xhkj77a, ru_wi);
  assign x1yjx1ygbxz3itn4unk[5] = k6e0_yza67v2jxtpu04dj6;
  assign sv83e3r3rq0uml1xp2ye7lra[5] = x2njxm7h7_nd6g2d_a00mvhzw;
  
  wire qz8n1j9eu82e13d8onz_;
  wire eqdh7ou2reaxdfus_jt7f5m = m0zd4aiaewfuvxrmvnw;
  wire a4pjlqbludrs7pan_gq8ty9 = d3zb3re2q1lc9oe & vf5xcr67bqhzlo43_[4];
  wire zs7ro8th45lctnezp5ilrl = eqdh7ou2reaxdfus_jt7f5m | a4pjlqbludrs7pan_gq8ty9;
  wire tnkipa54ueegg817530v = eqdh7ou2reaxdfus_jt7f5m & (~a4pjlqbludrs7pan_gq8ty9);
  ux607_gnrl_dfflr #(1) zwp_kff9z6exso317hgwa0a (zs7ro8th45lctnezp5ilrl, tnkipa54ueegg817530v, qz8n1j9eu82e13d8onz_, dk2xhkj77a, ru_wi);
  assign x1yjx1ygbxz3itn4unk[4] = qz8n1j9eu82e13d8onz_;
  assign sv83e3r3rq0uml1xp2ye7lra[4] = eqdh7ou2reaxdfus_jt7f5m;
  
  wire f3kwoj1931ziz5gnmtmxm94;
  wire sniy99ile4_f_silo26v0rmh = n5_szpwk_qwn65mqad;
  wire c7tap7nacs8uhyeisly2z4sx9 = d3zb3re2q1lc9oe & vf5xcr67bqhzlo43_[3];
  wire f27x6_ecvb5087annbgkog = sniy99ile4_f_silo26v0rmh | c7tap7nacs8uhyeisly2z4sx9;
  wire qnckz3g0jkfu84og1i1e = sniy99ile4_f_silo26v0rmh & (~c7tap7nacs8uhyeisly2z4sx9);
  ux607_gnrl_dfflr #(1) kemzr8h2umvylg1qr7oeuacrw (f27x6_ecvb5087annbgkog, qnckz3g0jkfu84og1i1e, f3kwoj1931ziz5gnmtmxm94, dk2xhkj77a, ru_wi);
  assign x1yjx1ygbxz3itn4unk[3] = f3kwoj1931ziz5gnmtmxm94;
  assign sv83e3r3rq0uml1xp2ye7lra[3] = sniy99ile4_f_silo26v0rmh;
  
  wire e5w3rdmlcmkrzp;
  wire nks4bgq3hjc4__xdrb = epcc1cvm2vllui4l;
  wire m6ktofruovkgbewctgevc = d3zb3re2q1lc9oe & vf5xcr67bqhzlo43_[2];
  wire po9mcm11udmp62v27 = nks4bgq3hjc4__xdrb | m6ktofruovkgbewctgevc;
  wire igh4ytj9iaitohpzng = 1'b0;
  ux607_gnrl_dfflr #(1) kz0_gxzmni98j76o7gurnbc (po9mcm11udmp62v27, igh4ytj9iaitohpzng, e5w3rdmlcmkrzp, gf33atgy, ru_wi);
  assign x1yjx1ygbxz3itn4unk[2] = e5w3rdmlcmkrzp;
  assign sv83e3r3rq0uml1xp2ye7lra[2] = nks4bgq3hjc4__xdrb;
  
  wire akb51beipsnqu;
  wire km0h_nhay_tegg86 = gpbhuvuyoc812d;
  wire eqw4ezqkmn6yp5gh = d3zb3re2q1lc9oe & vf5xcr67bqhzlo43_[0];
  wire pnzi9xh98300vqsxhv = km0h_nhay_tegg86 | eqw4ezqkmn6yp5gh;
  wire vn9r186wgz46sj3f28i = 1'b0;
  ux607_gnrl_dfflr #(1) fjn9y5k38wp94l2i5ndc (pnzi9xh98300vqsxhv, vn9r186wgz46sj3f28i, akb51beipsnqu, dk2xhkj77a, ru_wi);
  assign x1yjx1ygbxz3itn4unk[0] = akb51beipsnqu;
  assign sv83e3r3rq0uml1xp2ye7lra[0] = km0h_nhay_tegg86;
  
  assign x1yjx1ygbxz3itn4unk[31:7] = 25'b0;
  assign x1yjx1ygbxz3itn4unk[1] = 1'b0;
  
  assign sv83e3r3rq0uml1xp2ye7lra[31:7] = 25'b0;
  assign sv83e3r3rq0uml1xp2ye7lra[1] = 1'b0;
  
  
  wire [64-1:0] zylgiquxa5w        = bf27qv9x0e066;
  wire [64-1:0] ng7ft8ubwunj0lw      = h6t4j73gprqefaq03;
  wire [64-1:0] rc4v4mra6xuzgsxak5h  = pswr19y981daoeip06 ;
  wire [64-1:0] l8lnz796ln0mp8wb_ue  = ztnj98izh201_rom5xq8 ;
  wire [64-1:0] p2cbnkfxru9siuzmv6d  = l4s95jgdzel2lkmw94oc ;
  wire [64-1:0] abzpwx2is4xfioivt  = mx972bswiveneg0m3 ;
  wire [64-1:0] ftb953i514       = 64'b0; 
  wire [64-1:0] zcmenvygvs1tr7521     = 64'b0; 
  wire [64-1:0] b9v7h2vv4h5fgo4e = 64'b0; 
  wire [64-1:0] kd3g8vmacvpv2rvw1tf = 64'b0; 
  wire [64-1:0] c78inuigncqbtkf7sbp = 64'b0; 
  wire [64-1:0] jdkn85tb8sg_rwh8v3 = 64'b0; 
  
  wire [64-1:0] enhbns5z         = {k9jntnqwqp, ij_sgq3rtvw2};  
  wire [64-1:0] b1elz0eiw        = 64'b0;



  
  wire ofo2vvxrvlt9zy8 = ezm_pxkn5ocw0gh3a;
  wire [31:0] efc2znel8f5s_2d_;
  wire [31:0] iebtivwzxi3g_2ovi = {29'b0,vf5xcr67bqhzlo43_[2:0]};
  ux607_gnrl_dfflr #(32) uae39qbh9qtcrgtp (ofo2vvxrvlt9zy8, iebtivwzxi3g_2ovi, efc2znel8f5s_2d_, gf33atgy, ru_wi);
  assign zh5di64w3lxurvyr3b = efc2znel8f5s_2d_;
  
  wire d_foibnc5c0n5z4 = duvtv2rabgkvc6sr;
  wire [31:0] hqotlninf4u0xerhi;
  wire [31:0] fu0ahl2ekxxepw1v = {29'b0,vf5xcr67bqhzlo43_[2:0]};
  ux607_gnrl_dfflr #(32) llneyaw5qx3f43v3nfky (d_foibnc5c0n5z4, fu0ahl2ekxxepw1v, hqotlninf4u0xerhi, gf33atgy, ru_wi);
  assign skdz4fjkpq7ac0zq = hqotlninf4u0xerhi;
  
  wire n6k6_6werpw6mdojovc = a6zawvzasoonc9m;
  wire [31:0] p1e23t0ctg0ecxy8;
  wire [31:0] ah8c_kj5joxno4k = 32'b0;
  ux607_gnrl_dfflr #(32) s1qk37tntkg_0e1ayz (n6k6_6werpw6mdojovc, ah8c_kj5joxno4k, p1e23t0ctg0ecxy8, gf33atgy, ru_wi);
  assign ow9fve_mr7bvw_wtmgl7 = p1e23t0ctg0ecxy8;
 
  
  wire gt9ptrfsp8g3abmz7vgjp = owkf2vvzq562oym6txue;
  wire [31:0] nd4oyy8plwg2913kb4;
  wire [31:0] t19n7x98x494chy030h1 = 32'b0;
  ux607_gnrl_dfflr #(32) a9wv2vkrjq04iogc4u719r (gt9ptrfsp8g3abmz7vgjp, t19n7x98x494chy030h1, nd4oyy8plwg2913kb4, gf33atgy, ru_wi);
  assign zo6ft__dlnzl7dkr5qugp = nd4oyy8plwg2913kb4;
  
  wire g0r4hng9oumk8l4v541y = d42is86eedn26d0canw05y;
  wire [31:0] cpnh498hmivugspo;
  wire [31:0] vk1rwwjwqt4vxzjpjsr0ab = 32'b0;
  ux607_gnrl_dfflr #(32) l8k0_zo8le2u3j0t4j3k5a03 (g0r4hng9oumk8l4v541y, vk1rwwjwqt4vxzjpjsr0ab, cpnh498hmivugspo, gf33atgy, ru_wi);
  assign zwyd7w908csrxdqcda = cpnh498hmivugspo;

  
  
  

  assign n8wchbzg_bh0842ixfy   = ow9fve_mr7bvw_wtmgl7[0];
  assign w1cxh8pavpq2q547w7s   = ow9fve_mr7bvw_wtmgl7[2];
  assign s7n9pzp2_lkcxidvvlx3 = ow9fve_mr7bvw_wtmgl7[3];
  assign nr49mmvj0b7u6pwigbs_c = ow9fve_mr7bvw_wtmgl7[4];
  assign ld5yq_b89a6sygy4db = ow9fve_mr7bvw_wtmgl7[5];
  assign r4xqox_3f9vnymda3s = ow9fve_mr7bvw_wtmgl7[6];

  assign kqlt5dn5j_9ssgd4c_6r   = zo6ft__dlnzl7dkr5qugp[0];
  assign gjuz0xoojxqebmufd   = zo6ft__dlnzl7dkr5qugp[2];
  assign g6pqxgmhk51jqwlulfg_8s = zo6ft__dlnzl7dkr5qugp[3];
  assign gxdw47lxivtnooi_lskx = zo6ft__dlnzl7dkr5qugp[4];
  assign btvvfzv564gvdraohzba0 = zo6ft__dlnzl7dkr5qugp[5];
  assign w3e2huzmkc56w0h7beu0qb = zo6ft__dlnzl7dkr5qugp[6];

  assign pt59ki6znxmbz3ghc6w   = zwyd7w908csrxdqcda[0];
  assign rtydd5c8x9iyr93kh   = zwyd7w908csrxdqcda[2];
  assign hptxny5nc0vmhpggj2c = zwyd7w908csrxdqcda[3];
  assign rsifu2upb5ml53lssvgzbe = zwyd7w908csrxdqcda[4];
  assign qhyfb11m9idvddngwcmhlg = zwyd7w908csrxdqcda[5];
  assign sbkvckx34gx323tsogkphx = zwyd7w908csrxdqcda[6];


  assign l0hrd_ubxbkay3zy8yz = |(fu0bzqm3dpnn7r42aqz & sv83e3r3rq0uml1xp2ye7lra);

  wire rby_e01aj9mayt   = zh5di64w3lxurvyr3b[0];
  wire wy3w2aq98iuq6w   = zh5di64w3lxurvyr3b[1];
  wire x6zcn2iwg4w04   = zh5di64w3lxurvyr3b[2];
  wire edebxw2_52r74i4yub5n = zh5di64w3lxurvyr3b[3];
  wire n0a7cmohxqtifv1u_wo = zh5di64w3lxurvyr3b[4];
  wire jo9y8uxpmti4rhw6z = zh5di64w3lxurvyr3b[5];
  wire h_cfdp023jzvo4byhlbh = zh5di64w3lxurvyr3b[6];

  wire yvwjowlqpyzl2cdjmr   = skdz4fjkpq7ac0zq[0];
  wire eut3fa2784zt1m9g   = skdz4fjkpq7ac0zq[1];
  wire ra7birxz4b3gnigw   = skdz4fjkpq7ac0zq[2];
  wire mperzm5jjtfb4jk = skdz4fjkpq7ac0zq[3];
  wire gefz7vdqfjfmc7vx9p = skdz4fjkpq7ac0zq[4];
  wire gn663w5srr2mzrtvg = skdz4fjkpq7ac0zq[5];
  wire ed8kepqzl3lj7rms5l = skdz4fjkpq7ac0zq[6];






  assign {u2dvoyt5e7o_03z9z5, l9erxxpnphqd26vg9} = {1'b0,64'b0} 
                 | {rj6z05qy7n1gn3       , ({64{a2152sbihdib    }} & bf27qv9x0e066    )}
                 | {z9dm6e6fby2aqjhy     , ({64{ayvfv16uem7g44db  }} & h6t4j73gprqefaq03  )}
                 | {f_es_90qk00g6opdh6x , ({64{ugg4ygya0e7093647 }} & pswr19y981daoeip06 )}
                 | {fgzgnxejjal7h9rd , ({64{f__p9_za313d8e0r }} & ztnj98izh201_rom5xq8 )}
                 | {pcy6ei4r14x6ov28ryj , ({64{mhhil04nqg19efvv0_ }} & l4s95jgdzel2lkmw94oc )}
                 | {ocm0al346_oq8r_rk4saq , ({64{v9wd7zoiw_v9hv35ol }} & mx972bswiveneg0m3 )}
                 | {vsh2md0k8btsgo0fi   , ({64{lnt9d0tt4t2a3db  }} & {(64-1){1'b0}} )}
                 | {dy_4z613pc3tkdexyr2h7   , ({64{fac3zsi4lyeiytxhn7kf  }} & {(64-1){1'b0}} )}
                 | {xvlicu0ext8wdgxaxe   , ({64{t__8hl9hyxi3xvs4ny9b  }} & {(64-1){1'b0}} )}
                 | {jsopbsj58ttr78ayz  , ({64{iqgwv1j2_ep8qmzp5 }} & {(64-1){1'b0}} )}
                 | {nk5xjy4ed8_rbp4pzyoxd  , ({64{zxu8tncgm17k4ad6s6zht }} & {(64-1){1'b0}} )}
                 | {e5g_pgu_jge9y177bzkk  , ({64{knzxmbncn5juz_ce }} & {(64-1){1'b0}} )}
                 | {e2nua7o2jtyu0_g2gd  , ({64{tvij21_pu4txsd0y1cx }} & {(64-1){1'b0}} )}
                 | {it_k1w7q01tsk7pbr  , ({64{qxuijdu07rcenvnwbyv }} & {(64-1){1'b0}} )}
                 | {nzb9xw_eqn8iwu97rh1peh  , ({64{wnbxn_fxj6b_act11jh }} & {(64-1){1'b0}} )}
                 | {cw_4mgv8ahyjnni2ve  , ({64{bxs3fd5gqwpta8nzaokh3 }} & {(64-1){1'b0}} )}
                 | {sdm457413c0japs5y1a5g  , ({64{u_psvzndlof4onsd }} & {(64-1){1'b0}} )}
                 | {m4adp9ivz13luoy3p6n0  , ({64{x8jw220su9rl0jq_ }} & {(64-1){1'b0}} )}
                 | {ako6g9a473i_du0c3c  , ({64{a9ck7mbx5squ3a1lvhz2k }} & {(64-1){1'b0}} )}
                 | {i8k45cm1_hu1vr0yw  , ({64{ehvqob6usue9ira7hi0 }} & {(64-1){1'b0}} )}
                 | {gnn1m6xd1mfmldxgvkpcm  , ({64{k1pxlj3pkwavmz1ud }} & {(64-1){1'b0}} )}
                 | {pig91ircgpxokm21b0  , ({64{vyynogzp0y8paocqysgw6 }} & {(64-1){1'b0}} )}
                 | {zqi9hs4u7wi2xyenc  , ({64{xhdifl547wtmxewr }} & {(64-1){1'b0}} )}
                 | {rjhbpotkkuqex6ngypg4  , ({64{lz0bdiv1w155ykfxore }} & {(64-1){1'b0}} )}
                 | {sujv8mssps3r3c0yvsk  , ({64{nkc01_m88jm8yvuk }} & {(64-1){1'b0}} )}
                 | {x5z48ok_9ybuzzdqi  , ({64{ki3u2svcdfr7rqkq0t }} & {(64-1){1'b0}} )}
                 | {dwcebcicgji91syba9vx35  , ({64{ya_yx_os934avdybczhms }} & {(64-1){1'b0}} )}
                 | {znodfh_5p8v6vy6i_29  , ({64{z_oq7d2y6t47iv3mfg }} & {(64-1){1'b0}} )}
                 | {d0vcl63fuxsrv3a17eu  , ({64{g0eccm7oezzx707vxnpm }} & {(64-1){1'b0}} )}
                 | {bfix2k7kj4_cymu49h  , ({64{zfid8vodcdo8565p7si }} & {(64-1){1'b0}} )}
                 | {wh_whkedg1heijxqwe7ow  , ({64{oz7ge_4d2ujfqev27lrw }} & {(64-1){1'b0}} )}

                 | {bl3ql8yhyvm0j1hzey2  , ({64{q5ytndij3ua9ib1m }} & {(64-1){1'b0}} )}
                 | {szx_494r91n7lfktb50  , ({64{xk45vrbmnrwmmfot }} & {(64-1){1'b0}} )}
                 | {t8tz8_pdbmsiwmybl_6o  , ({64{cbv9gawz0e6r7q2l9knak }} & {(64-1){1'b0}} )}
                 | {ytbi6ubqw5j5__377nqb1 , ({64{zg1gmduc61biexqyjzo}} & {(64-1){1'b0}} )}
                 | {tw_epfx1m93ilyi1be2m2 , ({64{i4z3t0xqrj4n0k2r6yk_cx}} & {(64-1){1'b0}} )}
                 | {n5fuwx4idtuxc7tct809c , ({64{h6hkxd_ea12aa8c8sly}} & {(64-1){1'b0}} )}
                 | {fjx4uyep1wc4g3eu_vool , ({64{b_1_5ck6n6yueyl_2v9z5u}} & {(64-1){1'b0}} )}
                 | {sjxk0a2xndebcgiml86 , ({64{bmp_xtvz_jvv62qvbj}} & {(64-1){1'b0}} )}
                 | {g7iiqrs687lvtkb1ka , ({64{ntd7kr9mt1ebjpvfu4c}} & {(64-1){1'b0}} )}
                 | {gzsdi4bs7ub5271rfqw , ({64{z9muwxuqsv_ewu2r743d}} & {(64-1){1'b0}} )}
                 | {aeslm2tbru5a7_rixxj5m , ({64{nle9soi2avivz7gudyq}} & {(64-1){1'b0}} )}
                 | {p955_g_2i3jzj7cku4m , ({64{acziqc95enp6s8nr3cc}} & {(64-1){1'b0}} )}
                 | {od0n9fap1dx46bxku_vuyuw , ({64{mfm9kpan00kyxwlle48}} & {(64-1){1'b0}} )}
                 | {bpa8bumb36cks50x9nd , ({64{l6tdd8ye847wqwafh}} & {(64-1){1'b0}} )}
                 | {q_iz_w47hygrauver7g68 , ({64{vocnzx4d181giogclkir}} & {(64-1){1'b0}} )}
                 | {tmj8i01xw0hzor8gu7 , ({64{x2x6qypmfdxybe0j_eg_cw}} & {(64-1){1'b0}} )}
                 | {pn_h7mrr0xdv0pe7dbs , ({64{cr_vfwpe75_b5prq2vv}} & {(64-1){1'b0}} )}
                 | {mjbtpsfluunazpwqxsc5s7 , ({64{gld2hxb2y9qay27v7nh40w}} & {(64-1){1'b0}} )}
                 | {rmszohduwkl67ku12apqau , ({64{xuogz8gc9n6zxgpcw}} & {(64-1){1'b0}} )}
                 | {sx4gfxks7j_rndgzy65e , ({64{qm00ottp0gobf61ju_a}} & {(64-1){1'b0}} )}
                 | {lqicd_93ufdrb29kpr15ee , ({64{ubvjvn39xfkm6qq6o2cht}} & {(64-1){1'b0}} )}
                 | {gy7c8c0rxd6piv9j9e , ({64{dgtul488nhno8epbk5}} & {(64-1){1'b0}} )}
                 | {uvornd3dvu5bss_cr_ , ({64{s44cgwshmsan_5igy}} & {(64-1){1'b0}} )}
                 | {s_n6oz67gwnrvmq7tog5i_g , ({64{jy8uqowvshcdph_djto2}} & {(64-1){1'b0}} )}
                 | {b2fdgj9jx0wm3vc1_z , ({64{tt9wfj72e6ctzc9t08x}} & {(64-1){1'b0}} )}

                 | {bcel2b05bj4rashyehe, ({64{wtv9m96nm63mgnzs}} & {{(64-32){1'b0}}, yide5ljyfkky_y2g6ek}  )}
                 | {h8cnpp9r96r5jt3s , ({64{t6itxdn9xduvsw }} & {{(64-32){1'b0}}, zh5di64w3lxurvyr3b}  )}
                 | {yryyg8udb_4akvy , ({64{v9_rfvit5ecg18vn }} & {{(64-32){1'b0}}, skdz4fjkpq7ac0zq}  )}
                 | {f3nolyi4jv6dte      , ({64{etxyt17c      }} & zylgiquxa5w   )      }
                 | {exvzt_vf1mmht     , ({64{el4g39jr8hkit     }} & ftb953i514  )      }
                 | {e_kz098g       , ({64{z2euvwgdf       }} & enhbns5z    )      }
                 | {n0hf68fqn6tl      , ({64{ho_dmarc00      }} & b1elz0eiw   )      }
                 | {h0m0j6wupakd3zh    , ({64{vfr_4vmmkzbo6sp    }} & ng7ft8ubwunj0lw )      }
                 | {di0_fvfp1wszdubcc   , ({64{s1qp0h9wv806   }} & zcmenvygvs1tr7521)      }
                 | {w4w2ra2eqzikjlg , ({64{saua96jt58f2vheh6d }} & rc4v4mra6xuzgsxak5h )}
                 | {ek78h0rdvr2jbnet5d , ({64{vl3_0uq9ljyel49qm }} & l8lnz796ln0mp8wb_ue )}
                 | {u62i7sw55i0ixtfn , ({64{e1ggq2ytz6l382l3jg }} & p2cbnkfxru9siuzmv6d )}
                 | {b1u7q1bl0kcxqkk9lh , ({64{amzf3dktfg71xul98hi }} & abzpwx2is4xfioivt )}

                 | {ibihcuxenb1h85msj, ({64{m938n32g7ii_hd0xc6}} & b9v7h2vv4h5fgo4e)}
                 | {xiv4a67_96psl3rnqmp, ({64{fkut7_7ntf82jklyk}} & kd3g8vmacvpv2rvw1tf)}
                 | {wrwhm830pc1woxrw, ({64{dy7yna1cgh95r_h}} & c78inuigncqbtkf7sbp)}
                 | {cdtdn0g9ejv3kd5b, ({64{cnpslhb184w6eseyj}} & jdkn85tb8sg_rwh8v3)}

                 | {atqs6e48ujtlb69kq   , ({64{lrpcc6xutnlegsrctfe  }} & {(64-1){1'b0}} )}
                 | {m3s9phawcb5x9ggpi   , ({64{b7zcd2bw3av_my  }} & {(64-1){1'b0}} )}
                 | {bbupfe_9mnq91m2i5a2   , ({64{xaw7ey1s6xx5rnkr  }} & {(64-1){1'b0}} )}
                 | {msnj2ra1no6ygsuqoqp  , ({64{o22k49cqoesn2oo2 }} & {(64-1){1'b0}} )}
                 | {b9miqns7863wkebj4mx  , ({64{oska8h434cjp6zu6tiaq }} & {(64-1){1'b0}} )}
                 | {qwiayg271y7oeoc489  , ({64{ps7w4purbzr_i10x5i }} & {(64-1){1'b0}} )}
                 | {x15dpsgnj3pv30wcv29s3  , ({64{jjq1dceyzrzyes968 }} & {(64-1){1'b0}} )}
                 | {cward2fs662rfpiht  , ({64{u8l2wf2m78gyp4j }} & {(64-1){1'b0}} )}
                 | {gqsc7i4m_9qz5uj9y3  , ({64{ux1k115isiuamx1e }} & {(64-1){1'b0}} )}
                 | {d3j6m80dne1gc9mm1  , ({64{up6ar789i17u5ra3fgor }} & {(64-1){1'b0}} )}
                 | {o7105xr36ce4gs38vq85  , ({64{s8579tu61aj_f44 }} & {(64-1){1'b0}} )}
                 | {w8cnmp_jfu0jegjev  , ({64{hzabo0zo11yc4k37lqv }} & {(64-1){1'b0}} )}
                 | {zd_u7f6fwo9yzoh1lvgpz  , ({64{ez47ti1d8gb0d93aro }} & {(64-1){1'b0}} )}
                 | {ppoyy50dz_tg4_hb2w1h  , ({64{a3lqz8zf8izszn165yle }} & {(64-1){1'b0}} )}
                 | {f4ojjkposvudt33guq  , ({64{e5s0u0c3jx64fvp0 }} & {(64-1){1'b0}} )}
                 | {px4sutw16ys1h1dzhy90  , ({64{d3_m9cfog_c1tln5 }} & {(64-1){1'b0}} )}
                 | {uf6yc2ray6umf1z9y7ef  , ({64{wn9mt7zk595vn8p4mtxi }} & {(64-1){1'b0}} )}
                 | {xpxi0rp39arefykelf4  , ({64{bobarmb1ci8jsesfgm }} & {(64-1){1'b0}} )}
                 | {ia3bm9atiopwvx52n7fux  , ({64{ue1jhuvuqi2ezv9vkr0 }} & {(64-1){1'b0}} )}
                 | {kyby313yb5ca9djkzan  , ({64{ipcfszc_db2ggflm28l }} & {(64-1){1'b0}} )}
                 | {firzx78r_e7t287kr  , ({64{rvc03sew724c0hn9 }} & {(64-1){1'b0}} )}
                 | {nje80kd1i1pqhczz04  , ({64{slbxk7eoe968is4m8 }} & {(64-1){1'b0}} )}
                 | {om2footjljs7rqp3  , ({64{aqn143sj8jq7a8ved }} & {(64-1){1'b0}} )}
                 | {gwxoxa0q52lbsnv7  , ({64{gbexxxkryjwqywc }} & {(64-1){1'b0}} )}
                 | {iip0_by0868bv1qtl71qa  , ({64{e0pc4vcinzwwn1jzcne }} & {(64-1){1'b0}} )}

                 | {ifxpvbmuyc_pwaz1l11  , ({64{anftxlsrefgv_3eqde5 }} & {(64-1){1'b0}} )}
                 | {da6ktvhw9k3es2c2d6ny  , ({64{siyau38verruc640hm }} & {(64-1){1'b0}} )}
                 | {szl7vw62u60k8_ec  , ({64{v7c7cqsl3pnqrtcl }} & {(64-1){1'b0}} )}
                 | {q6eajkfxmvgr7zezw , ({64{k5p4vm2nwlnln4zhb}} & {(64-1){1'b0}} )}
                 | {mt0yfe5jvmj3qq22q4gqv0 , ({64{knjj4hx9j_i8gnp_6s}} & {(64-1){1'b0}} )}
                 | {k2iy3iepnrq2p0jbdy7 , ({64{cv_j2aqjiabk8f1jq}} & {(64-1){1'b0}} )}
                 | {vb68g5becvacfb5vw , ({64{ypy2mxdxutdtq4oq1e}} & {(64-1){1'b0}} )}
                 | {cgsldj0fn4rv0jq9hgi3v , ({64{ulsb07fx57abjmdpn}} & {(64-1){1'b0}} )}
                 | {s7hwf0hvylsgsr_j6mxkj , ({64{sz4jk9vbnxc2616i}} & {(64-1){1'b0}} )}
                 | {ztgid5grbo8ocvbyx8ci , ({64{wn79nudil4f0lh9l4_t}} & {(64-1){1'b0}} )}
                 | {dxm9cwgp22i0alrice2k , ({64{vzl3dx5c5bzl5jxfx}} & {(64-1){1'b0}} )}
                 | {cs6dm4hhsohstk8nrq , ({64{hf_quo0pwq1ozp9d}} & {(64-1){1'b0}} )}
                 | {dkuckj4op4kdhw_5_t9j , ({64{fm56xxqzxuj614e6e4_ya}} & {(64-1){1'b0}} )}
                 | {zc_cweb5hhx8lixq4v , ({64{ldn075ya9eqsh88flm}} & {(64-1){1'b0}} )}
                 | {hkyq2ytin5akeb3ska , ({64{ix8orbld9wpp9jpvaqq}} & {(64-1){1'b0}} )}
                 | {cfvznyjjj_o6wjz5u , ({64{xrpb7eq89xqww5exjd3}} & {(64-1){1'b0}} )}
                 | {iy71b9ln5s4dil291qeif , ({64{gp36zq9cuerz4xycg}} & {(64-1){1'b0}} )}
                 | {s1l4lgtbnqtz70zkucinz9 , ({64{l079h3jnhz1d01_m60b}} & {(64-1){1'b0}} )}
                 | {vzlk0jh0n7gqlk3btw0 , ({64{hkcs1nwvb3_53sa2nekga}} & {(64-1){1'b0}} )}
                 | {e5uiim0onnmny13k15sm , ({64{orkdamsky5y7oop2h549x}} & {(64-1){1'b0}} )}
                 | {snxumt7xwllnqlz3z , ({64{ezbjbo9sr98uecjc}} & {(64-1){1'b0}} )}
                 | {bxrvg7zifn8rg8_9pcb6 , ({64{yhe9g6ovhg_zvw173}} & {(64-1){1'b0}} )}
                 | {vkf55sffofrevohin4uc , ({64{r9ioxzwla4_gvskfx61nj}} & {(64-1){1'b0}} )}
                 | {o55a67_plzpw6ma0_ , ({64{jaw5sg6l42tk92f_u0ims}} & {(64-1){1'b0}} )}
                 | {he4pomdstab68w18rn43_a , ({64{vr_23ujl4y5nf7tmp}} & {(64-1){1'b0}} )}

              ;



    wire s32nr2e9a6f4hrqy4n775or =
                   atqs6e48ujtlb69kq  
                 | m3s9phawcb5x9ggpi  
                 | bbupfe_9mnq91m2i5a2  
                 | msnj2ra1no6ygsuqoqp 
                 | b9miqns7863wkebj4mx 
                 | qwiayg271y7oeoc489 
                 | x15dpsgnj3pv30wcv29s3 
                 | cward2fs662rfpiht 
                 | gqsc7i4m_9qz5uj9y3 
                 | d3j6m80dne1gc9mm1 
                 | o7105xr36ce4gs38vq85 
                 | w8cnmp_jfu0jegjev 
                 | zd_u7f6fwo9yzoh1lvgpz 
                 | ppoyy50dz_tg4_hb2w1h 
                 | f4ojjkposvudt33guq 
                 | px4sutw16ys1h1dzhy90 
                 | uf6yc2ray6umf1z9y7ef 
                 | xpxi0rp39arefykelf4 
                 | ia3bm9atiopwvx52n7fux 
                 | kyby313yb5ca9djkzan 
                 | firzx78r_e7t287kr 
                 | nje80kd1i1pqhczz04 
                 | om2footjljs7rqp3 
                 | gwxoxa0q52lbsnv7 
                 | iip0_by0868bv1qtl71qa 

                 | ifxpvbmuyc_pwaz1l11 
                 | da6ktvhw9k3es2c2d6ny 
                 | szl7vw62u60k8_ec 
                 | q6eajkfxmvgr7zezw
                 | mt0yfe5jvmj3qq22q4gqv0
                 | k2iy3iepnrq2p0jbdy7
                 | vb68g5becvacfb5vw
                 | cgsldj0fn4rv0jq9hgi3v
                 | s7hwf0hvylsgsr_j6mxkj
                 | ztgid5grbo8ocvbyx8ci
                 | dxm9cwgp22i0alrice2k
                 | cs6dm4hhsohstk8nrq
                 | dkuckj4op4kdhw_5_t9j
                 | zc_cweb5hhx8lixq4v
                 | hkyq2ytin5akeb3ska
                 | cfvznyjjj_o6wjz5u
                 | iy71b9ln5s4dil291qeif
                 | s1l4lgtbnqtz70zkucinz9
                 | vzlk0jh0n7gqlk3btw0
                 | e5uiim0onnmny13k15sm
                 | snxumt7xwllnqlz3z
                 | bxrvg7zifn8rg8_9pcb6
                 | vkf55sffofrevohin4uc
                 | o55a67_plzpw6ma0_
                 | he4pomdstab68w18rn43_a;

  assign um1_bmln_sf2i4vzbya_ = ( 
                    f3nolyi4jv6dte
                  | exvzt_vf1mmht    
                  | e_kz098g
                  | n0hf68fqn6tl
                  | h0m0j6wupakd3zh   
                  | di0_fvfp1wszdubcc  
                  | w4w2ra2eqzikjlg 
                  | ek78h0rdvr2jbnet5d 
                  | u62i7sw55i0ixtfn 
                  | b1u7q1bl0kcxqkk9lh 

                  | ibihcuxenb1h85msj
                  | xiv4a67_96psl3rnqmp
                  | wrwhm830pc1woxrw
                  | cdtdn0g9ejv3kd5b

                  | s32nr2e9a6f4hrqy4n775or 
                 )
               ;


  
  assign i72_qcuo70vljgkcb0fbj = 
      
                     a94vd35etec4 &  
                   
               ( 
                    f3nolyi4jv6dte        
                  | exvzt_vf1mmht       
                  | e_kz098g      
                  | n0hf68fqn6tl    
                  | h0m0j6wupakd3zh      
                  | di0_fvfp1wszdubcc     
                  | w4w2ra2eqzikjlg  
                  | ibihcuxenb1h85msj 
                  | ek78h0rdvr2jbnet5d  
                  | xiv4a67_96psl3rnqmp 
                  | u62i7sw55i0ixtfn  
                  | wrwhm830pc1woxrw 
                  | b1u7q1bl0kcxqkk9lh  
                  | cdtdn0g9ejv3kd5b 

                  | s32nr2e9a6f4hrqy4n775or 
                 )
               ;


  assign chjt9v0na3idosi9_0j5fe = s36z1abpqp & el7_p8jit09 &  
                   
                   
               ( 
                    (((~rby_e01aj9mayt  ) | (~yvwjowlqpyzl2cdjmr  )) & f3nolyi4jv6dte        )
                  | (((~rby_e01aj9mayt  ) | (~yvwjowlqpyzl2cdjmr  )) & exvzt_vf1mmht       )
                  | (((~wy3w2aq98iuq6w  ) | (~eut3fa2784zt1m9g  )) & e_kz098g         )
                  | (((~wy3w2aq98iuq6w  ) | (~eut3fa2784zt1m9g  )) & n0hf68fqn6tl        )
                  | (((~x6zcn2iwg4w04  ) | (~ra7birxz4b3gnigw  )) & h0m0j6wupakd3zh      )
                  | (((~x6zcn2iwg4w04  ) | (~ra7birxz4b3gnigw  )) & di0_fvfp1wszdubcc     )
                  | (((~edebxw2_52r74i4yub5n) | (~mperzm5jjtfb4jk)) & w4w2ra2eqzikjlg  )
                  | (((~edebxw2_52r74i4yub5n) | (~mperzm5jjtfb4jk)) & ibihcuxenb1h85msj )
                  | (((~n0a7cmohxqtifv1u_wo) | (~gefz7vdqfjfmc7vx9p)) & ek78h0rdvr2jbnet5d  )
                  | (((~n0a7cmohxqtifv1u_wo) | (~gefz7vdqfjfmc7vx9p)) & xiv4a67_96psl3rnqmp )
                  | (((~jo9y8uxpmti4rhw6z) | (~gn663w5srr2mzrtvg)) & u62i7sw55i0ixtfn  )
                  | (((~jo9y8uxpmti4rhw6z) | (~gn663w5srr2mzrtvg)) & wrwhm830pc1woxrw )
                  | (((~h_cfdp023jzvo4byhlbh) | (~ed8kepqzl3lj7rms5l)) & b1u7q1bl0kcxqkk9lh  )
                  | (((~h_cfdp023jzvo4byhlbh) | (~ed8kepqzl3lj7rms5l)) & cdtdn0g9ejv3kd5b )

                  | s32nr2e9a6f4hrqy4n775or 
                 )
               ;



  assign gjyhd0u2t3wy11drm07 = um1_bmln_sf2i4vzbya_ | yryyg8udb_4akvy;
  assign e280ym1w614qoep160njy = i72_qcuo70vljgkcb0fbj;
  assign an0s8c6hcabd901wob_8zo = y8_gkxsfle & (~pydatzxqqi) & el7_p8jit09 &  
                   
                   
               ( 
                    ((~rby_e01aj9mayt) & f3nolyi4jv6dte        )
                  | ((~rby_e01aj9mayt) & exvzt_vf1mmht       )
                  | ((~wy3w2aq98iuq6w) & e_kz098g         )
                  | ((~wy3w2aq98iuq6w) & n0hf68fqn6tl        )
                  | ((~x6zcn2iwg4w04) & h0m0j6wupakd3zh      )
                  | ((~x6zcn2iwg4w04) & di0_fvfp1wszdubcc     )
                  | ((~edebxw2_52r74i4yub5n)  & w4w2ra2eqzikjlg  )
                  | ((~edebxw2_52r74i4yub5n)  & ibihcuxenb1h85msj )
                  | ((~n0a7cmohxqtifv1u_wo)  & ek78h0rdvr2jbnet5d  )
                  | ((~n0a7cmohxqtifv1u_wo)  & xiv4a67_96psl3rnqmp )
                  | ((~jo9y8uxpmti4rhw6z)  & u62i7sw55i0ixtfn  )
                  | ((~jo9y8uxpmti4rhw6z)  & wrwhm830pc1woxrw )
                  | ((~h_cfdp023jzvo4byhlbh)  & b1u7q1bl0kcxqkk9lh  )
                  | ((~h_cfdp023jzvo4byhlbh)  & cdtdn0g9ejv3kd5b )

                  | s32nr2e9a6f4hrqy4n775or 
                 )
               ;


endmodule




















module ihs34rgb4pudd03(
  input xoauecm4__2ehfjw,
  input [64-1:0] vf5xcr67bqhzlo43_,

  input atqel3v0fzjjsz,
  output [64-1:0] wuke41p8s ,
  output hk9dhg3ue,

  input  dk2xhkj77a,
  input  ru_wi

  );


  wire [64-1:0] s6er21uf;
  wire l4ylal_gzpjxcqxv = ((s6er21uf == (~(64'b0))));
  wire t_fdz268gdu4    = xoauecm4__2ehfjw    |
                      (~atqel3v0fzjjsz)
                      ;
  
  wire [64-1:0] qd_0tqy7a    = xoauecm4__2ehfjw    ? vf5xcr67bqhzlo43_ : (s6er21uf  + {{64-1{1'b0}},1'b1});

  
  ux607_gnrl_dfflr #(64) pyjjf7_txbyb (t_fdz268gdu4, qd_0tqy7a, s6er21uf   , dk2xhkj77a, ru_wi);
  assign wuke41p8s    = s6er21uf;



  
  
  assign hk9dhg3ue = 1'b1
                     & l4ylal_gzpjxcqxv 
                     & (~xoauecm4__2ehfjw)
                     & (~atqel3v0fzjjsz)
                     ;

endmodule









































module whvqleuvihduw(

  input           gf33atgy,
  input           ru_wi,

  input           th06du2c8e2_b7k,
  output          irjoi8wvo25u209f_5,
  input  [32-1:0] zvk11dhgg2s67mkq, 
  input           zxe59xihintdqfy9d, 
  input  [32-1:0] u4r4b_6kp09q767q,

  output          klkflmsyyf5w7ar,
  input           wy36iirxspfw56864,
  output [32-1:0] h7f6k_ims_9p3,

  output          iqg2bp31t,
  output          gf9zfb8tq9sv,
  output          de1sbr3kjbswue, 


  output [32-1:0] olks1id,  
  output [32-1:0] rhpeh82g, 
  output          swohhsf_wlqj,
  output          f9xsdhw9rmwvtyi,

  input           v384utu4po2
);

  localparam zgwo0o2mbyu_fw7k_ci      = 16'hFFC     ;
  localparam vphttp38yp4             = 16'hFF8            ;
  localparam sx1illxej8b4gdl0at1    = 16'h0   ;
  localparam mq7bykaoqmzd0717wdpoi1v3    = 16'h4   ;
  localparam q0h8q2b3r95d_5vzxnc8rj = 16'h8;
  localparam rj1eq4aawwhd0p15saq2u04yu = 16'hC;
  localparam vmy0082birsmo98           = 16'hFF0          ;

  localparam wiw59xg5m2b8rigm6xnr5xpz      = 16'h1000     ;
  localparam r25qkppgc1vzeas4nxisqa65ef    = 16'hCFF8   ;
  localparam mb7e3axg90hck330t24hvmv    = 16'hCFFC   ;
  localparam imf7pim20ydr6h7en5gkymf_97 = 16'h5000;
  localparam x5ippqzy6szbaay_dr0ltreuiu3vp = 16'h5004;

  wire h5maomnmovgqtb7    = th06du2c8e2_b7k & irjoi8wvo25u209f_5;
  wire fz_isl8q3blzlbl2zzf = h5maomnmovgqtb7 & (~zxe59xihintdqfy9d); 
  wire dh1lon9y8avka453f7vc = h5maomnmovgqtb7 & zxe59xihintdqfy9d; 


  wire rbdq13ad1iflzgcxt      = (zvk11dhgg2s67mkq[16-1:0] == zgwo0o2mbyu_fw7k_ci)
                         | (zvk11dhgg2s67mkq[16-1:0] == wiw59xg5m2b8rigm6xnr5xpz)
                         ;
  wire itfo45nl8ccl9ho6anqy = (zvk11dhgg2s67mkq[16-1:0] == q0h8q2b3r95d_5vzxnc8rj)
                         | (zvk11dhgg2s67mkq[16-1:0] == imf7pim20ydr6h7en5gkymf_97)
                         ;
  wire fyv92axrq_nqf47o8p8p = (zvk11dhgg2s67mkq[16-1:0] == rj1eq4aawwhd0p15saq2u04yu)
                         | (zvk11dhgg2s67mkq[16-1:0] == x5ippqzy6szbaay_dr0ltreuiu3vp)
                         ;
  wire rxhdmd1_iqvdqy8s    = (zvk11dhgg2s67mkq[16-1:0] == sx1illxej8b4gdl0at1)
                         | (zvk11dhgg2s67mkq[16-1:0] == r25qkppgc1vzeas4nxisqa65ef)
                         ;
  wire lq2ijol665jfql_    = (zvk11dhgg2s67mkq[16-1:0] == mq7bykaoqmzd0717wdpoi1v3)
                         | (zvk11dhgg2s67mkq[16-1:0] == mb7e3axg90hck330t24hvmv)
                         ;
  wire u5tgrjl_vkffwc      = (zvk11dhgg2s67mkq[16-1:0] == vphttp38yp4);
  wire ftzkpyxxdu0xw56   = (zvk11dhgg2s67mkq[16-1:0] == vmy0082birsmo98);



  wire [32-1:0] y7hno0     ;
  wire [32-1:0] bci8vm0     ;
  wire [32-1:0] z30tlpe25_l;
  wire [32-1:0] zwoqlvqk974w;
  wire          rri79w57er4mc  ;

  wire [32-1:0] vf_r9hn9ty7axn = 
                     ({32{rbdq13ad1iflzgcxt     }} & y7hno0     )
                   | ({32{u5tgrjl_vkffwc     }} & bci8vm0     )
                   | ({32{itfo45nl8ccl9ho6anqy}} & z30tlpe25_l)
                   | ({32{fyv92axrq_nqf47o8p8p}} & zwoqlvqk974w)
                   | ({32{rxhdmd1_iqvdqy8s   }} & olks1id   )
                   | ({32{lq2ijol665jfql_   }} & rhpeh82g   )
                   | ({32{ftzkpyxxdu0xw56  }} & {rri79w57er4mc,31'b0});




  wire [32-1:0] owhv15w4y;
  wire x39yugtyz_ = fz_isl8q3blzlbl2zzf & u5tgrjl_vkffwc;
  assign owhv15w4y = {29'b0, u4r4b_6kp09q767q[2:0]};
  ux607_gnrl_dfflr #(32) bc6y97yaexc(x39yugtyz_, owhv15w4y, bci8vm0, gf33atgy, ru_wi);

  assign swohhsf_wlqj = bci8vm0[0];
  wire   oukjr0g0mvt9x5_b = bci8vm0[1];
  assign f9xsdhw9rmwvtyi = bci8vm0[2];



  wire [32-1:0] s0z0trof9;
  wire o9mswcyrhfg = fz_isl8q3blzlbl2zzf & rbdq13ad1iflzgcxt;
  assign s0z0trof9 = {31'b0, u4r4b_6kp09q767q[0]};
  ux607_gnrl_dfflr #(32) eq8wikscsg5(o9mswcyrhfg, s0z0trof9, y7hno0, gf33atgy, ru_wi);

  assign gf9zfb8tq9sv = y7hno0[0];


  wire [32-1:0] meexm9i6bxn817wfl;
  wire [32-1:0] cmx9w5jaxnxitrwy;

  wire [32-1:0] x81cfbipkcmhbrc;
  wire dpn69ps2tdrv88 = fz_isl8q3blzlbl2zzf & rxhdmd1_iqvdqy8s;
  wire ekm_hx_g545 = v384utu4po2;
  wire omast0gdm271p = oukjr0g0mvt9x5_b & iqg2bp31t;
  wire ftn8negiuj4cay = dpn69ps2tdrv88 | ekm_hx_g545 | omast0gdm271p;
  assign x81cfbipkcmhbrc = omast0gdm271p ? 32'b0 : dpn69ps2tdrv88 ? u4r4b_6kp09q767q : meexm9i6bxn817wfl;
  ux607_gnrl_dfflr #(32) crhtbc0l4ffy6(ftn8negiuj4cay, x81cfbipkcmhbrc, olks1id, gf33atgy, ru_wi);



  wire [32-1:0] w85m2_8h5lnk8;
  wire e9jryho67z9v = fz_isl8q3blzlbl2zzf & lq2ijol665jfql_;
  wire okwx10__iw = v384utu4po2;
  wire fa_idem1me0hmvv = omast0gdm271p;
  wire ckbztq1ujez9c = e9jryho67z9v | okwx10__iw | fa_idem1me0hmvv;
  assign w85m2_8h5lnk8 = fa_idem1me0hmvv ? 32'b0 : e9jryho67z9v ? u4r4b_6kp09q767q : cmx9w5jaxnxitrwy;
  ux607_gnrl_dfflr #(32) ptj04z8i2bigsylb_(ckbztq1ujez9c, w85m2_8h5lnk8, rhpeh82g, gf33atgy, ru_wi);




  assign {cmx9w5jaxnxitrwy, meexm9i6bxn817wfl} = {rhpeh82g, olks1id} + 64'b1;







  wire [32-1:0] fbapnnhj2hy97;
  wire ol94nll6c7s5n3fi = fz_isl8q3blzlbl2zzf & itfo45nl8ccl9ho6anqy;
  wire ej2q30w47kt2zc = ol94nll6c7s5n3fi;
  assign fbapnnhj2hy97 = u4r4b_6kp09q767q;

  ux607_gnrl_dfflrs #(32) rz013tx7y9mqx99afl3(ej2q30w47kt2zc, fbapnnhj2hy97, z30tlpe25_l, gf33atgy, ru_wi);



  wire [32-1:0] z4i7kceklhm_ozy0fk;
  wire fjkpradyunbjdkx5 = fz_isl8q3blzlbl2zzf & fyv92axrq_nqf47o8p8p;
  wire yen1vpxa06lib = fjkpradyunbjdkx5;
  assign z4i7kceklhm_ozy0fk = u4r4b_6kp09q767q;

  ux607_gnrl_dfflrs #(32) bf7xn1dyo9emrt8h(yen1vpxa06lib, z4i7kceklhm_ozy0fk, zwoqlvqk974w, gf33atgy, ru_wi);



  wire wtrj_xr_9ig73h;
  wire srrb8cjprkuezz = fz_isl8q3blzlbl2zzf & (u4r4b_6kp09q767q == 32'h80000a5f) & ftzkpyxxdu0xw56;
  wire z0nap6fndmfzxkik = srrb8cjprkuezz; 
  assign  wtrj_xr_9ig73h = srrb8cjprkuezz;
  ux607_gnrl_dfflr #(1) jkicwazwrw5dz6v9f(z0nap6fndmfzxkik, wtrj_xr_9ig73h, rri79w57er4mc, gf33atgy, ru_wi);

  assign iqg2bp31t = ({rhpeh82g, olks1id} >= {zwoqlvqk974w, z30tlpe25_l});
  assign de1sbr3kjbswue = rri79w57er4mc;


  assign klkflmsyyf5w7ar = th06du2c8e2_b7k;
  assign irjoi8wvo25u209f_5 = wy36iirxspfw56864;
  assign h7f6k_ims_9p3 = vf_r9hn9ty7axn;


endmodule























module ux607_tmr_top(
  output  tmr_active,
  input   clk_aon,
  input   clk,

  input   rst_n,

  input           i_icb_cmd_valid,
  output          i_icb_cmd_ready,
  input  [32-1:0] i_icb_cmd_addr, 
  input           i_icb_cmd_read, 
  input  [32-1:0] i_icb_cmd_wdata,
  input  [4 -1:0] i_icb_cmd_wmask,


  input           i_icb_cmd_mmode,
  input           i_icb_cmd_smode,
  input           i_icb_cmd_dmode, 

  output          i_icb_rsp_valid,
  input           i_icb_rsp_ready,
  output [32-1:0] i_icb_rsp_rdata,
  output          i_icb_rsp_err,

  output [31:0]   mtime,
  output [31:0]   mtimeh,

  output  tmr_irq,
  output  sft_irq,
  output  sft_rst_req,

  input   rtc_toggle_a,

  input   dbg_stoptime 
);

  wire          swohhsf_wlqj; 
  wire          f9xsdhw9rmwvtyi;

  wire          klkflmsyyf5w7ar;
  wire          wy36iirxspfw56864;
  wire [32-1:0] h7f6k_ims_9p3;

     
  assign wy36iirxspfw56864   = i_icb_rsp_ready;
  assign i_icb_rsp_valid = klkflmsyyf5w7ar;
  assign i_icb_rsp_rdata = h7f6k_ims_9p3;


  wire t_o10omz8u1qas6 = swohhsf_wlqj | dbg_stoptime;

  wire yjbgz3d9idgo15x6;

  ux607_gnrl_sync # (
  .DP(2),
  .DW(1)
  ) wfnbvh7mhj0x113sg(
      .din_a    (rtc_toggle_a),
      .dout     (yjbgz3d9idgo15x6),
      .clk      (clk_aon     ),
      .rst_n    (rst_n) 
  );


  wire hbstxas6ddt1 = yjbgz3d9idgo15x6;


  wire zd6jck3utr = hbstxas6ddt1 & (~t_o10omz8u1qas6);

  wire f17rj5pr; 

  ux607_gnrl_dffr #(1) t1d_mpleop2p (zd6jck3utr, f17rj5pr, clk_aon, rst_n);
  wire sgq8uw3gw03 = zd6jck3utr ^ f17rj5pr; 
  wire wz7x7tls = f9xsdhw9rmwvtyi ? (~t_o10omz8u1qas6) : sgq8uw3gw03;


  whvqleuvihduw  je6a0d77jwuf6fox99(

  .gf33atgy             (clk),
  .ru_wi           (rst_n  ),

  .th06du2c8e2_b7k   (i_icb_cmd_valid), 
  .irjoi8wvo25u209f_5   (i_icb_cmd_ready),
  .zvk11dhgg2s67mkq    (i_icb_cmd_addr ),
  .zxe59xihintdqfy9d    (i_icb_cmd_read ),
  .u4r4b_6kp09q767q   (i_icb_cmd_wdata),

  .klkflmsyyf5w7ar   (klkflmsyyf5w7ar),
  .wy36iirxspfw56864   (wy36iirxspfw56864),
  .h7f6k_ims_9p3   (h7f6k_ims_9p3),

  .olks1id         (mtime),
  .rhpeh82g        (mtimeh),
  .swohhsf_wlqj        (swohhsf_wlqj), 
  .f9xsdhw9rmwvtyi      (f9xsdhw9rmwvtyi),

  .gf9zfb8tq9sv         (sft_irq),
  .de1sbr3kjbswue     (sft_rst_req),
  .iqg2bp31t         (tmr_irq),
  .v384utu4po2      (wz7x7tls) 

  );

  assign tmr_active = i_icb_cmd_valid | i_icb_rsp_valid |  klkflmsyyf5w7ar |
                     ((~t_o10omz8u1qas6) & wz7x7tls);
  assign i_icb_rsp_err = 1'b0;

endmodule




















module zu3cpta_6amki_tj3nyfxw7 (

  input [64-1:0]  x6eruzvd5,

  
  

  input j2f1_e0en,
  input aw82i964do,
  input y8_gkxsfle,

  input kw2010ymt1iz5,
  input yeo38qe8mley55,
  input rvfxw53dft5,
  input r6dop3ru22,
    
  input [64*4-1:0] n6a0r_0zddzrme8,
  input [64*4-1:0] azll7rq5fab5ou,

  output coeuovgdaw1,
  output o_gen1so7__xgr3pw2,

  input gf33atgy,
  input ru_wi
  );

  
  wire [64-1:0] chp26_u95[0:4-1];
  wire [64-1:0] t6smjlrvsmz9cf[0:4-1];
  wire [64-1:0] ra_jg19sao28hcbk40imc3[0:4-1];
  
  wire [64-1:0] oozxn9oahfs[0:4-1];

  wire [4-1:0] rex4gxxixhigl;
  wire [4-1:0] uwmh9ibjhdww9lx;
  wire [4-1:0] rffq00v3nls9;
  wire [4-1:0] szhb198zgi;
  wire [4-1:0] xnmuifu1k94;
  wire [4-1:0] posoetp4resy;
  wire [4-1:0] es08_js9uv3;
  wire [4-1:0] yww0wmwdmuor__;
  wire [4-1:0] dyjl_ygidv1sb_ewz;
  wire [4-1:0] fe_ct99wyw3xf8zk;
  wire [4-1:0] o5_eyxx7i0cpwlmz;
  wire [6-1:0] rl3eibl4dzj7qma [4-1:0];
  wire [4-1:0] p0c8tgdma7gpbo_z0s;
  wire [4-1:0] ajb9pmoqwq8m;
  wire [4-1:0] rwdtxow9zmnysx;
  wire [4-1:0] xzfghka20fqvcz8ejsb;
  wire [4-1:0] qnnetqriq5ujaq2p8lz;
  wire [4-1:0] i7yzy90dwot7yv4aps135gip;
  wire [64-1:0] vfcxvf6all4svq [4-1:0];
  wire [64-1:0] n0qo9nodyynt [4-1:0];
  wire [64-1:0] e3ibtx9ft7rgyhl39za [4-1:0];
  wire [64-1:0] yzuopx8dmcz [4-1:0];

  wire [4-1:0] v87q0gcwk;
  wire [4-1:0] ngarog4ifb;

  
  
  


  genvar i;
  genvar j;

  generate 
  for(i=0; i<4; i=i+1) begin: v2qtfc2yoa 
      
    assign chp26_u95[i] = n6a0r_0zddzrme8[64*i +: 64]; 
    assign oozxn9oahfs[i] = azll7rq5fab5ou[64*i +: 64]; 


    assign rex4gxxixhigl [i] = oozxn9oahfs[i][0];
    assign uwmh9ibjhdww9lx [i] = oozxn9oahfs[i][1];
    assign rffq00v3nls9 [i] = oozxn9oahfs[i][2];
    assign szhb198zgi  [i] = oozxn9oahfs[i][3];
    assign xnmuifu1k94  [i] = oozxn9oahfs[i][4];
    assign posoetp4resy  [i] = oozxn9oahfs[i][6];
    assign dyjl_ygidv1sb_ewz [i] = (oozxn9oahfs[i][10:7] == 4'd0);
    assign fe_ct99wyw3xf8zk [i] = (oozxn9oahfs[i][10:7] == 4'd1);
    assign o5_eyxx7i0cpwlmz [i] = oozxn9oahfs[i][11];
    assign es08_js9uv3[i] = (oozxn9oahfs[i][17:12] == 6'd1);
    assign yww0wmwdmuor__[i] = (oozxn9oahfs[i][59]);
    assign rl3eibl4dzj7qma [i] = oozxn9oahfs[i][64-6:64-11];
    assign p0c8tgdma7gpbo_z0s[i] = (oozxn9oahfs[i][64-1:64-4] == 4'd2);

      
      
    assign vfcxvf6all4svq[i] = ~(64'b0);

      
      
      
      
      
      
      
      
      
      
      
      
      
      

    assign t6smjlrvsmz9cf[i] = {chp26_u95[i][64-2:0], 1'b1};
    assign ra_jg19sao28hcbk40imc3[i] = (~t6smjlrvsmz9cf[i]);
    for(j=0; j<64; j=j+1) begin: vxbvrafws 
      
        assign e3ibtx9ft7rgyhl39za[i][j] = |ra_jg19sao28hcbk40imc3[i][j:0]; 
    end
      
    assign n0qo9nodyynt[i] = {{(64-12){1'b1}}, e3ibtx9ft7rgyhl39za[i][11:0]};

    assign yzuopx8dmcz[i] = dyjl_ygidv1sb_ewz[i] ?  vfcxvf6all4svq[i] :
                           fe_ct99wyw3xf8zk[i] ?  n0qo9nodyynt[i] :
                                                (~(64'h0));
    
    
    


    assign ajb9pmoqwq8m[i] = (dyjl_ygidv1sb_ewz[i] |  fe_ct99wyw3xf8zk[i]) & 
                           ((x6eruzvd5 & yzuopx8dmcz[i][64-1:0]) == (chp26_u95[i][64-1:0] & yzuopx8dmcz[i][64-1:0])); 

    assign xzfghka20fqvcz8ejsb[i] = ( 
                           (p0c8tgdma7gpbo_z0s[i] & rex4gxxixhigl[i] & (kw2010ymt1iz5 | rvfxw53dft5)) 
                         | (p0c8tgdma7gpbo_z0s[i] & uwmh9ibjhdww9lx[i] & (yeo38qe8mley55 | rvfxw53dft5)) 
                         | (p0c8tgdma7gpbo_z0s[i] & rffq00v3nls9[i] & (r6dop3ru22)) 
                         );

    assign rwdtxow9zmnysx[i] = (aw82i964do ? posoetp4resy[i] : y8_gkxsfle ? xnmuifu1k94[i] : szhb198zgi[i])  & xzfghka20fqvcz8ejsb[i];

    assign qnnetqriq5ujaq2p8lz[i] = ajb9pmoqwq8m[i] & rwdtxow9zmnysx[i];

    assign i7yzy90dwot7yv4aps135gip[i] =   qnnetqriq5ujaq2p8lz[i];
    assign v87q0gcwk[i]   =   es08_js9uv3[i]  & i7yzy90dwot7yv4aps135gip[i] 
                          
                          & yww0wmwdmuor__[i];
    assign ngarog4ifb[i] = (~es08_js9uv3[i]) & i7yzy90dwot7yv4aps135gip[i];

  end
  endgenerate

  assign coeuovgdaw1   = (~j2f1_e0en) & (|v87q0gcwk);
  assign o_gen1so7__xgr3pw2 = (~j2f1_e0en) & (|ngarog4ifb);


endmodule





















module qy_752rpwt4qqgs1gejira_te (
    
  input [64*4-1:0] azll7rq5fab5ou,

  input  j2f1_e0en,
  input  aw82i964do,
  input  y8_gkxsfle,

  output dd8pb3i1ec_uv5,
  output s62ahm8e0we20r 
  );

  
  wire [64-1:0] dwt4xr7nj[0:4-1];

  wire [4-1:0] szhb198zgi;
  wire [4-1:0] xnmuifu1k94;
  wire [4-1:0] posoetp4resy;
  wire [4-1:0] es08_js9uv3;
  wire [4-1:0] wg0v_ml1wpp72y;
  wire [4-1:0] yww0wmwdmuor__;
  wire [4-1:0] cgrmm8bl47usi_c58ak5;

  wire [4-1:0] nag3soi;
  wire [4-1:0] v87q0gcwk;
  wire [4-1:0] ngarog4ifb;

  genvar i;

  generate 
  for(i=0; i<4; i=i+1) begin: v2qtfc2yoa 
      
    assign dwt4xr7nj[i] = azll7rq5fab5ou[64*i +: 64]; 


    assign es08_js9uv3[i] = (dwt4xr7nj[i][5:0] == 6'd1);
    assign szhb198zgi  [i] = dwt4xr7nj[i][6];
    assign xnmuifu1k94  [i] = dwt4xr7nj[i][7];
    assign posoetp4resy  [i] = dwt4xr7nj[i][9];
    assign wg0v_ml1wpp72y  [i] = dwt4xr7nj[i][10];
    assign yww0wmwdmuor__  [i] = dwt4xr7nj[i][59];
    assign cgrmm8bl47usi_c58ak5[i] = (dwt4xr7nj[i][64-1:64-4] == 4'd3);


    assign nag3soi[i] = (aw82i964do ? posoetp4resy[i] : y8_gkxsfle ? xnmuifu1k94[i] : szhb198zgi[i]) & 
                      cgrmm8bl47usi_c58ak5[i]   
                      
                      ;


    assign v87q0gcwk[i]   =   es08_js9uv3[i]  & nag3soi[i] 
                          
                          & yww0wmwdmuor__[i];
    assign ngarog4ifb[i] = (~es08_js9uv3[i]) & nag3soi[i];

  end
  endgenerate

  assign dd8pb3i1ec_uv5   = (~j2f1_e0en) & (|v87q0gcwk);
  assign s62ahm8e0we20r = (~j2f1_e0en) & (|ngarog4ifb);


endmodule





















module vx6hu6m3c9ub1xbqu6okmcqh6_ (
  input j2f1_e0en,
  input aw82i964do,
  input y8_gkxsfle,

  input dn8riluj40uunvq5,

  input [4:0] hh49o83xz9_uu,
  input [9:0] g1fa4tixb,

  input lmu064oe20,
  input qemnpyvmwrt,

    
  input [64*4-1:0] n6a0r_0zddzrme8,
  input [64*4-1:0] azll7rq5fab5ou,

  output coeuovgdaw1,
  output o_gen1so7__xgr3pw2 

  );

  
  wire [64-1:0] chp26_u95[0:4-1];
  
  wire [64-1:0] oozxn9oahfs[0:4-1];

  wire [4-1:0] es08_js9uv3;
  wire [4-1:0] szhb198zgi;
  wire [4-1:0] xnmuifu1k94;
  wire [4-1:0] posoetp4resy;
  wire [4-1:0] ex9hadotf0v6i96xrt;
  wire [4-1:0] wpmkxis2ol1jrqrwjo;
  wire [4-1:0] bgnys0xjuky70;
  wire [4-1:0] wu4wg9dj1dkxuk5;
  wire [4-1:0] jy904cz9x4dnfxmti9ek0;
  wire [4-1:0] t50ns65cya9amnkw;
  wire [4-1:0] sn1ikupg_0fn254crskt;
  wire [4-1:0] bihvo853v2swpd_w;
  wire [4-1:0] yww0wmwdmuor__;

  wire [4-1:0] v87q0gcwk;
  wire [4-1:0] ngarog4ifb;
  wire [4-1:0] nag3soi;

  genvar i;

  generate 
  for(i=0; i<4; i=i+1) begin: v2qtfc2yoa 
      
    assign chp26_u95[i] = n6a0r_0zddzrme8[64*i +: 64]; 
    assign oozxn9oahfs[i] = azll7rq5fab5ou[64*i +: 64]; 


    assign es08_js9uv3[i] = (oozxn9oahfs[i][5:0] == 6'd1);
    assign szhb198zgi  [i] = oozxn9oahfs[i][6];
    assign xnmuifu1k94  [i] = oozxn9oahfs[i][7];
    assign posoetp4resy  [i] = oozxn9oahfs[i][9];

    assign ex9hadotf0v6i96xrt[i] = (oozxn9oahfs[i][64-1:64-4] == 4'd4);
    assign wpmkxis2ol1jrqrwjo[i] = (oozxn9oahfs[i][64-1:64-4] == 4'd5);

    assign yww0wmwdmuor__  [i] = oozxn9oahfs[i][59];

    assign bgnys0xjuky70[i] = chp26_u95[i][hh49o83xz9_uu]; 


    
    
    
    
    
    assign jy904cz9x4dnfxmti9ek0[i] = chp26_u95[i][g1fa4tixb[4:0]]; 

    assign sn1ikupg_0fn254crskt[i] = chp26_u95[i][0]  & (chp26_u95[i][10:1]  == g1fa4tixb); 
    assign bihvo853v2swpd_w[i] = chp26_u95[i][16] & (chp26_u95[i][26:17] == g1fa4tixb); 

    assign t50ns65cya9amnkw[i] = (sn1ikupg_0fn254crskt[i] | bihvo853v2swpd_w[i]);

    assign wu4wg9dj1dkxuk5[i] = dn8riluj40uunvq5 ? t50ns65cya9amnkw[i] : jy904cz9x4dnfxmti9ek0[i];


    assign nag3soi[i] = (aw82i964do ? posoetp4resy[i] : y8_gkxsfle ? xnmuifu1k94[i] : szhb198zgi[i]) & ( 
                         | (ex9hadotf0v6i96xrt[i] & qemnpyvmwrt & wu4wg9dj1dkxuk5[i]) 
                         | (wpmkxis2ol1jrqrwjo[i] & lmu064oe20 & bgnys0xjuky70[i]) 
                         );

    assign v87q0gcwk[i]   =   es08_js9uv3[i]  & nag3soi[i] 
                          
                          & yww0wmwdmuor__[i];
    assign ngarog4ifb[i] = (~es08_js9uv3[i]) & nag3soi[i];

  end
  endgenerate

  assign coeuovgdaw1   = (~j2f1_e0en) & (|v87q0gcwk);
  assign o_gen1so7__xgr3pw2 = (~j2f1_e0en) & (|ngarog4ifb);


endmodule





























module n9qdnl9_3k0n2m1yo4pxt(
  input                                   ru_wi,
  input                                   gf33atgy,

  input                                   g3ljqli3ukatw2132ssx,
  
  input                                   fkuqlh34r,
  input [16-1:0]            hnc10arn_rd,
  input                                   rm1dxjejhq7dh3q5m,
  input [1:0]                             st2zalpx0uf,
  input                                   ni01kj42oob2x,
  input                                   ah8kjlmvnaxzbi,
  input [1:0]                             toox2fc0snvsr_n,                        
  
  
  
  output                                  f_yktlpn8eslyt9akam,
  output                                  lf2bvnvn_k5yqtn5od,
  output                                  vy13vm0dqfvofi_2dp09,
  output                                  klkyy__rhf1ui9omvg,
  output [66-1:0]       wqhbmg7dvocz1j9wy9,
  output [66-1:0]       tp8gw47qpcwgagtuvei,
  output [6-1:0]      jw_o9pbzjnqwneo0t,
  input  [66-1:0]       qbksws8auoc48qp3sb,
  input  [66-1:0]       xyeddoohku7q6ja9pvnp,
  
  
  
  input                                   kbi8qdl8tmgm5j0uu1p1xu0, 
  input                                   on37whxvtxni09my52drx, 
  input                                   ntychvakx3t8mzzgh8_ev, 
  input [27-1:0]            k11nc9vg2x3_cg_semdn, 
  input [27-1:0]            y0__7wpxqx83r42pl, 
 

  output                                  w9_jhj6c4a6df_4pxyyb,
  output [55-1:0]      oh3gt3hus6shq_f5p7d,
  output                                  zs5xuhg0c8f60zy_nv1v987v74,
  
  
  output                                  ezhgcskig85uffd7xor0c,
  output [51-1:0]      tbassexmaytz0vwwh79gt,
  output                                  ibq_47zipoy6cbbw2uwa2jy_1o,
  
  
  output                                  nvupfco9fb64lzc1ej,
  output                                  hi_bckth818lxu0y4nnr6xzf,

  output                                  xhehq_1td3fs,                        
  output                                  m0rgjbiqu6nadc33k5,
  
  
  
  input                                   m01i4z2a2meu,
  input                                   mou2g2qz02878jxn,
  input                                   yyz7lhabpe7x17h10y,
  input [16-1:0]            j3d84gxpt2b4pd8,
  output                                  ew6x7412r46,
  
  
  
  
  
  input                                   b3ymasxx4cnt,
  input                                   pffig1fl4xtnw,
  input                                   j48quvipiuwft,
  input                                   rxosbn3wj_1o6y20fv,
  input                                   w90yio82brq3k1uvzp57esy,
  input                                   kbv_rf0mvydplzwef_3qe,

  input [20-1:0]              kpl3digtonftoyh,
  input [1:0]                             ermcr77dq4jhq99jq,
  input                                   mnac5hr2jmri8kx5xj,
  input                                   o44hlt5z77imds2,
  input                                   he47fcvawyr15g,
  input                                   oclzmsyeij5bw,
  input                                   vv_afyrrunvcjbtl2_,
  input                                   n9qmjt3s04yv75d,
  input                                   cf1ozmszcxohbmdmqv,


  
  output [27-1:0]           uhegwov_bgw,
  output                                  b0l_kaqp,
  output                                  tlygxd1cs0w,
  output                                  i3o6jvv3t7i,
  output                                  xwd9yye9seo2l,
  
  output                                  d4ab_e8ynn1a53_52a3
  
  );
 

   
  wire sd4rdwq_5i7fe5;
  
  wire c4ughu0qm5sfai;
  ux607_gnrl_dffrs #(1) dbvgqgz185u8yqz4kvb4g ( 1'b0, c4ughu0qm5sfai, gf33atgy, ru_wi);
  
  wire ld42chldsdyksa9;
  wire t523n0nf23b9vzzq = (~ld42chldsdyksa9) & c4ughu0qm5sfai & (~g3ljqli3ukatw2132ssx);
  wire sr1rrv8mkq8ype = ld42chldsdyksa9 & sd4rdwq_5i7fe5;
  wire y2xlaa97t8eslcu1e = t523n0nf23b9vzzq | sr1rrv8mkq8ype;
  wire mk7m52sz5niya27 = t523n0nf23b9vzzq | ~sr1rrv8mkq8ype;
  ux607_gnrl_dfflr #(1) jwi0n6alhl8fjgnpgos (y2xlaa97t8eslcu1e, mk7m52sz5niya27, ld42chldsdyksa9, gf33atgy, ru_wi);

  wire x3h2m98yhzqwpra5q0q = ld42chldsdyksa9;

  
  localparam l4e4x5iuocpq14dam9ucku = 3;
  
  wire [l4e4x5iuocpq14dam9ucku-1:0] v0qy_p3s0bq9bqj0mz;
  wire [l4e4x5iuocpq14dam9ucku-1:0] q5xw1oq2dyd3_r9;
  wire e8ay6vzax1puil9e;
  ux607_gnrl_dfflr #(l4e4x5iuocpq14dam9ucku) bcvq19zb8g2rn0m33r4 (e8ay6vzax1puil9e, v0qy_p3s0bq9bqj0mz, q5xw1oq2dyd3_r9, gf33atgy, ru_wi);


  localparam klcv32s524noj675s         = 3'd0;
  localparam qi8j2njkyk3a22m95kc8jquq       = 3'd1;
  localparam ai81jjukhk7_uoovfndq690s   = 3'd2;
  localparam x2yiem7xqi4jww3op6siel        = 3'd3;
  localparam r_h500kxshad5gkq4zgdswta      = 3'd4;
  localparam qka__s7my8mvb4j5dhd071      = 3'd5;
  localparam iosvpnl0hccumt4jze71nkq0d    = 3'd6;
  localparam ghxu50th5tej1yhl8zrb7lticj     = 3'd7;
  
  
  wire [l4e4x5iuocpq14dam9ucku-1:0] u99tnldu986760c5;
  wire [l4e4x5iuocpq14dam9ucku-1:0] nhzryulpguznnnqmzgn0;
  wire [l4e4x5iuocpq14dam9ucku-1:0] jlnkd6qhsmjqw47tf1t64byci;
  wire [l4e4x5iuocpq14dam9ucku-1:0] s67r7tvcckkpgs9;
  wire [l4e4x5iuocpq14dam9ucku-1:0] x4lgrwp6fc79b0ehv9;
  wire [l4e4x5iuocpq14dam9ucku-1:0] dbw_jljmitz3e_zmp;
  wire [l4e4x5iuocpq14dam9ucku-1:0] u9fc6nt5deod0x3wvfv;
  wire [l4e4x5iuocpq14dam9ucku-1:0] v0gpnd2kvonwrxb2d1;
  
  wire wfoen161d4r42bkqp34lj;
  wire dqc3ngr_5saws_sp75dkhv;
  wire wd2v3s292zarv6r_qtszoymxjmnb9b;
  wire igbfek2f8xd5vcozwc6mvu;
  wire kqoce2mai7legb67b3_l3ofi1v;
  wire mqxidx634c8oo3gea0__8s;
  wire vr63zqx6y0ffx32ubvl670vs9m6qf;
  wire wydnyq82nhj8gfglsmtj8ffh;
  
  wire fi5j2nq20y39ylylwhs         = (q5xw1oq2dyd3_r9 == klcv32s524noj675s      );
  wire vikfdhomdfhf7ewfaitsy_gj       = (q5xw1oq2dyd3_r9 == qi8j2njkyk3a22m95kc8jquq    );
  wire fpsdt9vdjcwssz9tezden07r7   = (q5xw1oq2dyd3_r9 == ai81jjukhk7_uoovfndq690s);
  wire b7z98rnx88w42eg6952nx8x        = (q5xw1oq2dyd3_r9 == x2yiem7xqi4jww3op6siel     );
  wire nme7un7hr7uwq6h4qmctk_srkw      = (q5xw1oq2dyd3_r9 == r_h500kxshad5gkq4zgdswta   );
  wire d3o9i8v1m3g16rvwhai2wh7      = (q5xw1oq2dyd3_r9 == qka__s7my8mvb4j5dhd071   );
  wire qhcnhctsg82wxcyhu80cuex4c    = (q5xw1oq2dyd3_r9 == iosvpnl0hccumt4jze71nkq0d );
  wire oadttvx13julmicav817mtk5jev     = (q5xw1oq2dyd3_r9 == ghxu50th5tej1yhl8zrb7lticj  );
  
  assign e8ay6vzax1puil9e = wfoen161d4r42bkqp34lj
                          | dqc3ngr_5saws_sp75dkhv
                          | wd2v3s292zarv6r_qtszoymxjmnb9b
                          | igbfek2f8xd5vcozwc6mvu
                          | kqoce2mai7legb67b3_l3ofi1v
                          | mqxidx634c8oo3gea0__8s
                          | vr63zqx6y0ffx32ubvl670vs9m6qf
                          | wydnyq82nhj8gfglsmtj8ffh
                          ;
  

  assign v0qy_p3s0bq9bqj0mz = ({l4e4x5iuocpq14dam9ucku{fi5j2nq20y39ylylwhs      }} & u99tnldu986760c5      )
                          | ({l4e4x5iuocpq14dam9ucku{vikfdhomdfhf7ewfaitsy_gj    }} & nhzryulpguznnnqmzgn0    )
                          | ({l4e4x5iuocpq14dam9ucku{fpsdt9vdjcwssz9tezden07r7}} & jlnkd6qhsmjqw47tf1t64byci)
                          | ({l4e4x5iuocpq14dam9ucku{b7z98rnx88w42eg6952nx8x     }} & s67r7tvcckkpgs9     )
                          | ({l4e4x5iuocpq14dam9ucku{nme7un7hr7uwq6h4qmctk_srkw   }} & x4lgrwp6fc79b0ehv9   )
                          | ({l4e4x5iuocpq14dam9ucku{d3o9i8v1m3g16rvwhai2wh7   }} & dbw_jljmitz3e_zmp   )
                          | ({l4e4x5iuocpq14dam9ucku{qhcnhctsg82wxcyhu80cuex4c }} & u9fc6nt5deod0x3wvfv )
                          | ({l4e4x5iuocpq14dam9ucku{oadttvx13julmicav817mtk5jev  }} & v0gpnd2kvonwrxb2d1  )
                          ;

 
  wire o32vpum2sraiyu3dl       = (v0qy_p3s0bq9bqj0mz == klcv32s524noj675s      ) & e8ay6vzax1puil9e;
  wire xf53wre_7y6eulqc3z1     = (v0qy_p3s0bq9bqj0mz == qi8j2njkyk3a22m95kc8jquq    ) & e8ay6vzax1puil9e;
  wire tg7zajgb1p_43zyczn8ui0jqwt1 = (v0qy_p3s0bq9bqj0mz == ai81jjukhk7_uoovfndq690s) & e8ay6vzax1puil9e;
  wire ukeqsfnih_s1o_0dk_w8els      = (v0qy_p3s0bq9bqj0mz == x2yiem7xqi4jww3op6siel     ) & e8ay6vzax1puil9e;
  wire x2kluxpzwo7e4bojx6w9ph3    = (v0qy_p3s0bq9bqj0mz == r_h500kxshad5gkq4zgdswta   ) & e8ay6vzax1puil9e;
  wire ab9up1x30lvk2h8t3f89ads    = (v0qy_p3s0bq9bqj0mz == qka__s7my8mvb4j5dhd071   ) & e8ay6vzax1puil9e;
  wire mw35p42od2rj_je2r6w0fdsh  = (v0qy_p3s0bq9bqj0mz == iosvpnl0hccumt4jze71nkq0d ) & e8ay6vzax1puil9e;
  wire mvdyagaaq6p17_49ubja_i   = (v0qy_p3s0bq9bqj0mz == ghxu50th5tej1yhl8zrb7lticj  ) & e8ay6vzax1puil9e;
  
  assign d4ab_e8ynn1a53_52a3 = (v0qy_p3s0bq9bqj0mz != klcv32s524noj675s | q5xw1oq2dyd3_r9 != klcv32s524noj675s | t523n0nf23b9vzzq);
  
  wire qzvusaw9lyc30cqsig7tl18w = ab9up1x30lvk2h8t3f89ads | mw35p42od2rj_je2r6w0fdsh | mvdyagaaq6p17_49ubja_i;

  wire ra07vicltr81_z8;
  wire g_7nc4dw6abcm;
  wire wi0fxe4_7r_vmld14fes8;
  wire n56r23zad9uraj_56o5;
  wire cmbd5g6aephposs;

  wire vcrfj57jgo3_pfo6v7kc;
  wire eolarjcu8sj7ukw3z221 = qzvusaw9lyc30cqsig7tl18w;
  wire lr4kbcbmh553jxuqn1x6f7v = o32vpum2sraiyu3dl;
  wire cf0hcezcjw6tj35omcawkeu9k = eolarjcu8sj7ukw3z221 | ~lr4kbcbmh553jxuqn1x6f7v;
  wire mzv88i8pr6n26vqf5_twzv = eolarjcu8sj7ukw3z221 |  lr4kbcbmh553jxuqn1x6f7v;
  ux607_gnrl_dfflr #(1) eamdwvn9urivtulg38uhp11be (mzv88i8pr6n26vqf5_twzv, cf0hcezcjw6tj35omcawkeu9k, vcrfj57jgo3_pfo6v7kc, gf33atgy, ru_wi);
 
 
  wire fd08zi5rybh6vf54gwko2;
  wire vq31_o6tysljm1xafo_ = xf53wre_7y6eulqc3z1 & wi0fxe4_7r_vmld14fes8;
  wire b5etb0sfypx9bqbcl7j85 = o32vpum2sraiyu3dl | qzvusaw9lyc30cqsig7tl18w | (xf53wre_7y6eulqc3z1 & n56r23zad9uraj_56o5)
                             | (b0l_kaqp & fd08zi5rybh6vf54gwko2);
  wire uk1424xmyv6x032rcgt83o5 = vq31_o6tysljm1xafo_ | ~b5etb0sfypx9bqbcl7j85;
  wire mqwqhnwxw0yfg3kjgux62fe = vq31_o6tysljm1xafo_ |  b5etb0sfypx9bqbcl7j85;
  ux607_gnrl_dfflr #(1) bf50_oine070crftx_4e9fpn (mqwqhnwxw0yfg3kjgux62fe, uk1424xmyv6x032rcgt83o5, fd08zi5rybh6vf54gwko2, gf33atgy, ru_wi);
  assign m0rgjbiqu6nadc33k5   = fd08zi5rybh6vf54gwko2;


  wire g2s1v1ri9nldpeph;
  wire dw0p79b1rf939hlll6 = b0l_kaqp & (fd08zi5rybh6vf54gwko2 | wi0fxe4_7r_vmld14fes8);
  wire ri446c3ih_jjkv1p = g2s1v1ri9nldpeph & (pffig1fl4xtnw | j48quvipiuwft);
  wire o63476a_nj59fir4 = dw0p79b1rf939hlll6 | ~ri446c3ih_jjkv1p;
  wire ms_ak_pb6xlzqw0ytp0sc = dw0p79b1rf939hlll6 |  ri446c3ih_jjkv1p;
  ux607_gnrl_dfflr #(1) uo6kz7awhf3ohpw8_ukg24 (ms_ak_pb6xlzqw0ytp0sc, o63476a_nj59fir4, g2s1v1ri9nldpeph, gf33atgy, ru_wi);
  assign xhehq_1td3fs   = g2s1v1ri9nldpeph;

  wire ryl6cvoaujvg6lri3e;
  wire e4o3z9p2mcnv45_8689dc = xf53wre_7y6eulqc3z1 & n56r23zad9uraj_56o5;
  wire s_k9i3yr4co1idhz3uw = o32vpum2sraiyu3dl | qzvusaw9lyc30cqsig7tl18w | (xf53wre_7y6eulqc3z1 & wi0fxe4_7r_vmld14fes8) 
                             | (b0l_kaqp & ryl6cvoaujvg6lri3e);
  wire p32tne7wbmf1a2xfedzn = e4o3z9p2mcnv45_8689dc | ~s_k9i3yr4co1idhz3uw;
  wire iqmu4_hmnmtd7akp_eepcw = e4o3z9p2mcnv45_8689dc |  s_k9i3yr4co1idhz3uw;
  ux607_gnrl_dfflr #(1) wyugazwhhsieip9h6abkor4e (iqmu4_hmnmtd7akp_eepcw, p32tne7wbmf1a2xfedzn, ryl6cvoaujvg6lri3e, gf33atgy, ru_wi);


  wire o6zs2age2tfbqxrs;
  wire vjma_e6hodrjml2oc7v3_ = b0l_kaqp & (ryl6cvoaujvg6lri3e | n56r23zad9uraj_56o5);
  wire jpp3ptuoo5zgglpz = o6zs2age2tfbqxrs & (pffig1fl4xtnw | j48quvipiuwft);
  wire mrhxkk_wy5dvgma22yeu = vjma_e6hodrjml2oc7v3_ | ~jpp3ptuoo5zgglpz;
  wire q_1y742wiob55eeirm16 = vjma_e6hodrjml2oc7v3_ |  jpp3ptuoo5zgglpz;
  ux607_gnrl_dfflr #(1) rshg27mrrbhe7iibfb7sk (q_1y742wiob55eeirm16, mrhxkk_wy5dvgma22yeu, o6zs2age2tfbqxrs, gf33atgy, ru_wi);


  wire j1bzjadadk5nl_fo89slx = ~vcrfj57jgo3_pfo6v7kc;
  assign ra07vicltr81_z8 = m01i4z2a2meu & j1bzjadadk5nl_fo89slx;
  
  wire wirum77y73a0kflzedlta7wsj2u = ~fd08zi5rybh6vf54gwko2 & ~g2s1v1ri9nldpeph & ~g_7nc4dw6abcm  
                                & ~ryl6cvoaujvg6lri3e; 
  assign wi0fxe4_7r_vmld14fes8 = kbi8qdl8tmgm5j0uu1p1xu0 & wirum77y73a0kflzedlta7wsj2u; 
  
  wire dt99g_aav1hs6emyjgs860 = ~ra07vicltr81_z8;
  assign g_7nc4dw6abcm = rxosbn3wj_1o6y20fv & dt99g_aav1hs6emyjgs860;

  wire uf7r7106uyloyo2m5b0gax9tds2 = ~ra07vicltr81_z8 & ~wi0fxe4_7r_vmld14fes8 & ~g_7nc4dw6abcm & ~ryl6cvoaujvg6lri3e & ~o6zs2age2tfbqxrs 
                                & ~fd08zi5rybh6vf54gwko2; 
  assign n56r23zad9uraj_56o5 = ntychvakx3t8mzzgh8_ev & uf7r7106uyloyo2m5b0gax9tds2;
  
  assign cmbd5g6aephposs = wi0fxe4_7r_vmld14fes8 | n56r23zad9uraj_56o5;


  
  
  
  

  wire ufyt0wbivcs5bjbl;  
  wire po6_33ky73vq870 = ra07vicltr81_z8 & ~mou2g2qz02878jxn & ~yyz7lhabpe7x17h10y; 
  wire sosk9cm52vulowzu3l = g_7nc4dw6abcm & pffig1fl4xtnw; 
  wire b_l7znzwzqo4w4x = po6_33ky73vq870 | ~sosk9cm52vulowzu3l;
  wire hk396ql949nz_eh = po6_33ky73vq870 | sosk9cm52vulowzu3l;
  ux607_gnrl_dfflrs #(1) yhu5possa265omubk (hk396ql949nz_eh, b_l7znzwzqo4w4x, ufyt0wbivcs5bjbl, gf33atgy, ru_wi);
  wire [1:0] ygrnmd7zc14ooux0; 
  wire [1:0] lz9tkah9a8uzawtmhpo8za;
  wire lp6ujhfxz8naf8fdovc;
  ux607_gnrl_dfflrs #(1) ns6ajy6cakaho1y4pvjryop (lp6ujhfxz8naf8fdovc, lz9tkah9a8uzawtmhpo8za[0], ygrnmd7zc14ooux0[0], gf33atgy, ru_wi);
  ux607_gnrl_dfflr #(1) txa7gwkrtk7l4yq9ez1dl1i01 (lp6ujhfxz8naf8fdovc, lz9tkah9a8uzawtmhpo8za[1], ygrnmd7zc14ooux0[1], gf33atgy, ru_wi);


  wire [l4e4x5iuocpq14dam9ucku-1:0] jrfy34s3g08z1b27 = mou2g2qz02878jxn      ? qka__s7my8mvb4j5dhd071  :  
                                                   yyz7lhabpe7x17h10y    ? iosvpnl0hccumt4jze71nkq0d:
                                                                          ghxu50th5tej1yhl8zrb7lticj ;

  
  
  assign wfoen161d4r42bkqp34lj = fi5j2nq20y39ylylwhs & (ra07vicltr81_z8 | wi0fxe4_7r_vmld14fes8 | n56r23zad9uraj_56o5 | g_7nc4dw6abcm | x3h2m98yhzqwpra5q0q);
  assign u99tnldu986760c5 = x3h2m98yhzqwpra5q0q             ? ghxu50th5tej1yhl8zrb7lticj:
                          ra07vicltr81_z8                    ? jrfy34s3g08z1b27     :
                          g_7nc4dw6abcm                   ? klcv32s524noj675s    :  
                          cmbd5g6aephposs & ~ufyt0wbivcs5bjbl ? qi8j2njkyk3a22m95kc8jquq  : 
                                                          klcv32s524noj675s    ;
  
  

  wire xk9onv5o60eyf9;
  wire udxk4gyp4kyi;
  wire e7x7c02tu7umslg729;


  
  assign dqc3ngr_5saws_sp75dkhv = vikfdhomdfhf7ewfaitsy_gj & (ra07vicltr81_z8 |  e7x7c02tu7umslg729 |xk9onv5o60eyf9 | udxk4gyp4kyi | g_7nc4dw6abcm);
  assign nhzryulpguznnnqmzgn0 = ra07vicltr81_z8                                       ? jrfy34s3g08z1b27       :
                            e7x7c02tu7umslg729                                   ? x2yiem7xqi4jww3op6siel     :
                            xk9onv5o60eyf9                                       ? ai81jjukhk7_uoovfndq690s:
                            udxk4gyp4kyi & g_7nc4dw6abcm                        ? klcv32s524noj675s   : 
                            udxk4gyp4kyi & (g2s1v1ri9nldpeph | o6zs2age2tfbqxrs)  ? r_h500kxshad5gkq4zgdswta   : 
                            udxk4gyp4kyi    ? klcv32s524noj675s      : 
                                             qi8j2njkyk3a22m95kc8jquq    ;


  
  assign wd2v3s292zarv6r_qtszoymxjmnb9b = fpsdt9vdjcwssz9tezden07r7;
  assign jlnkd6qhsmjqw47tf1t64byci = ra07vicltr81_z8                               ? jrfy34s3g08z1b27   :
                                g_7nc4dw6abcm                              ? qi8j2njkyk3a22m95kc8jquq: 
                                cmbd5g6aephposs                           ? qi8j2njkyk3a22m95kc8jquq:
                                                                           klcv32s524noj675s  ;

  
  assign igbfek2f8xd5vcozwc6mvu = b7z98rnx88w42eg6952nx8x;
  assign s67r7tvcckkpgs9 = ra07vicltr81_z8                               ? jrfy34s3g08z1b27   :
                           g_7nc4dw6abcm                              ? qi8j2njkyk3a22m95kc8jquq: 
                           cmbd5g6aephposs                           ? qi8j2njkyk3a22m95kc8jquq:
                                                                      klcv32s524noj675s  ;


  
  assign kqoce2mai7legb67b3_l3ofi1v = nme7un7hr7uwq6h4qmctk_srkw;
  assign x4lgrwp6fc79b0ehv9 = ra07vicltr81_z8                                 ? jrfy34s3g08z1b27   :
                             b3ymasxx4cnt | pffig1fl4xtnw | j48quvipiuwft ? qi8j2njkyk3a22m95kc8jquq : 
                                                                          r_h500kxshad5gkq4zgdswta;


  wire c5rsvjgxx0datlxovp6f;
  assign sd4rdwq_5i7fe5 = c5rsvjgxx0datlxovp6f & (d3o9i8v1m3g16rvwhai2wh7 | qhcnhctsg82wxcyhu80cuex4c | oadttvx13julmicav817mtk5jev);
  assign ew6x7412r46 = sd4rdwq_5i7fe5;
  
  assign mqxidx634c8oo3gea0__8s = d3o9i8v1m3g16rvwhai2wh7 & sd4rdwq_5i7fe5;
  assign dbw_jljmitz3e_zmp = klcv32s524noj675s;

  
  assign vr63zqx6y0ffx32ubvl670vs9m6qf = qhcnhctsg82wxcyhu80cuex4c & sd4rdwq_5i7fe5;
  assign u9fc6nt5deod0x3wvfv = klcv32s524noj675s;

  
  assign wydnyq82nhj8gfglsmtj8ffh = oadttvx13julmicav817mtk5jev & sd4rdwq_5i7fe5;
  assign v0gpnd2kvonwrxb2d1 = klcv32s524noj675s;

  





  
  localparam lvcpofkw_r     = 5;
  localparam ag6ywem9ln_z    = 5;
  localparam r3kzsezay2f8jnn  = ~ 32'b0;
  localparam e306hu2yanbe   = {1'b0,{6{1'b1}}};
  
  wire [7-1:0] hfi2y7aons_t      = lvcpofkw_r[7-1:0];
  wire [7-1:0] l_jrtjcsdy5s_     = ag6ywem9ln_z[7-1:0];
  wire [7-1:0] nqjl3s3cfs_tpo   = r3kzsezay2f8jnn[7-1:0];
  wire [7-1:0] zykarimzgmuoq    = e306hu2yanbe[7-1:0];

  wire [7-1:0] fivfh22sha8ppz;
  wire [7-1:0] uyqega7f8ezigfj9m4m = (
                                                      c5rsvjgxx0datlxovp6f  
                                                      | (vikfdhomdfhf7ewfaitsy_gj & g_7nc4dw6abcm & (xk9onv5o60eyf9 | e7x7c02tu7umslg729)) 
                                                      | (fpsdt9vdjcwssz9tezden07r7 | b7z98rnx88w42eg6952nx8x) 
                                                     ) ? {7{1'b0}} : (fivfh22sha8ppz + {{7-1{1'b0}},1'b1});
  wire ygxy_nacztbq4h6kob5 = (fpsdt9vdjcwssz9tezden07r7 | b7z98rnx88w42eg6952nx8x) 
                        | (vikfdhomdfhf7ewfaitsy_gj & ~(g_7nc4dw6abcm & pffig1fl4xtnw))
                        | (vikfdhomdfhf7ewfaitsy_gj & udxk4gyp4kyi) 
                        | d3o9i8v1m3g16rvwhai2wh7 | qhcnhctsg82wxcyhu80cuex4c | oadttvx13julmicav817mtk5jev;
  ux607_gnrl_dfflr #(7) vpiaphyhutlsllwli0fbw (ygxy_nacztbq4h6kob5, uyqega7f8ezigfj9m4m, fivfh22sha8ppz, gf33atgy, ru_wi);

  wire [7-1:0] toomwmpbxsmlbhqtx0oi8y4pw =  vikfdhomdfhf7ewfaitsy_gj    ? hfi2y7aons_t    :
                                                            d3o9i8v1m3g16rvwhai2wh7   ? l_jrtjcsdy5s_   :
                                                            qhcnhctsg82wxcyhu80cuex4c ? nqjl3s3cfs_tpo :
                                                            oadttvx13julmicav817mtk5jev  ? zykarimzgmuoq  :
                                                                                      {7{1'b0}};

  assign c5rsvjgxx0datlxovp6f = (fivfh22sha8ppz == toomwmpbxsmlbhqtx0oi8y4pw);
  

  
  
  
  
  
  
  wire hj0v28frzjss37;
  wire e2vq9uu_okytxq;
  wire [1:0] zkrae_ghfjkro2af = ygrnmd7zc14ooux0;

  wire [1:0] hajgx9_kx9125g = ({2{ygrnmd7zc14ooux0 == 2'b00}} & 2'b01)
                           | ({2{ygrnmd7zc14ooux0 == 2'b01}} & 2'b00)
                           | ({2{ygrnmd7zc14ooux0 == 2'b10}} & 2'b00)
                           ;

  wire [1:0] rdu0huute6u3tv4u = ({2{ygrnmd7zc14ooux0 == 2'b00}} & 2'b10)
                           | ({2{ygrnmd7zc14ooux0 == 2'b01}} & 2'b10)
                           | ({2{ygrnmd7zc14ooux0 == 2'b10}} & 2'b01)
                           ;

  wire [1:0] crdbk04fibhyphv = ({2{fivfh22sha8ppz[2:1] == 2'b00}} & zkrae_ghfjkro2af)
                         | ({2{fivfh22sha8ppz[2:1] == 2'b01}} & hajgx9_kx9125g)
                         | ({2{fivfh22sha8ppz[2:1] == 2'b10}} & rdu0huute6u3tv4u)
                         ;
 
  wire [27-1:0] uiigu5mk12 = (vcrfj57jgo3_pfo6v7kc | fd08zi5rybh6vf54gwko2) ? k11nc9vg2x3_cg_semdn : y0__7wpxqx83r42pl;

  wire [6-1:0] r3ud3glj937o4_ = ({6{crdbk04fibhyphv == 2'b00}} & uiigu5mk12[6-1:0    ])
                                                | ({6{crdbk04fibhyphv == 2'b01}} & uiigu5mk12[6-1+9:9  ]) 
                                                | ({6{crdbk04fibhyphv == 2'b10}} & uiigu5mk12[6-1+18:18]) 
                                                ;
  

  wire ec9ae2r_4n0dqq8xd73im = ~fivfh22sha8ppz[0]; 
  wire warib_3d5o1png93gezjz2 = ~fivfh22sha8ppz[0];
  wire ruuziixs92g5sudfr9ki = 1'b0;
  wire x197sqagslv9avl082ww = 1'b0;
  wire [66-1:0] ztixdkyplyl9m0b51_c0qha = {66{1'b0}};
  wire [66-1:0] ythnrofnodk8gj5gm0owzh = {66{1'b0}};
  wire [6-1:0] qj0rupp44fw6_cqrup1 = r3ud3glj937o4_;
  wire [66-1:0] hombiq_bhjjgnsmqu6k1bh = qbksws8auoc48qp3sb;
  wire [66-1:0] q6w031s_tfpr__jvavyl4wez6 = xyeddoohku7q6ja9pvnp;

  wire wamg6_ub3yboo4       = hombiq_bhjjgnsmqu6k1bh[0:0];
  wire w8jc05jmo7k4cu1csud  = hombiq_bhjjgnsmqu6k1bh[1:1];
  wire dvgtpjau3srjx68f8q    = hombiq_bhjjgnsmqu6k1bh[2:2];
  wire ordss3f1jraq8uh3x    = hombiq_bhjjgnsmqu6k1bh[3:3];
  wire k3s02jf92kope8b90       = hombiq_bhjjgnsmqu6k1bh[4:4];
  wire uke__x98g6o37        = hombiq_bhjjgnsmqu6k1bh[5:5];
  wire t9mzd13l1ozfo7lkf      = hombiq_bhjjgnsmqu6k1bh[6:6];
  wire [1:0                       ] o_dq7s9iqfyodwne8411u = hombiq_bhjjgnsmqu6k1bh[8:7];
  wire [16-1:0      ] ha0z9pxiveln47mn4m      = hombiq_bhjjgnsmqu6k1bh[24:9];
  wire [20-1:0        ] k_w1g2qu45yvxf       = hombiq_bhjjgnsmqu6k1bh[44:25];
  wire [21-1:0] btt1j9ogtns        = hombiq_bhjjgnsmqu6k1bh[65:45];


  wire t9gdufsox031zlci6d       = q6w031s_tfpr__jvavyl4wez6[0:0];
  wire egcy0ygmvlb_3ul1z7ttso  = q6w031s_tfpr__jvavyl4wez6[1:1];
  wire nq34u_g0r21b_d3th    = q6w031s_tfpr__jvavyl4wez6[2:2];
  wire ajmz0zyeikdq59ltt_7    = q6w031s_tfpr__jvavyl4wez6[3:3];
  wire l8qaaplst40ukqs_h       = q6w031s_tfpr__jvavyl4wez6[4:4];
  wire r3w0ndgscxl6i2fj        = q6w031s_tfpr__jvavyl4wez6[5:5];
  wire b3jr6fc2nimoowyktn5      = q6w031s_tfpr__jvavyl4wez6[6:6];
  wire [1:0                       ] j5yuuochvphc58tzu29i = q6w031s_tfpr__jvavyl4wez6[8:7];
  wire [16-1:0      ] qgfk9ulbi6ib7sp      = q6w031s_tfpr__jvavyl4wez6[24:9];
  wire [20-1:0        ] dvp8fjkox7t_y2       = q6w031s_tfpr__jvavyl4wez6[44:25];
  wire [21-1:0] lh0ro02ju2ra8vh        = q6w031s_tfpr__jvavyl4wez6[65:45];

  wire [21-1:0] lftuqy9et97rb30lh9 = ({21{crdbk04fibhyphv == 2'b00}} & {21{1'b1}})
                                                    | ({21{crdbk04fibhyphv == 2'b01}} & {{21-9 {1'b1}},  9'b0})
                                                    | ({21{crdbk04fibhyphv == 2'b10}} & {{21-18{1'b1}}, 18'b0})
                                                    ;

  wire [21-1:0] nj8advwe4r3iefjlp = uiigu5mk12[27-1:6] & lftuqy9et97rb30lh9;


  wire or2jrhp2d5b1798bveca = (nj8advwe4r3iefjlp == btt1j9ogtns);
  wire llqi__ojtcawwmml0 = (nj8advwe4r3iefjlp == lh0ro02ju2ra8vh);
  wire q9a976q8fdpkb_cuyx18gr57 = (crdbk04fibhyphv == o_dq7s9iqfyodwne8411u);
  wire q9xr0vqthnop3ifjrvfwyvbvcs4vv = (crdbk04fibhyphv == j5yuuochvphc58tzu29i);

  wire uzgdmfu0z6qg2vr_d363mx0v3z16vc = (j3d84gxpt2b4pd8 == ha0z9pxiveln47mn4m) & ~t9mzd13l1ozfo7lkf; 
  wire xmusnbfgqnhl529_izdr6u5tv7ky = (j3d84gxpt2b4pd8 == qgfk9ulbi6ib7sp) & ~b3jr6fc2nimoowyktn5;

  wire sabys6s2q2y_ecnfqfw9 = (hnc10arn_rd == ha0z9pxiveln47mn4m);
  wire ck4rswltzjdgr0bs9op4hm = (hnc10arn_rd == qgfk9ulbi6ib7sp);
 
 
  wire cgewm1crv6gxm6h7r = wamg6_ub3yboo4 & or2jrhp2d5b1798bveca & q9a976q8fdpkb_cuyx18gr57 & (sabys6s2q2y_ecnfqfw9 | t9mzd13l1ozfo7lkf);
  wire iwxf98mwbvgvf3dd4u5 = t9gdufsox031zlci6d & llqi__ojtcawwmml0 & q9xr0vqthnop3ifjrvfwyvbvcs4vv & (ck4rswltzjdgr0bs9op4hm | b3jr6fc2nimoowyktn5);
  wire jii9roub28fcas     = (cgewm1crv6gxm6h7r | iwxf98mwbvgvf3dd4u5) & fivfh22sha8ppz[0] & vikfdhomdfhf7ewfaitsy_gj & e2vq9uu_okytxq; 
  
  assign xk9onv5o60eyf9 = jii9roub28fcas & ~e7x7c02tu7umslg729;
  assign udxk4gyp4kyi = c5rsvjgxx0datlxovp6f & ~xk9onv5o60eyf9;
 
  wire p90_43ok_ek4ch69      = 1'b1; 
  wire en1yucx5gpxpk_dgbhz = cgewm1crv6gxm6h7r ? w8jc05jmo7k4cu1csud : egcy0ygmvlb_3ul1z7ttso;
  wire gn5qnj2atfazc8hhq   = cgewm1crv6gxm6h7r ? dvgtpjau3srjx68f8q : nq34u_g0r21b_d3th;
  wire g6ra3jt_jkiw58fxov   = cgewm1crv6gxm6h7r ? ordss3f1jraq8uh3x : ajmz0zyeikdq59ltt_7;
  wire wmsb_vgasb6751vio      = cgewm1crv6gxm6h7r ? k3s02jf92kope8b90 : l8qaaplst40ukqs_h;
  wire hyrmhupqn6h7       = cgewm1crv6gxm6h7r ? uke__x98g6o37 : r3w0ndgscxl6i2fj;
  wire j0u4fh_zs2avw5dd     = cgewm1crv6gxm6h7r ? t9mzd13l1ozfo7lkf : b3jr6fc2nimoowyktn5;
  wire [1:0                       ] wqigu3jp6nr52maoxma = cgewm1crv6gxm6h7r ? o_dq7s9iqfyodwne8411u : j5yuuochvphc58tzu29i;
  wire [16-1:0      ] c7felg6fri354v      = cgewm1crv6gxm6h7r ? ha0z9pxiveln47mn4m : qgfk9ulbi6ib7sp;
  wire [20-1:0        ] eulvtosq2vlauykz       = cgewm1crv6gxm6h7r ? k_w1g2qu45yvxf : dvp8fjkox7t_y2;
  wire [21-1:0] uwhuvcsr1ocz        = cgewm1crv6gxm6h7r ? btt1j9ogtns : lh0ro02ju2ra8vh;
  
  wire [66-1:0] wsjju32txk0_f4u51cf = {
                                                       uwhuvcsr1ocz,
                                                       eulvtosq2vlauykz,
                                                       c7felg6fri354v,
                                                       wqigu3jp6nr52maoxma,
                                                       j0u4fh_zs2avw5dd,
                                                       hyrmhupqn6h7,
                                                       wmsb_vgasb6751vio,
                                                       g6ra3jt_jkiw58fxov,
                                                       gn5qnj2atfazc8hhq,
                                                       en1yucx5gpxpk_dgbhz,
                                                       p90_43ok_ek4ch69
                                                     };

  wire [66-1:0] vy1fm7h4jitsqpc669;
  wire fdj_rumy116244c8e = xk9onv5o60eyf9 & vikfdhomdfhf7ewfaitsy_gj;
  ux607_gnrl_dfflr #(66) bo28lkq0pvimbwqy568z (fdj_rumy116244c8e, wsjju32txk0_f4u51cf, vy1fm7h4jitsqpc669, gf33atgy, ru_wi);

  
  wire c7sq9i2s8;
  wire qux9r2p2iev = iwxf98mwbvgvf3dd4u5;
  wire xqi3gtxuh3hu3lg0 = xk9onv5o60eyf9 & vikfdhomdfhf7ewfaitsy_gj;
  ux607_gnrl_dfflr #(1) iuh1ieh4oqb0py_ (xqi3gtxuh3hu3lg0, qux9r2p2iev, c7sq9i2s8, gf33atgy, ru_wi);

  assign lp6ujhfxz8naf8fdovc = xk9onv5o60eyf9;
  assign lz9tkah9a8uzawtmhpo8za = wqigu3jp6nr52maoxma;
  
  
  wire [1:0] dewq6i6jchg2nhnxp = (rm1dxjejhq7dh3q5m & fd08zi5rybh6vf54gwko2) ? st2zalpx0uf : toox2fc0snvsr_n;


  
  wire ngvtudt6cbj1f2jivms_2v68xzv = jii9roub28fcas & fd08zi5rybh6vf54gwko2 & ~on37whxvtxni09my52drx & ~wmsb_vgasb6751vio;

  
  wire g05s70mnpo5aoa7bm_mzna7q = jii9roub28fcas & fd08zi5rybh6vf54gwko2 & ~on37whxvtxni09my52drx & ~gn5qnj2atfazc8hhq;

  
  wire qug5b6ehslx92r_4ko8qojhvi = jii9roub28fcas & fd08zi5rybh6vf54gwko2 &  on37whxvtxni09my52drx & ~g6ra3jt_jkiw58fxov & (~ni01kj42oob2x | (~en1yucx5gpxpk_dgbhz & ni01kj42oob2x));

  
  wire y5e42uisfvamoofa5wwv5hx4_477f = jii9roub28fcas & ryl6cvoaujvg6lri3e & ~en1yucx5gpxpk_dgbhz;
  
  
  wire yp7t_qd1qr9zw91ucj04s1c4 = jii9roub28fcas & (dewq6i6jchg2nhnxp == 2'b00) & ~hyrmhupqn6h7;

  
  wire br7hk4brb090w93_9hki68oz = jii9roub28fcas & (dewq6i6jchg2nhnxp == 2'b01) &  hyrmhupqn6h7 & (ryl6cvoaujvg6lri3e | fd08zi5rybh6vf54gwko2 & ~ah8kjlmvnaxzbi);

  assign e7x7c02tu7umslg729 = 1'b0
                        | ngvtudt6cbj1f2jivms_2v68xzv 
                        | g05s70mnpo5aoa7bm_mzna7q
                        | qug5b6ehslx92r_4ko8qojhvi
                        | y5e42uisfvamoofa5wwv5hx4_477f
                        | yp7t_qd1qr9zw91ucj04s1c4
                        | br7hk4brb090w93_9hki68oz
                        ;

  wire einnn_ogj8zi41_ymq0;
  wire vk16l9d1hagkpnu1m6b8r3xibw = vikfdhomdfhf7ewfaitsy_gj & fivfh22sha8ppz[0] & e7x7c02tu7umslg729 & e2vq9uu_okytxq;
  wire xr1l8cxhibtemkqzsugctw_ = ~vikfdhomdfhf7ewfaitsy_gj;
  wire qrv46o8vrmhbgum5iqhox = vk16l9d1hagkpnu1m6b8r3xibw | ~xr1l8cxhibtemkqzsugctw_;
  wire oklb8iebvitzjs0a8pjx6qej7 = vk16l9d1hagkpnu1m6b8r3xibw |  xr1l8cxhibtemkqzsugctw_;
  ux607_gnrl_dfflr #(1) nuw6pc54vneju1yvueua3vhacuej (oklb8iebvitzjs0a8pjx6qej7, qrv46o8vrmhbgum5iqhox, einnn_ogj8zi41_ymq0, gf33atgy, ru_wi);


  
  
  
  
  
  
  wire z3g4qkmuiyg_xfbwf7a2r = fd08zi5rybh6vf54gwko2;
  wire be_urjfihso_vqebnp9heqpi = ryl6cvoaujvg6lri3e;
  wire [55-1:0] lmvxjn5zlc78w16q73_ybu47 = {55{1'b0}};
  wire [51-1:0] h2zqfgvjbnma19r37rn9s = {51{1'b0}};
  wire zz2s0dg_zi49zvpaj8tygzbbpi = 1'b0;
  wire ba9aqillrmgw1eh2as1fhaja02rx6 = 1'b0;

  wire m7oe8scer3o7hu_v3ct5xtbe = einnn_ogj8zi41_ymq0;
  wire vudlml4_g7imvjcp1o18uo = 1'b0;

  
  
  
  
  

  wire t5n0cdht9qz0      = 1'b1; 
  wire q6chl10rx0r6sbnek_ = vy1fm7h4jitsqpc669[1:1];
  wire ior8m0p_l8iwxlwqk   = vy1fm7h4jitsqpc669[2:2];
  wire xglu0pzbtmtkekf   = vy1fm7h4jitsqpc669[3:3];
  wire gupypwowvqcf6b      = vy1fm7h4jitsqpc669[4:4];
  wire nn4zx06ycyciewu       = vy1fm7h4jitsqpc669[5:5];
  
  wire [1:0                 ] syjrm2mxj5tb9bhyqkx12 = vy1fm7h4jitsqpc669[8:7];
  
  wire [20-1:0  ] evv374je2a154hj       = vy1fm7h4jitsqpc669[44:25];
  
  
  wire [27-1:0] r23l7tyg0dluw3tzwox = ({27{syjrm2mxj5tb9bhyqkx12 == 2'b00}} & {27{1'b1}}) 
                                                | ({27{syjrm2mxj5tb9bhyqkx12 == 2'b01}} & {{27-9{1'b1}}  , 9'b0})
                                                | ({27{syjrm2mxj5tb9bhyqkx12 == 2'b10}} & {{27-18{1'b1}} , 18'b0});
  wire [27-1:0] lce7w9vhg8u      = uiigu5mk12 & r23l7tyg0dluw3tzwox;

  wire yw6x0r1j6uhow9nf5qu1 = fd08zi5rybh6vf54gwko2;
  wire je1s58zp9x4crpu7sd0_c_md2 = ryl6cvoaujvg6lri3e;
  wire [55-1:0] lj_9z8lqgvo5bet98sorzh = {
                                                           lce7w9vhg8u,
                                                           evv374je2a154hj,
                                                           syjrm2mxj5tb9bhyqkx12,
                                                           nn4zx06ycyciewu,
                                                           gupypwowvqcf6b,
                                                           xglu0pzbtmtkekf,
                                                           ior8m0p_l8iwxlwqk,
                                                           q6chl10rx0r6sbnek_,
                                                           t5n0cdht9qz0
                                                          };

  wire [51-1:0] gr7kjbwg55_sgsv87k0z = {
                                                           lce7w9vhg8u,
                                                           evv374je2a154hj,
                                                           syjrm2mxj5tb9bhyqkx12,
                                                           nn4zx06ycyciewu,
                                                           t5n0cdht9qz0
                                                          };
  wire mhu5ty6fyi1g5i40jtfpgkenhfn = fd08zi5rybh6vf54gwko2;
  wire d35npx0cpwxc6siaubaf_mx76i3nbqk = ryl6cvoaujvg6lri3e;

  wire vbb4gb1qjbfm7yzd98_7t26 = 1'b0;
  wire rq1ykv7_2goh27c1eo3u3jyynj62 = 1'b0;

  
  
  
  
  
  
  
  wire [27-1:0] a896qcozpsi1ek5tm9;
  assign b0l_kaqp = ((fi5j2nq20y39ylylwhs & cmbd5g6aephposs & ufyt0wbivcs5bjbl)  
                    | (vikfdhomdfhf7ewfaitsy_gj & udxk4gyp4kyi)) 
                   & (b3ymasxx4cnt | pffig1fl4xtnw | j48quvipiuwft);  
  assign uhegwov_bgw = g2s1v1ri9nldpeph ?  k11nc9vg2x3_cg_semdn : y0__7wpxqx83r42pl;
  assign a896qcozpsi1ek5tm9 = g2s1v1ri9nldpeph ? k11nc9vg2x3_cg_semdn : y0__7wpxqx83r42pl;
  assign tlygxd1cs0w = (fd08zi5rybh6vf54gwko2 | wi0fxe4_7r_vmld14fes8) & on37whxvtxni09my52drx;
  assign i3o6jvv3t7i = (fd08zi5rybh6vf54gwko2 | wi0fxe4_7r_vmld14fes8) & ~on37whxvtxni09my52drx;
  assign xwd9yye9seo2l = o6zs2age2tfbqxrs;


  
  
  
  
  
  
  
  wire [6-1:0] g5cld0_xqbmy2o0oiio_4 = ({6{ermcr77dq4jhq99jq == 2'b00}} & a896qcozpsi1ek5tm9[6-1:0])
                                                        | ({6{ermcr77dq4jhq99jq == 2'b01}} & a896qcozpsi1ek5tm9[6+ 9-1: 9])
                                                        | ({6{ermcr77dq4jhq99jq == 2'b10}} & a896qcozpsi1ek5tm9[6+18-1:18])
                                                        ;
  wire sbd346v940_sel = (g5cld0_xqbmy2o0oiio_4 == 6'd0);
  wire hmtqrdaxj0_sel = (r3ud3glj937o4_ == 6'd0);
  wire sbd346v941_sel = (g5cld0_xqbmy2o0oiio_4 == 6'd1);
  wire hmtqrdaxj1_sel = (r3ud3glj937o4_ == 6'd1);
  wire sbd346v942_sel = (g5cld0_xqbmy2o0oiio_4 == 6'd2);
  wire hmtqrdaxj2_sel = (r3ud3glj937o4_ == 6'd2);
  wire sbd346v943_sel = (g5cld0_xqbmy2o0oiio_4 == 6'd3);
  wire hmtqrdaxj3_sel = (r3ud3glj937o4_ == 6'd3);
  wire sbd346v944_sel = (g5cld0_xqbmy2o0oiio_4 == 6'd4);
  wire hmtqrdaxj4_sel = (r3ud3glj937o4_ == 6'd4);
  wire sbd346v945_sel = (g5cld0_xqbmy2o0oiio_4 == 6'd5);
  wire hmtqrdaxj5_sel = (r3ud3glj937o4_ == 6'd5);
  wire sbd346v946_sel = (g5cld0_xqbmy2o0oiio_4 == 6'd6);
  wire hmtqrdaxj6_sel = (r3ud3glj937o4_ == 6'd6);
  wire sbd346v947_sel = (g5cld0_xqbmy2o0oiio_4 == 6'd7);
  wire hmtqrdaxj7_sel = (r3ud3glj937o4_ == 6'd7);
  wire sbd346v948_sel = (g5cld0_xqbmy2o0oiio_4 == 6'd8);
  wire hmtqrdaxj8_sel = (r3ud3glj937o4_ == 6'd8);
  wire sbd346v949_sel = (g5cld0_xqbmy2o0oiio_4 == 6'd9);
  wire hmtqrdaxj9_sel = (r3ud3glj937o4_ == 6'd9);
  wire sbd346v9410_sel = (g5cld0_xqbmy2o0oiio_4 == 6'd10);
  wire hmtqrdaxj10_sel = (r3ud3glj937o4_ == 6'd10);
  wire sbd346v9411_sel = (g5cld0_xqbmy2o0oiio_4 == 6'd11);
  wire hmtqrdaxj11_sel = (r3ud3glj937o4_ == 6'd11);
  wire sbd346v9412_sel = (g5cld0_xqbmy2o0oiio_4 == 6'd12);
  wire hmtqrdaxj12_sel = (r3ud3glj937o4_ == 6'd12);
  wire sbd346v9413_sel = (g5cld0_xqbmy2o0oiio_4 == 6'd13);
  wire hmtqrdaxj13_sel = (r3ud3glj937o4_ == 6'd13);
  wire sbd346v9414_sel = (g5cld0_xqbmy2o0oiio_4 == 6'd14);
  wire hmtqrdaxj14_sel = (r3ud3glj937o4_ == 6'd14);
  wire sbd346v9415_sel = (g5cld0_xqbmy2o0oiio_4 == 6'd15);
  wire hmtqrdaxj15_sel = (r3ud3glj937o4_ == 6'd15);
  wire sbd346v9416_sel = (g5cld0_xqbmy2o0oiio_4 == 6'd16);
  wire hmtqrdaxj16_sel = (r3ud3glj937o4_ == 6'd16);
  wire sbd346v9417_sel = (g5cld0_xqbmy2o0oiio_4 == 6'd17);
  wire hmtqrdaxj17_sel = (r3ud3glj937o4_ == 6'd17);
  wire sbd346v9418_sel = (g5cld0_xqbmy2o0oiio_4 == 6'd18);
  wire hmtqrdaxj18_sel = (r3ud3glj937o4_ == 6'd18);
  wire sbd346v9419_sel = (g5cld0_xqbmy2o0oiio_4 == 6'd19);
  wire hmtqrdaxj19_sel = (r3ud3glj937o4_ == 6'd19);
  wire sbd346v9420_sel = (g5cld0_xqbmy2o0oiio_4 == 6'd20);
  wire hmtqrdaxj20_sel = (r3ud3glj937o4_ == 6'd20);
  wire sbd346v9421_sel = (g5cld0_xqbmy2o0oiio_4 == 6'd21);
  wire hmtqrdaxj21_sel = (r3ud3glj937o4_ == 6'd21);
  wire sbd346v9422_sel = (g5cld0_xqbmy2o0oiio_4 == 6'd22);
  wire hmtqrdaxj22_sel = (r3ud3glj937o4_ == 6'd22);
  wire sbd346v9423_sel = (g5cld0_xqbmy2o0oiio_4 == 6'd23);
  wire hmtqrdaxj23_sel = (r3ud3glj937o4_ == 6'd23);
  wire sbd346v9424_sel = (g5cld0_xqbmy2o0oiio_4 == 6'd24);
  wire hmtqrdaxj24_sel = (r3ud3glj937o4_ == 6'd24);
  wire sbd346v9425_sel = (g5cld0_xqbmy2o0oiio_4 == 6'd25);
  wire hmtqrdaxj25_sel = (r3ud3glj937o4_ == 6'd25);
  wire sbd346v9426_sel = (g5cld0_xqbmy2o0oiio_4 == 6'd26);
  wire hmtqrdaxj26_sel = (r3ud3glj937o4_ == 6'd26);
  wire sbd346v9427_sel = (g5cld0_xqbmy2o0oiio_4 == 6'd27);
  wire hmtqrdaxj27_sel = (r3ud3glj937o4_ == 6'd27);
  wire sbd346v9428_sel = (g5cld0_xqbmy2o0oiio_4 == 6'd28);
  wire hmtqrdaxj28_sel = (r3ud3glj937o4_ == 6'd28);
  wire sbd346v9429_sel = (g5cld0_xqbmy2o0oiio_4 == 6'd29);
  wire hmtqrdaxj29_sel = (r3ud3glj937o4_ == 6'd29);
  wire sbd346v9430_sel = (g5cld0_xqbmy2o0oiio_4 == 6'd30);
  wire hmtqrdaxj30_sel = (r3ud3glj937o4_ == 6'd30);
  wire sbd346v9431_sel = (g5cld0_xqbmy2o0oiio_4 == 6'd31);
  wire hmtqrdaxj31_sel = (r3ud3glj937o4_ == 6'd31);
  wire sbd346v9432_sel = (g5cld0_xqbmy2o0oiio_4 == 6'd32);
  wire hmtqrdaxj32_sel = (r3ud3glj937o4_ == 6'd32);
  wire sbd346v9433_sel = (g5cld0_xqbmy2o0oiio_4 == 6'd33);
  wire hmtqrdaxj33_sel = (r3ud3glj937o4_ == 6'd33);
  wire sbd346v9434_sel = (g5cld0_xqbmy2o0oiio_4 == 6'd34);
  wire hmtqrdaxj34_sel = (r3ud3glj937o4_ == 6'd34);
  wire sbd346v9435_sel = (g5cld0_xqbmy2o0oiio_4 == 6'd35);
  wire hmtqrdaxj35_sel = (r3ud3glj937o4_ == 6'd35);
  wire sbd346v9436_sel = (g5cld0_xqbmy2o0oiio_4 == 6'd36);
  wire hmtqrdaxj36_sel = (r3ud3glj937o4_ == 6'd36);
  wire sbd346v9437_sel = (g5cld0_xqbmy2o0oiio_4 == 6'd37);
  wire hmtqrdaxj37_sel = (r3ud3glj937o4_ == 6'd37);
  wire sbd346v9438_sel = (g5cld0_xqbmy2o0oiio_4 == 6'd38);
  wire hmtqrdaxj38_sel = (r3ud3glj937o4_ == 6'd38);
  wire sbd346v9439_sel = (g5cld0_xqbmy2o0oiio_4 == 6'd39);
  wire hmtqrdaxj39_sel = (r3ud3glj937o4_ == 6'd39);
  wire sbd346v9440_sel = (g5cld0_xqbmy2o0oiio_4 == 6'd40);
  wire hmtqrdaxj40_sel = (r3ud3glj937o4_ == 6'd40);
  wire sbd346v9441_sel = (g5cld0_xqbmy2o0oiio_4 == 6'd41);
  wire hmtqrdaxj41_sel = (r3ud3glj937o4_ == 6'd41);
  wire sbd346v9442_sel = (g5cld0_xqbmy2o0oiio_4 == 6'd42);
  wire hmtqrdaxj42_sel = (r3ud3glj937o4_ == 6'd42);
  wire sbd346v9443_sel = (g5cld0_xqbmy2o0oiio_4 == 6'd43);
  wire hmtqrdaxj43_sel = (r3ud3glj937o4_ == 6'd43);
  wire sbd346v9444_sel = (g5cld0_xqbmy2o0oiio_4 == 6'd44);
  wire hmtqrdaxj44_sel = (r3ud3glj937o4_ == 6'd44);
  wire sbd346v9445_sel = (g5cld0_xqbmy2o0oiio_4 == 6'd45);
  wire hmtqrdaxj45_sel = (r3ud3glj937o4_ == 6'd45);
  wire sbd346v9446_sel = (g5cld0_xqbmy2o0oiio_4 == 6'd46);
  wire hmtqrdaxj46_sel = (r3ud3glj937o4_ == 6'd46);
  wire sbd346v9447_sel = (g5cld0_xqbmy2o0oiio_4 == 6'd47);
  wire hmtqrdaxj47_sel = (r3ud3glj937o4_ == 6'd47);
  wire sbd346v9448_sel = (g5cld0_xqbmy2o0oiio_4 == 6'd48);
  wire hmtqrdaxj48_sel = (r3ud3glj937o4_ == 6'd48);
  wire sbd346v9449_sel = (g5cld0_xqbmy2o0oiio_4 == 6'd49);
  wire hmtqrdaxj49_sel = (r3ud3glj937o4_ == 6'd49);
  wire sbd346v9450_sel = (g5cld0_xqbmy2o0oiio_4 == 6'd50);
  wire hmtqrdaxj50_sel = (r3ud3glj937o4_ == 6'd50);
  wire sbd346v9451_sel = (g5cld0_xqbmy2o0oiio_4 == 6'd51);
  wire hmtqrdaxj51_sel = (r3ud3glj937o4_ == 6'd51);
  wire sbd346v9452_sel = (g5cld0_xqbmy2o0oiio_4 == 6'd52);
  wire hmtqrdaxj52_sel = (r3ud3glj937o4_ == 6'd52);
  wire sbd346v9453_sel = (g5cld0_xqbmy2o0oiio_4 == 6'd53);
  wire hmtqrdaxj53_sel = (r3ud3glj937o4_ == 6'd53);
  wire sbd346v9454_sel = (g5cld0_xqbmy2o0oiio_4 == 6'd54);
  wire hmtqrdaxj54_sel = (r3ud3glj937o4_ == 6'd54);
  wire sbd346v9455_sel = (g5cld0_xqbmy2o0oiio_4 == 6'd55);
  wire hmtqrdaxj55_sel = (r3ud3glj937o4_ == 6'd55);
  wire sbd346v9456_sel = (g5cld0_xqbmy2o0oiio_4 == 6'd56);
  wire hmtqrdaxj56_sel = (r3ud3glj937o4_ == 6'd56);
  wire sbd346v9457_sel = (g5cld0_xqbmy2o0oiio_4 == 6'd57);
  wire hmtqrdaxj57_sel = (r3ud3glj937o4_ == 6'd57);
  wire sbd346v9458_sel = (g5cld0_xqbmy2o0oiio_4 == 6'd58);
  wire hmtqrdaxj58_sel = (r3ud3glj937o4_ == 6'd58);
  wire sbd346v9459_sel = (g5cld0_xqbmy2o0oiio_4 == 6'd59);
  wire hmtqrdaxj59_sel = (r3ud3glj937o4_ == 6'd59);
  wire sbd346v9460_sel = (g5cld0_xqbmy2o0oiio_4 == 6'd60);
  wire hmtqrdaxj60_sel = (r3ud3glj937o4_ == 6'd60);
  wire sbd346v9461_sel = (g5cld0_xqbmy2o0oiio_4 == 6'd61);
  wire hmtqrdaxj61_sel = (r3ud3glj937o4_ == 6'd61);
  wire sbd346v9462_sel = (g5cld0_xqbmy2o0oiio_4 == 6'd62);
  wire hmtqrdaxj62_sel = (r3ud3glj937o4_ == 6'd62);
  wire sbd346v9463_sel = (g5cld0_xqbmy2o0oiio_4 == 6'd63);
  wire hmtqrdaxj63_sel = (r3ud3glj937o4_ == 6'd63);

  wire sbd346v940_r;
  wire sbd346v940_nxt = pffig1fl4xtnw ? ~sbd346v940_r : ~c7sq9i2s8;
  wire sbd346v940_ena = (sbd346v940_sel & pffig1fl4xtnw) | (hmtqrdaxj0_sel & fpsdt9vdjcwssz9tezden07r7);
  ux607_gnrl_dfflr #(1) sbd346v940_dfflr (sbd346v940_ena, sbd346v940_nxt, sbd346v940_r, gf33atgy, ru_wi );
  wire sbd346v940_way0_we = sbd346v940_sel & ~sbd346v940_r;
  wire sbd346v940_way1_we = sbd346v940_sel &  sbd346v940_r;

  wire sbd346v941_r;
  wire sbd346v941_nxt = pffig1fl4xtnw ? ~sbd346v941_r : ~c7sq9i2s8;
  wire sbd346v941_ena = (sbd346v941_sel & pffig1fl4xtnw) | (hmtqrdaxj1_sel & fpsdt9vdjcwssz9tezden07r7);
  ux607_gnrl_dfflr #(1) sbd346v941_dfflr (sbd346v941_ena, sbd346v941_nxt, sbd346v941_r, gf33atgy, ru_wi );
  wire sbd346v941_way0_we = sbd346v941_sel & ~sbd346v941_r;
  wire sbd346v941_way1_we = sbd346v941_sel &  sbd346v941_r;

  wire sbd346v942_r;
  wire sbd346v942_nxt = pffig1fl4xtnw ? ~sbd346v942_r : ~c7sq9i2s8;
  wire sbd346v942_ena = (sbd346v942_sel & pffig1fl4xtnw) | (hmtqrdaxj2_sel & fpsdt9vdjcwssz9tezden07r7);
  ux607_gnrl_dfflr #(1) sbd346v942_dfflr (sbd346v942_ena, sbd346v942_nxt, sbd346v942_r, gf33atgy, ru_wi );
  wire sbd346v942_way0_we = sbd346v942_sel & ~sbd346v942_r;
  wire sbd346v942_way1_we = sbd346v942_sel &  sbd346v942_r;

  wire sbd346v943_r;
  wire sbd346v943_nxt = pffig1fl4xtnw ? ~sbd346v943_r : ~c7sq9i2s8;
  wire sbd346v943_ena = (sbd346v943_sel & pffig1fl4xtnw) | (hmtqrdaxj3_sel & fpsdt9vdjcwssz9tezden07r7);
  ux607_gnrl_dfflr #(1) sbd346v943_dfflr (sbd346v943_ena, sbd346v943_nxt, sbd346v943_r, gf33atgy, ru_wi );
  wire sbd346v943_way0_we = sbd346v943_sel & ~sbd346v943_r;
  wire sbd346v943_way1_we = sbd346v943_sel &  sbd346v943_r;

  wire sbd346v944_r;
  wire sbd346v944_nxt = pffig1fl4xtnw ? ~sbd346v944_r : ~c7sq9i2s8;
  wire sbd346v944_ena = (sbd346v944_sel & pffig1fl4xtnw) | (hmtqrdaxj4_sel & fpsdt9vdjcwssz9tezden07r7);
  ux607_gnrl_dfflr #(1) sbd346v944_dfflr (sbd346v944_ena, sbd346v944_nxt, sbd346v944_r, gf33atgy, ru_wi );
  wire sbd346v944_way0_we = sbd346v944_sel & ~sbd346v944_r;
  wire sbd346v944_way1_we = sbd346v944_sel &  sbd346v944_r;

  wire sbd346v945_r;
  wire sbd346v945_nxt = pffig1fl4xtnw ? ~sbd346v945_r : ~c7sq9i2s8;
  wire sbd346v945_ena = (sbd346v945_sel & pffig1fl4xtnw) | (hmtqrdaxj5_sel & fpsdt9vdjcwssz9tezden07r7);
  ux607_gnrl_dfflr #(1) sbd346v945_dfflr (sbd346v945_ena, sbd346v945_nxt, sbd346v945_r, gf33atgy, ru_wi );
  wire sbd346v945_way0_we = sbd346v945_sel & ~sbd346v945_r;
  wire sbd346v945_way1_we = sbd346v945_sel &  sbd346v945_r;

  wire sbd346v946_r;
  wire sbd346v946_nxt = pffig1fl4xtnw ? ~sbd346v946_r : ~c7sq9i2s8;
  wire sbd346v946_ena = (sbd346v946_sel & pffig1fl4xtnw) | (hmtqrdaxj6_sel & fpsdt9vdjcwssz9tezden07r7);
  ux607_gnrl_dfflr #(1) sbd346v946_dfflr (sbd346v946_ena, sbd346v946_nxt, sbd346v946_r, gf33atgy, ru_wi );
  wire sbd346v946_way0_we = sbd346v946_sel & ~sbd346v946_r;
  wire sbd346v946_way1_we = sbd346v946_sel &  sbd346v946_r;

  wire sbd346v947_r;
  wire sbd346v947_nxt = pffig1fl4xtnw ? ~sbd346v947_r : ~c7sq9i2s8;
  wire sbd346v947_ena = (sbd346v947_sel & pffig1fl4xtnw) | (hmtqrdaxj7_sel & fpsdt9vdjcwssz9tezden07r7);
  ux607_gnrl_dfflr #(1) sbd346v947_dfflr (sbd346v947_ena, sbd346v947_nxt, sbd346v947_r, gf33atgy, ru_wi );
  wire sbd346v947_way0_we = sbd346v947_sel & ~sbd346v947_r;
  wire sbd346v947_way1_we = sbd346v947_sel &  sbd346v947_r;

  wire sbd346v948_r;
  wire sbd346v948_nxt = pffig1fl4xtnw ? ~sbd346v948_r : ~c7sq9i2s8;
  wire sbd346v948_ena = (sbd346v948_sel & pffig1fl4xtnw) | (hmtqrdaxj8_sel & fpsdt9vdjcwssz9tezden07r7);
  ux607_gnrl_dfflr #(1) sbd346v948_dfflr (sbd346v948_ena, sbd346v948_nxt, sbd346v948_r, gf33atgy, ru_wi );
  wire sbd346v948_way0_we = sbd346v948_sel & ~sbd346v948_r;
  wire sbd346v948_way1_we = sbd346v948_sel &  sbd346v948_r;

  wire sbd346v949_r;
  wire sbd346v949_nxt = pffig1fl4xtnw ? ~sbd346v949_r : ~c7sq9i2s8;
  wire sbd346v949_ena = (sbd346v949_sel & pffig1fl4xtnw) | (hmtqrdaxj9_sel & fpsdt9vdjcwssz9tezden07r7);
  ux607_gnrl_dfflr #(1) sbd346v949_dfflr (sbd346v949_ena, sbd346v949_nxt, sbd346v949_r, gf33atgy, ru_wi );
  wire sbd346v949_way0_we = sbd346v949_sel & ~sbd346v949_r;
  wire sbd346v949_way1_we = sbd346v949_sel &  sbd346v949_r;

  wire sbd346v9410_r;
  wire sbd346v9410_nxt = pffig1fl4xtnw ? ~sbd346v9410_r : ~c7sq9i2s8;
  wire sbd346v9410_ena = (sbd346v9410_sel & pffig1fl4xtnw) | (hmtqrdaxj10_sel & fpsdt9vdjcwssz9tezden07r7);
  ux607_gnrl_dfflr #(1) sbd346v9410_dfflr (sbd346v9410_ena, sbd346v9410_nxt, sbd346v9410_r, gf33atgy, ru_wi );
  wire sbd346v9410_way0_we = sbd346v9410_sel & ~sbd346v9410_r;
  wire sbd346v9410_way1_we = sbd346v9410_sel &  sbd346v9410_r;

  wire sbd346v9411_r;
  wire sbd346v9411_nxt = pffig1fl4xtnw ? ~sbd346v9411_r : ~c7sq9i2s8;
  wire sbd346v9411_ena = (sbd346v9411_sel & pffig1fl4xtnw) | (hmtqrdaxj11_sel & fpsdt9vdjcwssz9tezden07r7);
  ux607_gnrl_dfflr #(1) sbd346v9411_dfflr (sbd346v9411_ena, sbd346v9411_nxt, sbd346v9411_r, gf33atgy, ru_wi );
  wire sbd346v9411_way0_we = sbd346v9411_sel & ~sbd346v9411_r;
  wire sbd346v9411_way1_we = sbd346v9411_sel &  sbd346v9411_r;

  wire sbd346v9412_r;
  wire sbd346v9412_nxt = pffig1fl4xtnw ? ~sbd346v9412_r : ~c7sq9i2s8;
  wire sbd346v9412_ena = (sbd346v9412_sel & pffig1fl4xtnw) | (hmtqrdaxj12_sel & fpsdt9vdjcwssz9tezden07r7);
  ux607_gnrl_dfflr #(1) sbd346v9412_dfflr (sbd346v9412_ena, sbd346v9412_nxt, sbd346v9412_r, gf33atgy, ru_wi );
  wire sbd346v9412_way0_we = sbd346v9412_sel & ~sbd346v9412_r;
  wire sbd346v9412_way1_we = sbd346v9412_sel &  sbd346v9412_r;

  wire sbd346v9413_r;
  wire sbd346v9413_nxt = pffig1fl4xtnw ? ~sbd346v9413_r : ~c7sq9i2s8;
  wire sbd346v9413_ena = (sbd346v9413_sel & pffig1fl4xtnw) | (hmtqrdaxj13_sel & fpsdt9vdjcwssz9tezden07r7);
  ux607_gnrl_dfflr #(1) sbd346v9413_dfflr (sbd346v9413_ena, sbd346v9413_nxt, sbd346v9413_r, gf33atgy, ru_wi );
  wire sbd346v9413_way0_we = sbd346v9413_sel & ~sbd346v9413_r;
  wire sbd346v9413_way1_we = sbd346v9413_sel &  sbd346v9413_r;

  wire sbd346v9414_r;
  wire sbd346v9414_nxt = pffig1fl4xtnw ? ~sbd346v9414_r : ~c7sq9i2s8;
  wire sbd346v9414_ena = (sbd346v9414_sel & pffig1fl4xtnw) | (hmtqrdaxj14_sel & fpsdt9vdjcwssz9tezden07r7);
  ux607_gnrl_dfflr #(1) sbd346v9414_dfflr (sbd346v9414_ena, sbd346v9414_nxt, sbd346v9414_r, gf33atgy, ru_wi );
  wire sbd346v9414_way0_we = sbd346v9414_sel & ~sbd346v9414_r;
  wire sbd346v9414_way1_we = sbd346v9414_sel &  sbd346v9414_r;

  wire sbd346v9415_r;
  wire sbd346v9415_nxt = pffig1fl4xtnw ? ~sbd346v9415_r : ~c7sq9i2s8;
  wire sbd346v9415_ena = (sbd346v9415_sel & pffig1fl4xtnw) | (hmtqrdaxj15_sel & fpsdt9vdjcwssz9tezden07r7);
  ux607_gnrl_dfflr #(1) sbd346v9415_dfflr (sbd346v9415_ena, sbd346v9415_nxt, sbd346v9415_r, gf33atgy, ru_wi );
  wire sbd346v9415_way0_we = sbd346v9415_sel & ~sbd346v9415_r;
  wire sbd346v9415_way1_we = sbd346v9415_sel &  sbd346v9415_r;

  wire sbd346v9416_r;
  wire sbd346v9416_nxt = pffig1fl4xtnw ? ~sbd346v9416_r : ~c7sq9i2s8;
  wire sbd346v9416_ena = (sbd346v9416_sel & pffig1fl4xtnw) | (hmtqrdaxj16_sel & fpsdt9vdjcwssz9tezden07r7);
  ux607_gnrl_dfflr #(1) sbd346v9416_dfflr (sbd346v9416_ena, sbd346v9416_nxt, sbd346v9416_r, gf33atgy, ru_wi );
  wire sbd346v9416_way0_we = sbd346v9416_sel & ~sbd346v9416_r;
  wire sbd346v9416_way1_we = sbd346v9416_sel &  sbd346v9416_r;

  wire sbd346v9417_r;
  wire sbd346v9417_nxt = pffig1fl4xtnw ? ~sbd346v9417_r : ~c7sq9i2s8;
  wire sbd346v9417_ena = (sbd346v9417_sel & pffig1fl4xtnw) | (hmtqrdaxj17_sel & fpsdt9vdjcwssz9tezden07r7);
  ux607_gnrl_dfflr #(1) sbd346v9417_dfflr (sbd346v9417_ena, sbd346v9417_nxt, sbd346v9417_r, gf33atgy, ru_wi );
  wire sbd346v9417_way0_we = sbd346v9417_sel & ~sbd346v9417_r;
  wire sbd346v9417_way1_we = sbd346v9417_sel &  sbd346v9417_r;

  wire sbd346v9418_r;
  wire sbd346v9418_nxt = pffig1fl4xtnw ? ~sbd346v9418_r : ~c7sq9i2s8;
  wire sbd346v9418_ena = (sbd346v9418_sel & pffig1fl4xtnw) | (hmtqrdaxj18_sel & fpsdt9vdjcwssz9tezden07r7);
  ux607_gnrl_dfflr #(1) sbd346v9418_dfflr (sbd346v9418_ena, sbd346v9418_nxt, sbd346v9418_r, gf33atgy, ru_wi );
  wire sbd346v9418_way0_we = sbd346v9418_sel & ~sbd346v9418_r;
  wire sbd346v9418_way1_we = sbd346v9418_sel &  sbd346v9418_r;

  wire sbd346v9419_r;
  wire sbd346v9419_nxt = pffig1fl4xtnw ? ~sbd346v9419_r : ~c7sq9i2s8;
  wire sbd346v9419_ena = (sbd346v9419_sel & pffig1fl4xtnw) | (hmtqrdaxj19_sel & fpsdt9vdjcwssz9tezden07r7);
  ux607_gnrl_dfflr #(1) sbd346v9419_dfflr (sbd346v9419_ena, sbd346v9419_nxt, sbd346v9419_r, gf33atgy, ru_wi );
  wire sbd346v9419_way0_we = sbd346v9419_sel & ~sbd346v9419_r;
  wire sbd346v9419_way1_we = sbd346v9419_sel &  sbd346v9419_r;

  wire sbd346v9420_r;
  wire sbd346v9420_nxt = pffig1fl4xtnw ? ~sbd346v9420_r : ~c7sq9i2s8;
  wire sbd346v9420_ena = (sbd346v9420_sel & pffig1fl4xtnw) | (hmtqrdaxj20_sel & fpsdt9vdjcwssz9tezden07r7);
  ux607_gnrl_dfflr #(1) sbd346v9420_dfflr (sbd346v9420_ena, sbd346v9420_nxt, sbd346v9420_r, gf33atgy, ru_wi );
  wire sbd346v9420_way0_we = sbd346v9420_sel & ~sbd346v9420_r;
  wire sbd346v9420_way1_we = sbd346v9420_sel &  sbd346v9420_r;

  wire sbd346v9421_r;
  wire sbd346v9421_nxt = pffig1fl4xtnw ? ~sbd346v9421_r : ~c7sq9i2s8;
  wire sbd346v9421_ena = (sbd346v9421_sel & pffig1fl4xtnw) | (hmtqrdaxj21_sel & fpsdt9vdjcwssz9tezden07r7);
  ux607_gnrl_dfflr #(1) sbd346v9421_dfflr (sbd346v9421_ena, sbd346v9421_nxt, sbd346v9421_r, gf33atgy, ru_wi );
  wire sbd346v9421_way0_we = sbd346v9421_sel & ~sbd346v9421_r;
  wire sbd346v9421_way1_we = sbd346v9421_sel &  sbd346v9421_r;

  wire sbd346v9422_r;
  wire sbd346v9422_nxt = pffig1fl4xtnw ? ~sbd346v9422_r : ~c7sq9i2s8;
  wire sbd346v9422_ena = (sbd346v9422_sel & pffig1fl4xtnw) | (hmtqrdaxj22_sel & fpsdt9vdjcwssz9tezden07r7);
  ux607_gnrl_dfflr #(1) sbd346v9422_dfflr (sbd346v9422_ena, sbd346v9422_nxt, sbd346v9422_r, gf33atgy, ru_wi );
  wire sbd346v9422_way0_we = sbd346v9422_sel & ~sbd346v9422_r;
  wire sbd346v9422_way1_we = sbd346v9422_sel &  sbd346v9422_r;

  wire sbd346v9423_r;
  wire sbd346v9423_nxt = pffig1fl4xtnw ? ~sbd346v9423_r : ~c7sq9i2s8;
  wire sbd346v9423_ena = (sbd346v9423_sel & pffig1fl4xtnw) | (hmtqrdaxj23_sel & fpsdt9vdjcwssz9tezden07r7);
  ux607_gnrl_dfflr #(1) sbd346v9423_dfflr (sbd346v9423_ena, sbd346v9423_nxt, sbd346v9423_r, gf33atgy, ru_wi );
  wire sbd346v9423_way0_we = sbd346v9423_sel & ~sbd346v9423_r;
  wire sbd346v9423_way1_we = sbd346v9423_sel &  sbd346v9423_r;

  wire sbd346v9424_r;
  wire sbd346v9424_nxt = pffig1fl4xtnw ? ~sbd346v9424_r : ~c7sq9i2s8;
  wire sbd346v9424_ena = (sbd346v9424_sel & pffig1fl4xtnw) | (hmtqrdaxj24_sel & fpsdt9vdjcwssz9tezden07r7);
  ux607_gnrl_dfflr #(1) sbd346v9424_dfflr (sbd346v9424_ena, sbd346v9424_nxt, sbd346v9424_r, gf33atgy, ru_wi );
  wire sbd346v9424_way0_we = sbd346v9424_sel & ~sbd346v9424_r;
  wire sbd346v9424_way1_we = sbd346v9424_sel &  sbd346v9424_r;

  wire sbd346v9425_r;
  wire sbd346v9425_nxt = pffig1fl4xtnw ? ~sbd346v9425_r : ~c7sq9i2s8;
  wire sbd346v9425_ena = (sbd346v9425_sel & pffig1fl4xtnw) | (hmtqrdaxj25_sel & fpsdt9vdjcwssz9tezden07r7);
  ux607_gnrl_dfflr #(1) sbd346v9425_dfflr (sbd346v9425_ena, sbd346v9425_nxt, sbd346v9425_r, gf33atgy, ru_wi );
  wire sbd346v9425_way0_we = sbd346v9425_sel & ~sbd346v9425_r;
  wire sbd346v9425_way1_we = sbd346v9425_sel &  sbd346v9425_r;

  wire sbd346v9426_r;
  wire sbd346v9426_nxt = pffig1fl4xtnw ? ~sbd346v9426_r : ~c7sq9i2s8;
  wire sbd346v9426_ena = (sbd346v9426_sel & pffig1fl4xtnw) | (hmtqrdaxj26_sel & fpsdt9vdjcwssz9tezden07r7);
  ux607_gnrl_dfflr #(1) sbd346v9426_dfflr (sbd346v9426_ena, sbd346v9426_nxt, sbd346v9426_r, gf33atgy, ru_wi );
  wire sbd346v9426_way0_we = sbd346v9426_sel & ~sbd346v9426_r;
  wire sbd346v9426_way1_we = sbd346v9426_sel &  sbd346v9426_r;

  wire sbd346v9427_r;
  wire sbd346v9427_nxt = pffig1fl4xtnw ? ~sbd346v9427_r : ~c7sq9i2s8;
  wire sbd346v9427_ena = (sbd346v9427_sel & pffig1fl4xtnw) | (hmtqrdaxj27_sel & fpsdt9vdjcwssz9tezden07r7);
  ux607_gnrl_dfflr #(1) sbd346v9427_dfflr (sbd346v9427_ena, sbd346v9427_nxt, sbd346v9427_r, gf33atgy, ru_wi );
  wire sbd346v9427_way0_we = sbd346v9427_sel & ~sbd346v9427_r;
  wire sbd346v9427_way1_we = sbd346v9427_sel &  sbd346v9427_r;

  wire sbd346v9428_r;
  wire sbd346v9428_nxt = pffig1fl4xtnw ? ~sbd346v9428_r : ~c7sq9i2s8;
  wire sbd346v9428_ena = (sbd346v9428_sel & pffig1fl4xtnw) | (hmtqrdaxj28_sel & fpsdt9vdjcwssz9tezden07r7);
  ux607_gnrl_dfflr #(1) sbd346v9428_dfflr (sbd346v9428_ena, sbd346v9428_nxt, sbd346v9428_r, gf33atgy, ru_wi );
  wire sbd346v9428_way0_we = sbd346v9428_sel & ~sbd346v9428_r;
  wire sbd346v9428_way1_we = sbd346v9428_sel &  sbd346v9428_r;

  wire sbd346v9429_r;
  wire sbd346v9429_nxt = pffig1fl4xtnw ? ~sbd346v9429_r : ~c7sq9i2s8;
  wire sbd346v9429_ena = (sbd346v9429_sel & pffig1fl4xtnw) | (hmtqrdaxj29_sel & fpsdt9vdjcwssz9tezden07r7);
  ux607_gnrl_dfflr #(1) sbd346v9429_dfflr (sbd346v9429_ena, sbd346v9429_nxt, sbd346v9429_r, gf33atgy, ru_wi );
  wire sbd346v9429_way0_we = sbd346v9429_sel & ~sbd346v9429_r;
  wire sbd346v9429_way1_we = sbd346v9429_sel &  sbd346v9429_r;

  wire sbd346v9430_r;
  wire sbd346v9430_nxt = pffig1fl4xtnw ? ~sbd346v9430_r : ~c7sq9i2s8;
  wire sbd346v9430_ena = (sbd346v9430_sel & pffig1fl4xtnw) | (hmtqrdaxj30_sel & fpsdt9vdjcwssz9tezden07r7);
  ux607_gnrl_dfflr #(1) sbd346v9430_dfflr (sbd346v9430_ena, sbd346v9430_nxt, sbd346v9430_r, gf33atgy, ru_wi );
  wire sbd346v9430_way0_we = sbd346v9430_sel & ~sbd346v9430_r;
  wire sbd346v9430_way1_we = sbd346v9430_sel &  sbd346v9430_r;

  wire sbd346v9431_r;
  wire sbd346v9431_nxt = pffig1fl4xtnw ? ~sbd346v9431_r : ~c7sq9i2s8;
  wire sbd346v9431_ena = (sbd346v9431_sel & pffig1fl4xtnw) | (hmtqrdaxj31_sel & fpsdt9vdjcwssz9tezden07r7);
  ux607_gnrl_dfflr #(1) sbd346v9431_dfflr (sbd346v9431_ena, sbd346v9431_nxt, sbd346v9431_r, gf33atgy, ru_wi );
  wire sbd346v9431_way0_we = sbd346v9431_sel & ~sbd346v9431_r;
  wire sbd346v9431_way1_we = sbd346v9431_sel &  sbd346v9431_r;

  wire sbd346v9432_r;
  wire sbd346v9432_nxt = pffig1fl4xtnw ? ~sbd346v9432_r : ~c7sq9i2s8;
  wire sbd346v9432_ena = (sbd346v9432_sel & pffig1fl4xtnw) | (hmtqrdaxj32_sel & fpsdt9vdjcwssz9tezden07r7);
  ux607_gnrl_dfflr #(1) sbd346v9432_dfflr (sbd346v9432_ena, sbd346v9432_nxt, sbd346v9432_r, gf33atgy, ru_wi );
  wire sbd346v9432_way0_we = sbd346v9432_sel & ~sbd346v9432_r;
  wire sbd346v9432_way1_we = sbd346v9432_sel &  sbd346v9432_r;

  wire sbd346v9433_r;
  wire sbd346v9433_nxt = pffig1fl4xtnw ? ~sbd346v9433_r : ~c7sq9i2s8;
  wire sbd346v9433_ena = (sbd346v9433_sel & pffig1fl4xtnw) | (hmtqrdaxj33_sel & fpsdt9vdjcwssz9tezden07r7);
  ux607_gnrl_dfflr #(1) sbd346v9433_dfflr (sbd346v9433_ena, sbd346v9433_nxt, sbd346v9433_r, gf33atgy, ru_wi );
  wire sbd346v9433_way0_we = sbd346v9433_sel & ~sbd346v9433_r;
  wire sbd346v9433_way1_we = sbd346v9433_sel &  sbd346v9433_r;

  wire sbd346v9434_r;
  wire sbd346v9434_nxt = pffig1fl4xtnw ? ~sbd346v9434_r : ~c7sq9i2s8;
  wire sbd346v9434_ena = (sbd346v9434_sel & pffig1fl4xtnw) | (hmtqrdaxj34_sel & fpsdt9vdjcwssz9tezden07r7);
  ux607_gnrl_dfflr #(1) sbd346v9434_dfflr (sbd346v9434_ena, sbd346v9434_nxt, sbd346v9434_r, gf33atgy, ru_wi );
  wire sbd346v9434_way0_we = sbd346v9434_sel & ~sbd346v9434_r;
  wire sbd346v9434_way1_we = sbd346v9434_sel &  sbd346v9434_r;

  wire sbd346v9435_r;
  wire sbd346v9435_nxt = pffig1fl4xtnw ? ~sbd346v9435_r : ~c7sq9i2s8;
  wire sbd346v9435_ena = (sbd346v9435_sel & pffig1fl4xtnw) | (hmtqrdaxj35_sel & fpsdt9vdjcwssz9tezden07r7);
  ux607_gnrl_dfflr #(1) sbd346v9435_dfflr (sbd346v9435_ena, sbd346v9435_nxt, sbd346v9435_r, gf33atgy, ru_wi );
  wire sbd346v9435_way0_we = sbd346v9435_sel & ~sbd346v9435_r;
  wire sbd346v9435_way1_we = sbd346v9435_sel &  sbd346v9435_r;

  wire sbd346v9436_r;
  wire sbd346v9436_nxt = pffig1fl4xtnw ? ~sbd346v9436_r : ~c7sq9i2s8;
  wire sbd346v9436_ena = (sbd346v9436_sel & pffig1fl4xtnw) | (hmtqrdaxj36_sel & fpsdt9vdjcwssz9tezden07r7);
  ux607_gnrl_dfflr #(1) sbd346v9436_dfflr (sbd346v9436_ena, sbd346v9436_nxt, sbd346v9436_r, gf33atgy, ru_wi );
  wire sbd346v9436_way0_we = sbd346v9436_sel & ~sbd346v9436_r;
  wire sbd346v9436_way1_we = sbd346v9436_sel &  sbd346v9436_r;

  wire sbd346v9437_r;
  wire sbd346v9437_nxt = pffig1fl4xtnw ? ~sbd346v9437_r : ~c7sq9i2s8;
  wire sbd346v9437_ena = (sbd346v9437_sel & pffig1fl4xtnw) | (hmtqrdaxj37_sel & fpsdt9vdjcwssz9tezden07r7);
  ux607_gnrl_dfflr #(1) sbd346v9437_dfflr (sbd346v9437_ena, sbd346v9437_nxt, sbd346v9437_r, gf33atgy, ru_wi );
  wire sbd346v9437_way0_we = sbd346v9437_sel & ~sbd346v9437_r;
  wire sbd346v9437_way1_we = sbd346v9437_sel &  sbd346v9437_r;

  wire sbd346v9438_r;
  wire sbd346v9438_nxt = pffig1fl4xtnw ? ~sbd346v9438_r : ~c7sq9i2s8;
  wire sbd346v9438_ena = (sbd346v9438_sel & pffig1fl4xtnw) | (hmtqrdaxj38_sel & fpsdt9vdjcwssz9tezden07r7);
  ux607_gnrl_dfflr #(1) sbd346v9438_dfflr (sbd346v9438_ena, sbd346v9438_nxt, sbd346v9438_r, gf33atgy, ru_wi );
  wire sbd346v9438_way0_we = sbd346v9438_sel & ~sbd346v9438_r;
  wire sbd346v9438_way1_we = sbd346v9438_sel &  sbd346v9438_r;

  wire sbd346v9439_r;
  wire sbd346v9439_nxt = pffig1fl4xtnw ? ~sbd346v9439_r : ~c7sq9i2s8;
  wire sbd346v9439_ena = (sbd346v9439_sel & pffig1fl4xtnw) | (hmtqrdaxj39_sel & fpsdt9vdjcwssz9tezden07r7);
  ux607_gnrl_dfflr #(1) sbd346v9439_dfflr (sbd346v9439_ena, sbd346v9439_nxt, sbd346v9439_r, gf33atgy, ru_wi );
  wire sbd346v9439_way0_we = sbd346v9439_sel & ~sbd346v9439_r;
  wire sbd346v9439_way1_we = sbd346v9439_sel &  sbd346v9439_r;

  wire sbd346v9440_r;
  wire sbd346v9440_nxt = pffig1fl4xtnw ? ~sbd346v9440_r : ~c7sq9i2s8;
  wire sbd346v9440_ena = (sbd346v9440_sel & pffig1fl4xtnw) | (hmtqrdaxj40_sel & fpsdt9vdjcwssz9tezden07r7);
  ux607_gnrl_dfflr #(1) sbd346v9440_dfflr (sbd346v9440_ena, sbd346v9440_nxt, sbd346v9440_r, gf33atgy, ru_wi );
  wire sbd346v9440_way0_we = sbd346v9440_sel & ~sbd346v9440_r;
  wire sbd346v9440_way1_we = sbd346v9440_sel &  sbd346v9440_r;

  wire sbd346v9441_r;
  wire sbd346v9441_nxt = pffig1fl4xtnw ? ~sbd346v9441_r : ~c7sq9i2s8;
  wire sbd346v9441_ena = (sbd346v9441_sel & pffig1fl4xtnw) | (hmtqrdaxj41_sel & fpsdt9vdjcwssz9tezden07r7);
  ux607_gnrl_dfflr #(1) sbd346v9441_dfflr (sbd346v9441_ena, sbd346v9441_nxt, sbd346v9441_r, gf33atgy, ru_wi );
  wire sbd346v9441_way0_we = sbd346v9441_sel & ~sbd346v9441_r;
  wire sbd346v9441_way1_we = sbd346v9441_sel &  sbd346v9441_r;

  wire sbd346v9442_r;
  wire sbd346v9442_nxt = pffig1fl4xtnw ? ~sbd346v9442_r : ~c7sq9i2s8;
  wire sbd346v9442_ena = (sbd346v9442_sel & pffig1fl4xtnw) | (hmtqrdaxj42_sel & fpsdt9vdjcwssz9tezden07r7);
  ux607_gnrl_dfflr #(1) sbd346v9442_dfflr (sbd346v9442_ena, sbd346v9442_nxt, sbd346v9442_r, gf33atgy, ru_wi );
  wire sbd346v9442_way0_we = sbd346v9442_sel & ~sbd346v9442_r;
  wire sbd346v9442_way1_we = sbd346v9442_sel &  sbd346v9442_r;

  wire sbd346v9443_r;
  wire sbd346v9443_nxt = pffig1fl4xtnw ? ~sbd346v9443_r : ~c7sq9i2s8;
  wire sbd346v9443_ena = (sbd346v9443_sel & pffig1fl4xtnw) | (hmtqrdaxj43_sel & fpsdt9vdjcwssz9tezden07r7);
  ux607_gnrl_dfflr #(1) sbd346v9443_dfflr (sbd346v9443_ena, sbd346v9443_nxt, sbd346v9443_r, gf33atgy, ru_wi );
  wire sbd346v9443_way0_we = sbd346v9443_sel & ~sbd346v9443_r;
  wire sbd346v9443_way1_we = sbd346v9443_sel &  sbd346v9443_r;

  wire sbd346v9444_r;
  wire sbd346v9444_nxt = pffig1fl4xtnw ? ~sbd346v9444_r : ~c7sq9i2s8;
  wire sbd346v9444_ena = (sbd346v9444_sel & pffig1fl4xtnw) | (hmtqrdaxj44_sel & fpsdt9vdjcwssz9tezden07r7);
  ux607_gnrl_dfflr #(1) sbd346v9444_dfflr (sbd346v9444_ena, sbd346v9444_nxt, sbd346v9444_r, gf33atgy, ru_wi );
  wire sbd346v9444_way0_we = sbd346v9444_sel & ~sbd346v9444_r;
  wire sbd346v9444_way1_we = sbd346v9444_sel &  sbd346v9444_r;

  wire sbd346v9445_r;
  wire sbd346v9445_nxt = pffig1fl4xtnw ? ~sbd346v9445_r : ~c7sq9i2s8;
  wire sbd346v9445_ena = (sbd346v9445_sel & pffig1fl4xtnw) | (hmtqrdaxj45_sel & fpsdt9vdjcwssz9tezden07r7);
  ux607_gnrl_dfflr #(1) sbd346v9445_dfflr (sbd346v9445_ena, sbd346v9445_nxt, sbd346v9445_r, gf33atgy, ru_wi );
  wire sbd346v9445_way0_we = sbd346v9445_sel & ~sbd346v9445_r;
  wire sbd346v9445_way1_we = sbd346v9445_sel &  sbd346v9445_r;

  wire sbd346v9446_r;
  wire sbd346v9446_nxt = pffig1fl4xtnw ? ~sbd346v9446_r : ~c7sq9i2s8;
  wire sbd346v9446_ena = (sbd346v9446_sel & pffig1fl4xtnw) | (hmtqrdaxj46_sel & fpsdt9vdjcwssz9tezden07r7);
  ux607_gnrl_dfflr #(1) sbd346v9446_dfflr (sbd346v9446_ena, sbd346v9446_nxt, sbd346v9446_r, gf33atgy, ru_wi );
  wire sbd346v9446_way0_we = sbd346v9446_sel & ~sbd346v9446_r;
  wire sbd346v9446_way1_we = sbd346v9446_sel &  sbd346v9446_r;

  wire sbd346v9447_r;
  wire sbd346v9447_nxt = pffig1fl4xtnw ? ~sbd346v9447_r : ~c7sq9i2s8;
  wire sbd346v9447_ena = (sbd346v9447_sel & pffig1fl4xtnw) | (hmtqrdaxj47_sel & fpsdt9vdjcwssz9tezden07r7);
  ux607_gnrl_dfflr #(1) sbd346v9447_dfflr (sbd346v9447_ena, sbd346v9447_nxt, sbd346v9447_r, gf33atgy, ru_wi );
  wire sbd346v9447_way0_we = sbd346v9447_sel & ~sbd346v9447_r;
  wire sbd346v9447_way1_we = sbd346v9447_sel &  sbd346v9447_r;

  wire sbd346v9448_r;
  wire sbd346v9448_nxt = pffig1fl4xtnw ? ~sbd346v9448_r : ~c7sq9i2s8;
  wire sbd346v9448_ena = (sbd346v9448_sel & pffig1fl4xtnw) | (hmtqrdaxj48_sel & fpsdt9vdjcwssz9tezden07r7);
  ux607_gnrl_dfflr #(1) sbd346v9448_dfflr (sbd346v9448_ena, sbd346v9448_nxt, sbd346v9448_r, gf33atgy, ru_wi );
  wire sbd346v9448_way0_we = sbd346v9448_sel & ~sbd346v9448_r;
  wire sbd346v9448_way1_we = sbd346v9448_sel &  sbd346v9448_r;

  wire sbd346v9449_r;
  wire sbd346v9449_nxt = pffig1fl4xtnw ? ~sbd346v9449_r : ~c7sq9i2s8;
  wire sbd346v9449_ena = (sbd346v9449_sel & pffig1fl4xtnw) | (hmtqrdaxj49_sel & fpsdt9vdjcwssz9tezden07r7);
  ux607_gnrl_dfflr #(1) sbd346v9449_dfflr (sbd346v9449_ena, sbd346v9449_nxt, sbd346v9449_r, gf33atgy, ru_wi );
  wire sbd346v9449_way0_we = sbd346v9449_sel & ~sbd346v9449_r;
  wire sbd346v9449_way1_we = sbd346v9449_sel &  sbd346v9449_r;

  wire sbd346v9450_r;
  wire sbd346v9450_nxt = pffig1fl4xtnw ? ~sbd346v9450_r : ~c7sq9i2s8;
  wire sbd346v9450_ena = (sbd346v9450_sel & pffig1fl4xtnw) | (hmtqrdaxj50_sel & fpsdt9vdjcwssz9tezden07r7);
  ux607_gnrl_dfflr #(1) sbd346v9450_dfflr (sbd346v9450_ena, sbd346v9450_nxt, sbd346v9450_r, gf33atgy, ru_wi );
  wire sbd346v9450_way0_we = sbd346v9450_sel & ~sbd346v9450_r;
  wire sbd346v9450_way1_we = sbd346v9450_sel &  sbd346v9450_r;

  wire sbd346v9451_r;
  wire sbd346v9451_nxt = pffig1fl4xtnw ? ~sbd346v9451_r : ~c7sq9i2s8;
  wire sbd346v9451_ena = (sbd346v9451_sel & pffig1fl4xtnw) | (hmtqrdaxj51_sel & fpsdt9vdjcwssz9tezden07r7);
  ux607_gnrl_dfflr #(1) sbd346v9451_dfflr (sbd346v9451_ena, sbd346v9451_nxt, sbd346v9451_r, gf33atgy, ru_wi );
  wire sbd346v9451_way0_we = sbd346v9451_sel & ~sbd346v9451_r;
  wire sbd346v9451_way1_we = sbd346v9451_sel &  sbd346v9451_r;

  wire sbd346v9452_r;
  wire sbd346v9452_nxt = pffig1fl4xtnw ? ~sbd346v9452_r : ~c7sq9i2s8;
  wire sbd346v9452_ena = (sbd346v9452_sel & pffig1fl4xtnw) | (hmtqrdaxj52_sel & fpsdt9vdjcwssz9tezden07r7);
  ux607_gnrl_dfflr #(1) sbd346v9452_dfflr (sbd346v9452_ena, sbd346v9452_nxt, sbd346v9452_r, gf33atgy, ru_wi );
  wire sbd346v9452_way0_we = sbd346v9452_sel & ~sbd346v9452_r;
  wire sbd346v9452_way1_we = sbd346v9452_sel &  sbd346v9452_r;

  wire sbd346v9453_r;
  wire sbd346v9453_nxt = pffig1fl4xtnw ? ~sbd346v9453_r : ~c7sq9i2s8;
  wire sbd346v9453_ena = (sbd346v9453_sel & pffig1fl4xtnw) | (hmtqrdaxj53_sel & fpsdt9vdjcwssz9tezden07r7);
  ux607_gnrl_dfflr #(1) sbd346v9453_dfflr (sbd346v9453_ena, sbd346v9453_nxt, sbd346v9453_r, gf33atgy, ru_wi );
  wire sbd346v9453_way0_we = sbd346v9453_sel & ~sbd346v9453_r;
  wire sbd346v9453_way1_we = sbd346v9453_sel &  sbd346v9453_r;

  wire sbd346v9454_r;
  wire sbd346v9454_nxt = pffig1fl4xtnw ? ~sbd346v9454_r : ~c7sq9i2s8;
  wire sbd346v9454_ena = (sbd346v9454_sel & pffig1fl4xtnw) | (hmtqrdaxj54_sel & fpsdt9vdjcwssz9tezden07r7);
  ux607_gnrl_dfflr #(1) sbd346v9454_dfflr (sbd346v9454_ena, sbd346v9454_nxt, sbd346v9454_r, gf33atgy, ru_wi );
  wire sbd346v9454_way0_we = sbd346v9454_sel & ~sbd346v9454_r;
  wire sbd346v9454_way1_we = sbd346v9454_sel &  sbd346v9454_r;

  wire sbd346v9455_r;
  wire sbd346v9455_nxt = pffig1fl4xtnw ? ~sbd346v9455_r : ~c7sq9i2s8;
  wire sbd346v9455_ena = (sbd346v9455_sel & pffig1fl4xtnw) | (hmtqrdaxj55_sel & fpsdt9vdjcwssz9tezden07r7);
  ux607_gnrl_dfflr #(1) sbd346v9455_dfflr (sbd346v9455_ena, sbd346v9455_nxt, sbd346v9455_r, gf33atgy, ru_wi );
  wire sbd346v9455_way0_we = sbd346v9455_sel & ~sbd346v9455_r;
  wire sbd346v9455_way1_we = sbd346v9455_sel &  sbd346v9455_r;

  wire sbd346v9456_r;
  wire sbd346v9456_nxt = pffig1fl4xtnw ? ~sbd346v9456_r : ~c7sq9i2s8;
  wire sbd346v9456_ena = (sbd346v9456_sel & pffig1fl4xtnw) | (hmtqrdaxj56_sel & fpsdt9vdjcwssz9tezden07r7);
  ux607_gnrl_dfflr #(1) sbd346v9456_dfflr (sbd346v9456_ena, sbd346v9456_nxt, sbd346v9456_r, gf33atgy, ru_wi );
  wire sbd346v9456_way0_we = sbd346v9456_sel & ~sbd346v9456_r;
  wire sbd346v9456_way1_we = sbd346v9456_sel &  sbd346v9456_r;

  wire sbd346v9457_r;
  wire sbd346v9457_nxt = pffig1fl4xtnw ? ~sbd346v9457_r : ~c7sq9i2s8;
  wire sbd346v9457_ena = (sbd346v9457_sel & pffig1fl4xtnw) | (hmtqrdaxj57_sel & fpsdt9vdjcwssz9tezden07r7);
  ux607_gnrl_dfflr #(1) sbd346v9457_dfflr (sbd346v9457_ena, sbd346v9457_nxt, sbd346v9457_r, gf33atgy, ru_wi );
  wire sbd346v9457_way0_we = sbd346v9457_sel & ~sbd346v9457_r;
  wire sbd346v9457_way1_we = sbd346v9457_sel &  sbd346v9457_r;

  wire sbd346v9458_r;
  wire sbd346v9458_nxt = pffig1fl4xtnw ? ~sbd346v9458_r : ~c7sq9i2s8;
  wire sbd346v9458_ena = (sbd346v9458_sel & pffig1fl4xtnw) | (hmtqrdaxj58_sel & fpsdt9vdjcwssz9tezden07r7);
  ux607_gnrl_dfflr #(1) sbd346v9458_dfflr (sbd346v9458_ena, sbd346v9458_nxt, sbd346v9458_r, gf33atgy, ru_wi );
  wire sbd346v9458_way0_we = sbd346v9458_sel & ~sbd346v9458_r;
  wire sbd346v9458_way1_we = sbd346v9458_sel &  sbd346v9458_r;

  wire sbd346v9459_r;
  wire sbd346v9459_nxt = pffig1fl4xtnw ? ~sbd346v9459_r : ~c7sq9i2s8;
  wire sbd346v9459_ena = (sbd346v9459_sel & pffig1fl4xtnw) | (hmtqrdaxj59_sel & fpsdt9vdjcwssz9tezden07r7);
  ux607_gnrl_dfflr #(1) sbd346v9459_dfflr (sbd346v9459_ena, sbd346v9459_nxt, sbd346v9459_r, gf33atgy, ru_wi );
  wire sbd346v9459_way0_we = sbd346v9459_sel & ~sbd346v9459_r;
  wire sbd346v9459_way1_we = sbd346v9459_sel &  sbd346v9459_r;

  wire sbd346v9460_r;
  wire sbd346v9460_nxt = pffig1fl4xtnw ? ~sbd346v9460_r : ~c7sq9i2s8;
  wire sbd346v9460_ena = (sbd346v9460_sel & pffig1fl4xtnw) | (hmtqrdaxj60_sel & fpsdt9vdjcwssz9tezden07r7);
  ux607_gnrl_dfflr #(1) sbd346v9460_dfflr (sbd346v9460_ena, sbd346v9460_nxt, sbd346v9460_r, gf33atgy, ru_wi );
  wire sbd346v9460_way0_we = sbd346v9460_sel & ~sbd346v9460_r;
  wire sbd346v9460_way1_we = sbd346v9460_sel &  sbd346v9460_r;

  wire sbd346v9461_r;
  wire sbd346v9461_nxt = pffig1fl4xtnw ? ~sbd346v9461_r : ~c7sq9i2s8;
  wire sbd346v9461_ena = (sbd346v9461_sel & pffig1fl4xtnw) | (hmtqrdaxj61_sel & fpsdt9vdjcwssz9tezden07r7);
  ux607_gnrl_dfflr #(1) sbd346v9461_dfflr (sbd346v9461_ena, sbd346v9461_nxt, sbd346v9461_r, gf33atgy, ru_wi );
  wire sbd346v9461_way0_we = sbd346v9461_sel & ~sbd346v9461_r;
  wire sbd346v9461_way1_we = sbd346v9461_sel &  sbd346v9461_r;

  wire sbd346v9462_r;
  wire sbd346v9462_nxt = pffig1fl4xtnw ? ~sbd346v9462_r : ~c7sq9i2s8;
  wire sbd346v9462_ena = (sbd346v9462_sel & pffig1fl4xtnw) | (hmtqrdaxj62_sel & fpsdt9vdjcwssz9tezden07r7);
  ux607_gnrl_dfflr #(1) sbd346v9462_dfflr (sbd346v9462_ena, sbd346v9462_nxt, sbd346v9462_r, gf33atgy, ru_wi );
  wire sbd346v9462_way0_we = sbd346v9462_sel & ~sbd346v9462_r;
  wire sbd346v9462_way1_we = sbd346v9462_sel &  sbd346v9462_r;

  wire sbd346v9463_r;
  wire sbd346v9463_nxt = pffig1fl4xtnw ? ~sbd346v9463_r : ~c7sq9i2s8;
  wire sbd346v9463_ena = (sbd346v9463_sel & pffig1fl4xtnw) | (hmtqrdaxj63_sel & fpsdt9vdjcwssz9tezden07r7);
  ux607_gnrl_dfflr #(1) sbd346v9463_dfflr (sbd346v9463_ena, sbd346v9463_nxt, sbd346v9463_r, gf33atgy, ru_wi );
  wire sbd346v9463_way0_we = sbd346v9463_sel & ~sbd346v9463_r;
  wire sbd346v9463_way1_we = sbd346v9463_sel &  sbd346v9463_r;

  
  wire wlxoaneirix6ez6fhtyv3os9c3 = 1'b0 
                              | sbd346v940_way0_we 
                              | sbd346v941_way0_we 
                              | sbd346v942_way0_we 
                              | sbd346v943_way0_we 
                              | sbd346v944_way0_we 
                              | sbd346v945_way0_we 
                              | sbd346v946_way0_we 
                              | sbd346v947_way0_we 
                              | sbd346v948_way0_we 
                              | sbd346v949_way0_we 
                              | sbd346v9410_way0_we 
                              | sbd346v9411_way0_we 
                              | sbd346v9412_way0_we 
                              | sbd346v9413_way0_we 
                              | sbd346v9414_way0_we 
                              | sbd346v9415_way0_we 
                              | sbd346v9416_way0_we 
                              | sbd346v9417_way0_we 
                              | sbd346v9418_way0_we 
                              | sbd346v9419_way0_we 
                              | sbd346v9420_way0_we 
                              | sbd346v9421_way0_we 
                              | sbd346v9422_way0_we 
                              | sbd346v9423_way0_we 
                              | sbd346v9424_way0_we 
                              | sbd346v9425_way0_we 
                              | sbd346v9426_way0_we 
                              | sbd346v9427_way0_we 
                              | sbd346v9428_way0_we 
                              | sbd346v9429_way0_we 
                              | sbd346v9430_way0_we 
                              | sbd346v9431_way0_we 
                              | sbd346v9432_way0_we 
                              | sbd346v9433_way0_we 
                              | sbd346v9434_way0_we 
                              | sbd346v9435_way0_we 
                              | sbd346v9436_way0_we 
                              | sbd346v9437_way0_we 
                              | sbd346v9438_way0_we 
                              | sbd346v9439_way0_we 
                              | sbd346v9440_way0_we 
                              | sbd346v9441_way0_we 
                              | sbd346v9442_way0_we 
                              | sbd346v9443_way0_we 
                              | sbd346v9444_way0_we 
                              | sbd346v9445_way0_we 
                              | sbd346v9446_way0_we 
                              | sbd346v9447_way0_we 
                              | sbd346v9448_way0_we 
                              | sbd346v9449_way0_we 
                              | sbd346v9450_way0_we 
                              | sbd346v9451_way0_we 
                              | sbd346v9452_way0_we 
                              | sbd346v9453_way0_we 
                              | sbd346v9454_way0_we 
                              | sbd346v9455_way0_we 
                              | sbd346v9456_way0_we 
                              | sbd346v9457_way0_we 
                              | sbd346v9458_way0_we 
                              | sbd346v9459_way0_we 
                              | sbd346v9460_way0_we 
                              | sbd346v9461_way0_we 
                              | sbd346v9462_way0_we 
                              | sbd346v9463_way0_we 
                              ;

  wire vx9vkec2yijlr_jhrjx54o = 1'b0
                              | sbd346v940_way1_we
                              | sbd346v941_way1_we
                              | sbd346v942_way1_we
                              | sbd346v943_way1_we
                              | sbd346v944_way1_we
                              | sbd346v945_way1_we
                              | sbd346v946_way1_we
                              | sbd346v947_way1_we
                              | sbd346v948_way1_we
                              | sbd346v949_way1_we
                              | sbd346v9410_way1_we
                              | sbd346v9411_way1_we
                              | sbd346v9412_way1_we
                              | sbd346v9413_way1_we
                              | sbd346v9414_way1_we
                              | sbd346v9415_way1_we
                              | sbd346v9416_way1_we
                              | sbd346v9417_way1_we
                              | sbd346v9418_way1_we
                              | sbd346v9419_way1_we
                              | sbd346v9420_way1_we
                              | sbd346v9421_way1_we
                              | sbd346v9422_way1_we
                              | sbd346v9423_way1_we
                              | sbd346v9424_way1_we
                              | sbd346v9425_way1_we
                              | sbd346v9426_way1_we
                              | sbd346v9427_way1_we
                              | sbd346v9428_way1_we
                              | sbd346v9429_way1_we
                              | sbd346v9430_way1_we
                              | sbd346v9431_way1_we
                              | sbd346v9432_way1_we
                              | sbd346v9433_way1_we
                              | sbd346v9434_way1_we
                              | sbd346v9435_way1_we
                              | sbd346v9436_way1_we
                              | sbd346v9437_way1_we
                              | sbd346v9438_way1_we
                              | sbd346v9439_way1_we
                              | sbd346v9440_way1_we
                              | sbd346v9441_way1_we
                              | sbd346v9442_way1_we
                              | sbd346v9443_way1_we
                              | sbd346v9444_way1_we
                              | sbd346v9445_way1_we
                              | sbd346v9446_way1_we
                              | sbd346v9447_way1_we
                              | sbd346v9448_way1_we
                              | sbd346v9449_way1_we
                              | sbd346v9450_way1_we
                              | sbd346v9451_way1_we
                              | sbd346v9452_way1_we
                              | sbd346v9453_way1_we
                              | sbd346v9454_way1_we
                              | sbd346v9455_way1_we
                              | sbd346v9456_way1_we
                              | sbd346v9457_way1_we
                              | sbd346v9458_way1_we
                              | sbd346v9459_way1_we
                              | sbd346v9460_way1_we
                              | sbd346v9461_way1_we
                              | sbd346v9462_way1_we
                              | sbd346v9463_way1_we
                              ;
  
  wire emd52ti6nwoy8wmgl4ovad4 = wlxoaneirix6ez6fhtyv3os9c3;
  wire ag2lcgnjbjb6qsmz8nyfj8xo = vx9vkec2yijlr_jhrjx54o;


  wire [21-1:0] edzwk0f_72hrauna9np = ({21{ermcr77dq4jhq99jq==2'b00}} & {21{1'b1}})
                                                      | ({21{ermcr77dq4jhq99jq==2'b01}} & {{21- 9{1'b1}},9'b0})
                                                      | ({21{ermcr77dq4jhq99jq==2'b10}} & {{21-18{1'b1}},18'b0})
                                                      ;
                                                      

  wire [21-1:0] xm30ftlghlhimfgyj = a896qcozpsi1ek5tm9[27-1:6] & edzwk0f_72hrauna9np;



  wire [66-1:0] xpjbkfbf63tm66lzrn8iz0av8 = {
                                                                xm30ftlghlhimfgyj,
                                                                kpl3digtonftoyh,
                                                                hnc10arn_rd,
                                                                ermcr77dq4jhq99jq,
                                                                cf1ozmszcxohbmdmqv,
                                                                n9qmjt3s04yv75d,
                                                                vv_afyrrunvcjbtl2_,
                                                                oclzmsyeij5bw,
                                                                he47fcvawyr15g,
                                                                o44hlt5z77imds2,
                                                                mnac5hr2jmri8kx5xj
                                                              };

  wire [66-1:0] pzqax8ejy4hhndogcybi3a2sbceey = xpjbkfbf63tm66lzrn8iz0av8;
  
  
  wire [27-1:0] l63cfn2f2u8kf9sq7q4qroet3p = ({27{ermcr77dq4jhq99jq==2'b00}} & {27{1'b1}})
                                                      | ({27{ermcr77dq4jhq99jq==2'b01}} & {{27- 9{1'b1}}, 9'b0})
                                                      | ({27{ermcr77dq4jhq99jq==2'b10}} & {{27-18{1'b1}},18'b0})
                                                      ;
  wire [27-1:0] znuclykv4zmtqom7of8 = a896qcozpsi1ek5tm9 & l63cfn2f2u8kf9sq7q4qroet3p;

  wire [55-1:0] ys_6ym9zhq2nap8h6ic458 = {
                                                           znuclykv4zmtqom7of8, 
                                                           kpl3digtonftoyh,
                                                           ermcr77dq4jhq99jq,
                                                           n9qmjt3s04yv75d,
                                                           vv_afyrrunvcjbtl2_,
                                                           oclzmsyeij5bw,
                                                           he47fcvawyr15g,
                                                           o44hlt5z77imds2,
                                                           rxosbn3wj_1o6y20fv
                                                          };
  wire m8duke1scmp1j1b2gsxvd0kgwnth = 1'b1;
 
  wire [51-1:0] wb830emeqn9cg6xwqf8zyhmh = {
                                                           znuclykv4zmtqom7of8, 
                                                           kpl3digtonftoyh,
                                                           ermcr77dq4jhq99jq,
                                                           n9qmjt3s04yv75d,
                                                           rxosbn3wj_1o6y20fv
                                                          };
  wire we8bfdl7knt4u7tz_5j3yzk05za = 1'b1;

  wire bfq086wwiq2gcn35xu5ht_ = 1'b0;
  wire oq5a7kel6r6mfb94lmoku6mf2h = 1'b0;



  
  
  
  
  
  
  wire [55-1:0] d0cnik_anppky6tr4eq1_qh = 55'b0;
  wire fw07acfs_f933fiuzbzm_uos808p = 1'b0;

  wire [51-1:0] is3iuu91tdb5m94kq0ge = 51'b0;
  wire w22ftvp0b0wgmzsk047gs8psps58 = 1'b0;

  wire jf57e9ustr_m76k657bv7 = kbv_rf0mvydplzwef_3qe;
  wire o8bdntgotaqjaspa3fho6mx = w90yio82brq3k1uvzp57esy;


  
  
  
  
  
  
  
  wire z_k8w9px8ti01nrstqg8yja = or2jrhp2d5b1798bveca | ~mou2g2qz02878jxn;
  wire bwdihfhlm6ihh6wog_nncy = llqi__ojtcawwmml0 | ~mou2g2qz02878jxn;
  wire n36u23svjuwuqbrgjd7qus75 = uzgdmfu0z6qg2vr_d363mx0v3z16vc | ~yyz7lhabpe7x17h10y;
  wire dn4bjqivrjkkhpghd8r7x = xmusnbfgqnhl529_izdr6u5tv7ky | ~yyz7lhabpe7x17h10y;
  wire mvpexggyuu3q6okq1yf = z_k8w9px8ti01nrstqg8yja & n36u23svjuwuqbrgjd7qus75 & fivfh22sha8ppz[0];
  wire wzxfgymeeysdv9udmue = bwdihfhlm6ihh6wog_nncy & dn4bjqivrjkkhpghd8r7x & fivfh22sha8ppz[0];
  
  wire [6-1:0] gpcz4u7cii_qx2l3i64u2 = r3ud3glj937o4_;

  wire yv9y07j2gpf7td3hfhgk = ~fivfh22sha8ppz[0] | mvpexggyuu3q6okq1yf;
  wire h9rupeicwkhuuc_x9eyb = ~fivfh22sha8ppz[0] | wzxfgymeeysdv9udmue;
  wire m3vodq8e1ip22ea7d1hai =  fivfh22sha8ppz[0] & mvpexggyuu3q6okq1yf; 
  wire cogh1_67zoyj0e2v8hc8v =  fivfh22sha8ppz[0] & wzxfgymeeysdv9udmue; 
  wire [66-1:0] w_601ovw98i6s0w18dv24ta = 66'b0;
  wire [66-1:0] axhnownqpdcqm5zr0ljulot5oy = 66'b0;
  wire [6-1:0] bsfw1fpvv_iu7y6s5 = gpcz4u7cii_qx2l3i64u2;
  
  
  
  
  
  
  
  
  wire jrzwzcl1o4z7nm4lb2yv3 = ~fivfh22sha8ppz[0] | mvpexggyuu3q6okq1yf;
  wire pfbcvnfs6begexbt4_3wvz94_p = ~fivfh22sha8ppz[0] | wzxfgymeeysdv9udmue;
  wire a0exoan5hqn8q_xewop53c9 =  fivfh22sha8ppz[0] & mvpexggyuu3q6okq1yf;
  wire yyyy2iexny5ic6ctfgkbx =  fivfh22sha8ppz[0] & wzxfgymeeysdv9udmue;

  wire [66-1:0] wk6bks3mhazo5109xz1bmw8azl = 66'b0;
  wire [66-1:0] wsyep6576x493nhte6s9ngpc7zhw = 66'b0;
  wire [6-1:0] eb0xcpdsbwzz7dupo25i = fivfh22sha8ppz[6:1];


  
  
  
  
  
  wire wrr04r1umk6gubhknku7tpnb = 1'b1;
  wire k61j2i07_d9mxzb07jemhp7y = 1'b1;
  wire n9c9804vurfjx2m_1tolf_y = 1'b1; 
  wire i2sex0vzcri42vw75t6w_hzv = 1'b1;
  wire [66-1:0] zm9ilm420c04hep9p4zg3rppf1 = 66'b0;
  wire [66-1:0] t5c93ylv80oxb9ntphva4_llypo = 66'b0;
  wire [6-1:0] v9jhx3p9v0kkas567a9i = fivfh22sha8ppz[6-1:0];


  
  
  
  
  
  
  wire okduot7qrje6co_;
  wire uhsfi7nuqd3ylu4oc;

  assign okduot7qrje6co_ = vikfdhomdfhf7ewfaitsy_gj & ~uhsfi7nuqd3ylu4oc; 
  assign uhsfi7nuqd3ylu4oc = g_7nc4dw6abcm & pffig1fl4xtnw;
  wire r4chpfrvnjvn4kj5 = d3o9i8v1m3g16rvwhai2wh7;
  wire u_1dmhhp0oj7r18 = qhcnhctsg82wxcyhu80cuex4c;
  wire sgws6jzons2h3tlui = oadttvx13julmicav817mtk5jev;
  assign hj0v28frzjss37 = (f_yktlpn8eslyt9akam & ~vy13vm0dqfvofi_2dp09) | (lf2bvnvn_k5yqtn5od & ~klkyy__rhf1ui9omvg);
  ux607_gnrl_dffr #(1) zl7yjvjz6b4kzry1o385 (hj0v28frzjss37, e2vq9uu_okytxq, gf33atgy, ru_wi);

  

  assign f_yktlpn8eslyt9akam = okduot7qrje6co_ & ec9ae2r_4n0dqq8xd73im
                         | uhsfi7nuqd3ylu4oc & emd52ti6nwoy8wmgl4ovad4
                         | r4chpfrvnjvn4kj5 & yv9y07j2gpf7td3hfhgk
                         | u_1dmhhp0oj7r18 & jrzwzcl1o4z7nm4lb2yv3
                         | sgws6jzons2h3tlui & wrr04r1umk6gubhknku7tpnb
                         ;
 
  assign lf2bvnvn_k5yqtn5od = okduot7qrje6co_ & warib_3d5o1png93gezjz2
                         | uhsfi7nuqd3ylu4oc & ag2lcgnjbjb6qsmz8nyfj8xo
                         | r4chpfrvnjvn4kj5 & h9rupeicwkhuuc_x9eyb
                         | u_1dmhhp0oj7r18 & pfbcvnfs6begexbt4_3wvz94_p
                         | sgws6jzons2h3tlui & k61j2i07_d9mxzb07jemhp7y
                         ;

  assign vy13vm0dqfvofi_2dp09 = okduot7qrje6co_ & ruuziixs92g5sudfr9ki
                         | uhsfi7nuqd3ylu4oc & wlxoaneirix6ez6fhtyv3os9c3
                         | r4chpfrvnjvn4kj5 & m3vodq8e1ip22ea7d1hai
                         | u_1dmhhp0oj7r18 & a0exoan5hqn8q_xewop53c9
                         | sgws6jzons2h3tlui & n9c9804vurfjx2m_1tolf_y
                         ;

  
  assign klkyy__rhf1ui9omvg = okduot7qrje6co_ & x197sqagslv9avl082ww
                         | uhsfi7nuqd3ylu4oc & vx9vkec2yijlr_jhrjx54o
                         | r4chpfrvnjvn4kj5 & cogh1_67zoyj0e2v8hc8v
                         | u_1dmhhp0oj7r18 & yyyy2iexny5ic6ctfgkbx
                         | sgws6jzons2h3tlui & i2sex0vzcri42vw75t6w_hzv
                         ;
  

  assign  wqhbmg7dvocz1j9wy9 = ({66{okduot7qrje6co_}} & ztixdkyplyl9m0b51_c0qha    )
                             | ({66{uhsfi7nuqd3ylu4oc}} & xpjbkfbf63tm66lzrn8iz0av8)
                             | ({66{r4chpfrvnjvn4kj5}} & w_601ovw98i6s0w18dv24ta   )
                             | ({66{u_1dmhhp0oj7r18}} & wk6bks3mhazo5109xz1bmw8azl )
                             | ({66{sgws6jzons2h3tlui}} & zm9ilm420c04hep9p4zg3rppf1  )
                             ;
  
  
  assign  tp8gw47qpcwgagtuvei = ({66{okduot7qrje6co_}} & ythnrofnodk8gj5gm0owzh    )
                             | ({66{uhsfi7nuqd3ylu4oc}} & pzqax8ejy4hhndogcybi3a2sbceey)
                             | ({66{r4chpfrvnjvn4kj5}} & axhnownqpdcqm5zr0ljulot5oy   )
                             | ({66{u_1dmhhp0oj7r18}} & wsyep6576x493nhte6s9ngpc7zhw )
                             | ({66{sgws6jzons2h3tlui}} & t5c93ylv80oxb9ntphva4_llypo  )
                             ;
 
  
  assign jw_o9pbzjnqwneo0t = ({6{okduot7qrje6co_}} & qj0rupp44fw6_cqrup1    )
                       | ({6{uhsfi7nuqd3ylu4oc}} & g5cld0_xqbmy2o0oiio_4)
                       | ({6{r4chpfrvnjvn4kj5}} & bsfw1fpvv_iu7y6s5   )
                       | ({6{u_1dmhhp0oj7r18}} & eb0xcpdsbwzz7dupo25i )
                       | ({6{sgws6jzons2h3tlui}} & v9jhx3p9v0kkas567a9i  )
                       ;


  
  
  
  
  
  
  wire qammxfl2w_juh = b7z98rnx88w42eg6952nx8x & ~g_7nc4dw6abcm;  
  wire x52s82zhoyw = fpsdt9vdjcwssz9tezden07r7 & ~g_7nc4dw6abcm;
  wire rg2r09fg5o5 = g_7nc4dw6abcm & j48quvipiuwft;
  wire bmrlssdzm1jp3 = g_7nc4dw6abcm & pffig1fl4xtnw;

  assign w9_jhj6c4a6df_4pxyyb = qammxfl2w_juh & fd08zi5rybh6vf54gwko2 & z3g4qkmuiyg_xfbwf7a2r  
                          | x52s82zhoyw & fd08zi5rybh6vf54gwko2 & yw6x0r1j6uhow9nf5qu1
                          | rg2r09fg5o5 & g2s1v1ri9nldpeph
                          | bmrlssdzm1jp3 & g2s1v1ri9nldpeph
                          ;


  assign oh3gt3hus6shq_f5p7d = ({55{qammxfl2w_juh}} & lmvxjn5zlc78w16q73_ybu47 )
                          | ({55{x52s82zhoyw}} & lj_9z8lqgvo5bet98sorzh)
                          | ({55{rg2r09fg5o5}} & d0cnik_anppky6tr4eq1_qh )
                          | ({55{bmrlssdzm1jp3}} & ys_6ym9zhq2nap8h6ic458)
                          ;


  assign zs5xuhg0c8f60zy_nv1v987v74 = qammxfl2w_juh & fd08zi5rybh6vf54gwko2 & zz2s0dg_zi49zvpaj8tygzbbpi
                                | x52s82zhoyw & fd08zi5rybh6vf54gwko2 & mhu5ty6fyi1g5i40jtfpgkenhfn
                                | rg2r09fg5o5 & g2s1v1ri9nldpeph & fw07acfs_f933fiuzbzm_uos808p
                                | bmrlssdzm1jp3 & g2s1v1ri9nldpeph & m8duke1scmp1j1b2gsxvd0kgwnth
                                ;



  assign ezhgcskig85uffd7xor0c = qammxfl2w_juh & ryl6cvoaujvg6lri3e & be_urjfihso_vqebnp9heqpi
                          | x52s82zhoyw & ryl6cvoaujvg6lri3e & je1s58zp9x4crpu7sd0_c_md2
                          | rg2r09fg5o5 & o6zs2age2tfbqxrs
                          | bmrlssdzm1jp3 & o6zs2age2tfbqxrs
                          ;


  assign tbassexmaytz0vwwh79gt = ({51{qammxfl2w_juh}} & h2zqfgvjbnma19r37rn9s )
                          | ({51{x52s82zhoyw}} & gr7kjbwg55_sgsv87k0z)
                          | ({51{rg2r09fg5o5}} & is3iuu91tdb5m94kq0ge )
                          | ({51{bmrlssdzm1jp3}} & wb830emeqn9cg6xwqf8zyhmh)
                          ;
    

  assign ibq_47zipoy6cbbw2uwa2jy_1o = qammxfl2w_juh & ryl6cvoaujvg6lri3e & ba9aqillrmgw1eh2as1fhaja02rx6
                                | x52s82zhoyw & ryl6cvoaujvg6lri3e & d35npx0cpwxc6siaubaf_mx76i3nbqk
                                | rg2r09fg5o5 & o6zs2age2tfbqxrs & w22ftvp0b0wgmzsk047gs8psps58
                                | bmrlssdzm1jp3 & o6zs2age2tfbqxrs & we8bfdl7knt4u7tz_5j3yzk05za
                                ;
 
  assign nvupfco9fb64lzc1ej = qammxfl2w_juh & m7oe8scer3o7hu_v3ct5xtbe
                           | x52s82zhoyw & vbb4gb1qjbfm7yzd98_7t26
                           | rg2r09fg5o5 & jf57e9ustr_m76k657bv7
                           | bmrlssdzm1jp3 & bfq086wwiq2gcn35xu5ht_
                           ;

  assign hi_bckth818lxu0y4nnr6xzf = qammxfl2w_juh & vudlml4_g7imvjcp1o18uo
                             | x52s82zhoyw & rq1ykv7_2goh27c1eo3u3jyynj62
                             | rg2r09fg5o5 & o8bdntgotaqjaspa3fho6mx
                             | bmrlssdzm1jp3 & oq5a7kel6r6mfb94lmoku6mf2h
                             ;

endmodule






























module sgcljp8bjyetj1gfifd(
  input                                           ru_wi,
  input                                           gf33atgy,


  
  input                                           b0l_kaqp,
  input                                           tlygxd1cs0w,
  input                                           i3o6jvv3t7i,
  input                                           xwd9yye9seo2l,
  input [27-1:0]                    uhegwov_bgw,
  input                                           hhmod6mrlp,

  output                                          ata0drtuuh,
  output                                          se_0n3327r,
  output                                          k9ocj6wlczbbe2,
  output                                          rxosbn3wj_1o6y20fv,
  output                                          w90yio82brq3k1uvzp57esy,
  output                                          kbv_rf0mvydplzwef_3qe,
  output [20-1:0]                     kpl3digtonftoyh,
  output [1:0]                                    ermcr77dq4jhq99jq,
  output                                          mnac5hr2jmri8kx5xj,
  output                                          o44hlt5z77imds2,
  output                                          he47fcvawyr15g,
  output                                          oclzmsyeij5bw,
  output                                          vv_afyrrunvcjbtl2_,
  output                                          n9qmjt3s04yv75d,
  output                                          cf1ozmszcxohbmdmqv,


  
  output [32-1:0]                      fwt3o39z4wp7kgxvw1t,
  output                                          mvs_fsi6kfei3,
  output                                          pctmewhh2f_cwcf5s69,
  output                                          ulxix1i53xn713u9xj7,
  output                                          b5beplnhdi2bmdath3b7,

  input                                          fratob3hz3uz8_es,
  input                                           cpltrra0abys2mc67,


  input                                           wgzv30ij6tqvr1ykebebnmf,

  

  
  output                                          ax9vq1cjvpo685qhrq8y, 
  input                                           e7xoepkekhele1jha9, 
  output [32-1:0]                      qp_qdf85kgmrdv0g,
  output [1:0]                                    dulmf_uxmfqqtg2l,
  output                                          ypi9wk4jnw81_n4nch6,
  output                                          dyakcoiio7g_syixx88j,
  output                                          t0y69cfh1u7o0doo239h,
  output                                          mfpiw_tv_z1eky7kc85o_,
  input                                           s7l5s1wmqz91n6j1gc,
  output                                          yq4iwd6ozbphw48uqdu,
  input                                           ewtcvmi5tj2tjjcu,
  input [64-1:0]                          j8_netqgm7ehavktx6w1_,

  
  input [20-1:0]                      b2ulqcjb,
  input                                           rm1dxjejhq7dh3q5m,
  input [1:0]                                     st2zalpx0uf,
  input                                           ni01kj42oob2x,
  input                                           ah8kjlmvnaxzbi,
  input [1:0]                                     ih7iqx5fe57,

  
  output                                          r4_c53bcpygr5c

);

  localparam zm25xvw0veos8x8r = 3;
  
  wire [zm25xvw0veos8x8r-1:0] uie_swu60u4dfcfjp;
  wire [zm25xvw0veos8x8r-1:0] ehkj2kbe12420;
  wire mgar__kreltg1z76w;
  ux607_gnrl_dfflr #(zm25xvw0veos8x8r) oan760smbfan9qmv28e (mgar__kreltg1z76w, uie_swu60u4dfcfjp, ehkj2kbe12420, gf33atgy, ru_wi);


  localparam jj09e69g9izeh6     = 3'd0;
  localparam gj1cn_xluzljfvpth4l  = 3'd1;
  localparam za5rn0pvbe1ybbwl6f8y1  = 3'd2;
  localparam xmzlx96hi4patqwb1dvvd = 3'd3;
  localparam r9j41ay0icrdol8fhzk   = 3'd4;
  localparam u0bfe54adahta1ques    = 3'd5;
  

  wire [zm25xvw0veos8x8r-1:0] u99tnldu986760c5;
  wire [zm25xvw0veos8x8r-1:0] u_o1hryg6odw8kllden;
  wire [zm25xvw0veos8x8r-1:0] f6f9mxh047a9jnty87ri;
  wire [zm25xvw0veos8x8r-1:0] kquagc_yv6a6gsnk5aq9c1;
  wire [zm25xvw0veos8x8r-1:0] rybupy99nixwcjlvx;
  wire [zm25xvw0veos8x8r-1:0] s67r7tvcckkpgs9;

  wire wfoen161d4r42bkqp34lj;
  wire ogcg7kpm5ntmm5f5pnfxqpb;
  wire c_1t2is39wcxu_gxbmxf_xj;
  wire ybdyo99dw3jffmof74t8vv43aovp;
  wire dq55r5tfg7zc8x9nmmh7wza89;
  wire igbfek2f8xd5vcozwc6mvu;

  wire xbs6xqqdjn8qzdom      = (ehkj2kbe12420 == jj09e69g9izeh6    );
  wire k2qlgxv3oy5ppj8s3res   = (ehkj2kbe12420 == gj1cn_xluzljfvpth4l );
  wire h3wurte832ua3h76gqrp6l   = (ehkj2kbe12420 == za5rn0pvbe1ybbwl6f8y1 );
  wire lr2o95dm_bbktf7tl9hpwh6  = (ehkj2kbe12420 == xmzlx96hi4patqwb1dvvd);
  wire xh3vosowd226kams9y8k    = (ehkj2kbe12420 == r9j41ay0icrdol8fhzk  );
  wire rcmrrfxp3hfd_0ct5     = (ehkj2kbe12420 == u0bfe54adahta1ques   );

  assign mgar__kreltg1z76w = wfoen161d4r42bkqp34lj
                       | ogcg7kpm5ntmm5f5pnfxqpb
                       | c_1t2is39wcxu_gxbmxf_xj
                       | ybdyo99dw3jffmof74t8vv43aovp
                       | dq55r5tfg7zc8x9nmmh7wza89
                       | igbfek2f8xd5vcozwc6mvu
                       ;

  assign uie_swu60u4dfcfjp =  ({zm25xvw0veos8x8r{xbs6xqqdjn8qzdom     }} & u99tnldu986760c5     )
                        | ({zm25xvw0veos8x8r{k2qlgxv3oy5ppj8s3res  }} & u_o1hryg6odw8kllden  )
                        | ({zm25xvw0veos8x8r{h3wurte832ua3h76gqrp6l  }} & f6f9mxh047a9jnty87ri  )
                        | ({zm25xvw0veos8x8r{lr2o95dm_bbktf7tl9hpwh6 }} & kquagc_yv6a6gsnk5aq9c1 )
                        | ({zm25xvw0veos8x8r{xh3vosowd226kams9y8k   }} & rybupy99nixwcjlvx   )
                        | ({zm25xvw0veos8x8r{rcmrrfxp3hfd_0ct5    }} & s67r7tvcckkpgs9    )
                        ;



  wire o32vpum2sraiyu3dl    = (uie_swu60u4dfcfjp == jj09e69g9izeh6    ) & mgar__kreltg1z76w;
  wire p6mp3uoeuxd2dlhqz_4kvko = (uie_swu60u4dfcfjp == gj1cn_xluzljfvpth4l ) & mgar__kreltg1z76w;
  wire yelu0ifm01dok1xkz7i9sfd = (uie_swu60u4dfcfjp == za5rn0pvbe1ybbwl6f8y1 ) & mgar__kreltg1z76w;
  wire ks021sdv42uwjt2a4b7n50qpaf= (uie_swu60u4dfcfjp == xmzlx96hi4patqwb1dvvd) & mgar__kreltg1z76w;
  wire fkeje1miwa0oongga3jsvb2h  = (uie_swu60u4dfcfjp == r9j41ay0icrdol8fhzk  ) & mgar__kreltg1z76w;
  wire ukeqsfnih_s1o_0dk_w8els   = (uie_swu60u4dfcfjp == u0bfe54adahta1ques   ) & mgar__kreltg1z76w;


  assign r4_c53bcpygr5c     = (b0l_kaqp | ehkj2kbe12420 != jj09e69g9izeh6);

  assign ata0drtuuh   = xbs6xqqdjn8qzdom;
  assign se_0n3327r = xh3vosowd226kams9y8k;
  assign k9ocj6wlczbbe2  = rcmrrfxp3hfd_0ct5;
  assign rxosbn3wj_1o6y20fv = xh3vosowd226kams9y8k | rcmrrfxp3hfd_0ct5;

  
  assign wfoen161d4r42bkqp34lj = xbs6xqqdjn8qzdom & b0l_kaqp;
  assign u99tnldu986760c5 = gj1cn_xluzljfvpth4l;


  
  wire ywx9fbvnw_g8no;
  wire mrxv14k2syk5_0eo_prc3491vu2;
  wire gppkfp8cx1th0k6k4aoct3vdgmpav = wgzv30ij6tqvr1ykebebnmf & k2qlgxv3oy5ppj8s3res 
                                                         & ~ywx9fbvnw_g8no 
                                                         & ~mrxv14k2syk5_0eo_prc3491vu2; 
  
  wire bkya4oqgqax9ifdldc0dt = gppkfp8cx1th0k6k4aoct3vdgmpav | mrxv14k2syk5_0eo_prc3491vu2
                             ;
  wire oe46no4c38ljpbrgsdlpi6x7;

  assign ogcg7kpm5ntmm5f5pnfxqpb = k2qlgxv3oy5ppj8s3res;
  assign u_o1hryg6odw8kllden = hhmod6mrlp               ? jj09e69g9izeh6   :
                             bkya4oqgqax9ifdldc0dt       ? u0bfe54adahta1ques  :
                             oe46no4c38ljpbrgsdlpi6x7 ? r9j41ay0icrdol8fhzk :
                                                       za5rn0pvbe1ybbwl6f8y1;


  
  
  assign c_1t2is39wcxu_gxbmxf_xj = h3wurte832ua3h76gqrp6l & e7xoepkekhele1jha9;
  assign f6f9mxh047a9jnty87ri = xmzlx96hi4patqwb1dvvd;

  
  assign ybdyo99dw3jffmof74t8vv43aovp = lr2o95dm_bbktf7tl9hpwh6 & s7l5s1wmqz91n6j1gc;
  assign kquagc_yv6a6gsnk5aq9c1 = ewtcvmi5tj2tjjcu ? u0bfe54adahta1ques : gj1cn_xluzljfvpth4l;

  
  assign dq55r5tfg7zc8x9nmmh7wza89 = xh3vosowd226kams9y8k;
  assign rybupy99nixwcjlvx = b0l_kaqp ? gj1cn_xluzljfvpth4l : jj09e69g9izeh6; 

  
  assign igbfek2f8xd5vcozwc6mvu = rcmrrfxp3hfd_0ct5;
  assign s67r7tvcckkpgs9 = b0l_kaqp ? gj1cn_xluzljfvpth4l : jj09e69g9izeh6;


  
  
  
  
  
  
  wire ds_hd7yxf1ad426t = rxosbn3wj_1o6y20fv & b0l_kaqp;
  wire dkfyb96a0__8f0 = xbs6xqqdjn8qzdom & b0l_kaqp;

  wire dym9qcd2znn = ds_hd7yxf1ad426t | dkfyb96a0__8f0;

  
  
  

  wire i54f9nxqggp;
  wire fg920c5kt2m8 = tlygxd1cs0w;
  ux607_gnrl_dfflr #(1) pzzyechrbnl3joq (dym9qcd2znn, fg920c5kt2m8, i54f9nxqggp, gf33atgy, ru_wi);

  wire omxo8zjmjjw0p7;
  wire pvyko2wa_zf98q9e = i3o6jvv3t7i;
  ux607_gnrl_dfflr #(1) jg7aww06mlevgs97_ (dym9qcd2znn, pvyko2wa_zf98q9e, omxo8zjmjjw0p7, gf33atgy, ru_wi);

  wire u34jf86psbiakk;
  wire gi4_hly49c98avr; 
  wire xfr4nhe4e2osue741d = fratob3hz3uz8_es;
  ux607_gnrl_dfflr #(1) bjbxujs0mdw9qdoxlbd52 (u34jf86psbiakk, xfr4nhe4e2osue741d, gi4_hly49c98avr, gf33atgy, ru_wi);

  wire jhfh0wvubm4_3h_0llx;
  wire vxhxbjkk77spepxprlaqcnw6 = cpltrra0abys2mc67;
  ux607_gnrl_dfflr #(1) v4qxv43qg8qs1m5hne90k9h (dym9qcd2znn, vxhxbjkk77spepxprlaqcnw6, jhfh0wvubm4_3h_0llx, gf33atgy, ru_wi);

  wire [1:0] bnuk7i1r040vc;
  wire [1:0] mbxbkx9ksn0ztox = ih7iqx5fe57;
  ux607_gnrl_dfflr #(2) dgw6nthfddusc7tz (dym9qcd2znn, mbxbkx9ksn0ztox, bnuk7i1r040vc, gf33atgy, ru_wi);

  
  
  

  
  
  
  
  
  
  wire [1:0] z18yn0lrl6e;
  wire dge3eitzkr9uu = dym9qcd2znn | hhmod6mrlp; 
  wire jliarhcopu5fa = k2qlgxv3oy5ppj8s3res;
  wire [1:0] cfcimdv09enqnpb = dge3eitzkr9uu ? 2'b00 : (z18yn0lrl6e + 2'b01);
  wire iefz4bpjaqkhvb = dge3eitzkr9uu | jliarhcopu5fa;
  ux607_gnrl_dfflr #(2) rvvoja_gephu63atj (iefz4bpjaqkhvb, cfcimdv09enqnpb, z18yn0lrl6e, gf33atgy, ru_wi);



  
  
  
  
  
  
  wire [64-1:0] qllx20wfbwc;

  wire [64-1:0] f_ylpq2dt6tqar = qllx20wfbwc;
  wire [64-1:0] uc521p6zdkn7p02dbc22;
  wire whh06cku29tn0bl88w7c;

  wire [32-1:0] m01nkyoco0x75jz9u = qllx20wfbwc[32-1:0];
  wire [32-1:0] oo2x79ep1phizk7pg8;
  assign u34jf86psbiakk = k2qlgxv3oy5ppj8s3res & yelu0ifm01dok1xkz7i9sfd;

  wire [64-1:0] dz609dh6grkaxz4jd1x01 = qllx20wfbwc;
  wire [64-1:0] a42e6owkepqeqvj75skijuo;
  wire m0r9896_0s4rtwdglo = k2qlgxv3oy5ppj8s3res & fkeje1miwa0oongga3jsvb2h;


  wire [64-1:0] t5_17ey3993p1 = {64{whh06cku29tn0bl88w7c   }} & uc521p6zdkn7p02dbc22
                                      | {64{u34jf86psbiakk    }} & {{64-32{1'b0}},oo2x79ep1phizk7pg8}
                                      | {64{m0r9896_0s4rtwdglo}} & a42e6owkepqeqvj75skijuo
                                      ;

  wire cn1e5dcmpmz7a0 = whh06cku29tn0bl88w7c | u34jf86psbiakk | m0r9896_0s4rtwdglo;
  ux607_gnrl_dfflr #(64) os6t7p0w96rr1kgz (cn1e5dcmpmz7a0, t5_17ey3993p1, qllx20wfbwc, gf33atgy, ru_wi);

  wire [32-1:0] edi2fgoz3pny6rbsnbi1z = {32{z18yn0lrl6e == 2'b00}} & {b2ulqcjb, uhegwov_bgw[27-1:27-9], 3'b0}
                                               | {32{z18yn0lrl6e == 2'b01}} & {f_ylpq2dt6tqar[32-3:10], uhegwov_bgw[27-10:27-18], 3'b0}
                                               | {32{z18yn0lrl6e == 2'b10}} & {f_ylpq2dt6tqar[32-3:10], uhegwov_bgw[27-19:27-27], 3'b0}
                                               ;

  assign oo2x79ep1phizk7pg8 = edi2fgoz3pny6rbsnbi1z;

  
  
  
  
  
  
  wire [20-1:0] z1lbprjzso4w54 = f_ylpq2dt6tqar[32-3:10];
  wire [8:0] gq1slg3_z7q5n51ap = f_ylpq2dt6tqar[27:19];
  wire [8:0] x81n9uc9klblsq = f_ylpq2dt6tqar[18:10];
  wire lfmcd_zdpqp7_ = f_ylpq2dt6tqar[7];
  wire q4lqkjxi84 = f_ylpq2dt6tqar[6];
  wire mgobzatsr = f_ylpq2dt6tqar[5];
  wire zvxzy6m6__ = f_ylpq2dt6tqar[4];
  wire gc5uh5lxv1kn = f_ylpq2dt6tqar[3];
  wire gzr4fozal = f_ylpq2dt6tqar[2];
  wire txjq64_4j = f_ylpq2dt6tqar[1];
  wire jzo1k85m8alj9 = f_ylpq2dt6tqar[0];


  wire [1:0] kktbljjy1_bd8ah = rm1dxjejhq7dh3q5m ? st2zalpx0uf : ih7iqx5fe57;
  wire rdvtb5h5mlv3ax = (z18yn0lrl6e == 2'b00);

  assign ywx9fbvnw_g8no = jzo1k85m8alj9 & (txjq64_4j | gc5uh5lxv1kn) & ~rdvtb5h5mlv3ax;
  wire s7rkotljlza1 = jzo1k85m8alj9 & ~gc5uh5lxv1kn & ~txjq64_4j & ~rdvtb5h5mlv3ax;
  wire mhw568w_mjc6bfde0j73 = s7rkotljlza1 & z18yn0lrl6e[1] & z18yn0lrl6e[0]; 
  wire g1u70uo3y6wv8fk5 = jzo1k85m8alj9 & ~txjq64_4j & gzr4fozal & ~rdvtb5h5mlv3ax; 

  wire v1tga2lzktow7mxitu6u6d = mhw568w_mjc6bfde0j73 | g1u70uo3y6wv8fk5;
  wire vsmhcgdm9qjn8xhors1ris355a8e4 = ywx9fbvnw_g8no & ( z18yn0lrl6e == 2'b01 & (|{gq1slg3_z7q5n51ap, x81n9uc9klblsq})  
                                                  |z18yn0lrl6e == 2'b10 & (|x81n9uc9klblsq)  
                                                  );
  
  

  wire kz2cy0ussch7thg = ~rdvtb5h5mlv3ax & ~jzo1k85m8alj9;
  wire e98a3331mp3h7naj7 = ywx9fbvnw_g8no & ~q4lqkjxi84 ;  
  wire bkgicfme_groykm1uaf = ywx9fbvnw_g8no & ~lfmcd_zdpqp7_ & omxo8zjmjjw0p7;
  wire k0goimos2ax_a5e = ywx9fbvnw_g8no & ~txjq64_4j & i54f9nxqggp & ~(gc5uh5lxv1kn & ni01kj42oob2x);
  wire vtl8_2_rkhms90edg5 = ywx9fbvnw_g8no & ~gzr4fozal & omxo8zjmjjw0p7;
  wire jmn7iav7oigeh4bxmyi = ywx9fbvnw_g8no & ~gc5uh5lxv1kn & xwd9yye9seo2l;
  wire m04mpkuzs406yj2 = ywx9fbvnw_g8no & 
                         (
                          zvxzy6m6__ & (kktbljjy1_bd8ah == 2'b01) & ~xwd9yye9seo2l & ~ah8kjlmvnaxzbi
                          | zvxzy6m6__ & (ih7iqx5fe57 == 2'b01) & xwd9yye9seo2l
                          |~zvxzy6m6__ & (ih7iqx5fe57 == 2'b00) & xwd9yye9seo2l 
                          |~zvxzy6m6__ & (kktbljjy1_bd8ah == 2'b00) & ~xwd9yye9seo2l 
                         );


  assign mrxv14k2syk5_0eo_prc3491vu2 = k2qlgxv3oy5ppj8s3res & ( v1tga2lzktow7mxitu6u6d
                                                       | vsmhcgdm9qjn8xhors1ris355a8e4
                                                       | kz2cy0ussch7thg
                                                       | e98a3331mp3h7naj7
                                                       | bkgicfme_groykm1uaf
                                                       | k0goimos2ax_a5e
                                                       | vtl8_2_rkhms90edg5
                                                       | jmn7iav7oigeh4bxmyi
                                                       | m04mpkuzs406yj2 
                                                       );
                                
  

  assign fwt3o39z4wp7kgxvw1t   = edi2fgoz3pny6rbsnbi1z;
  assign mvs_fsi6kfei3     = k2qlgxv3oy5ppj8s3res;
  assign pctmewhh2f_cwcf5s69 = xwd9yye9seo2l;
  assign ulxix1i53xn713u9xj7   = i54f9nxqggp;
  assign b5beplnhdi2bmdath3b7  = omxo8zjmjjw0p7;
  wire [1:0] mmwgkw3juwfizpkr_46tzkf = (z18yn0lrl6e == 2'b01) ? 2'b10: 
                                   (z18yn0lrl6e == 2'b10) ? 2'b01: 
                                                          2'b00; 

  assign oe46no4c38ljpbrgsdlpi6x7 = ywx9fbvnw_g8no & ~bkya4oqgqax9ifdldc0dt; 
  
  wire cccikmxr43gbce3epq;
  wire urn4pvnsvvli7il8do4w9 = s7rkotljlza1 & mgobzatsr;
  wire bvek72xgw236z30786bt5 = dym9qcd2znn;
  wire labdrx2p3xz18ruvoy4te = urn4pvnsvvli7il8do4w9 & ~bvek72xgw236z30786bt5;
  wire sjnhkhpqnw7j1o8z5i6 = urn4pvnsvvli7il8do4w9 | bvek72xgw236z30786bt5;
  ux607_gnrl_dfflr #(1) w3skm5uzgkyd1sd_g41vdv (sjnhkhpqnw7j1o8z5i6, labdrx2p3xz18ruvoy4te, cccikmxr43gbce3epq, gf33atgy, ru_wi);


  localparam szsamxxlhq7zjjenpax9 = 20+2+7;

  
  
  
  wire [20-1:0] evv374je2a154hj = {20{1'b0}}
                                       | {20{z18yn0lrl6e == 2'b01}} & {f_ylpq2dt6tqar[32-3:28], 18'b0}
                                       | {20{z18yn0lrl6e == 2'b10}} & {f_ylpq2dt6tqar[32-3:19], 9'b0}
                                       | {20{z18yn0lrl6e == 2'b11}} & {f_ylpq2dt6tqar[32-3:10]}
                                       ;
  wire [1:0] syjrm2mxj5tb9bhyqkx12 = mmwgkw3juwfizpkr_46tzkf;
  wire ld7y9a38i_     = jzo1k85m8alj9      ;
  wire jb2r6ahdjf     = gc5uh5lxv1kn      ;
  wire nsmyiq9n6ar     = gzr4fozal      ;
  wire t7slufcb     = txjq64_4j      ;
  wire dyd2ogruie     = lfmcd_zdpqp7_      ;
  wire xxmevt09_e     = zvxzy6m6__      ;
  wire daxjzxtqgbmcc     = cccikmxr43gbce3epq | mgobzatsr; 


  assign a42e6owkepqeqvj75skijuo[szsamxxlhq7zjjenpax9-1:0] = { evv374je2a154hj,
                                                      syjrm2mxj5tb9bhyqkx12,
                                                      ld7y9a38i_,
                                                      jb2r6ahdjf,
                                                      nsmyiq9n6ar,
                                                      t7slufcb,
                                                      dyd2ogruie,
                                                      xxmevt09_e,
                                                      daxjzxtqgbmcc
                                                    };
  assign a42e6owkepqeqvj75skijuo[64-1:szsamxxlhq7zjjenpax9] = {64-szsamxxlhq7zjjenpax9{1'b0}};
  


  
  
  
  
  
  

  assign { kpl3digtonftoyh,
           ermcr77dq4jhq99jq,
           mnac5hr2jmri8kx5xj,
           o44hlt5z77imds2,
           he47fcvawyr15g,
           oclzmsyeij5bw,
           vv_afyrrunvcjbtl2_,
           n9qmjt3s04yv75d,
           cf1ozmszcxohbmdmqv } = dz609dh6grkaxz4jd1x01[szsamxxlhq7zjjenpax9-1:0];
  

  
  
  
  
  
  assign ax9vq1cjvpo685qhrq8y = h3wurte832ua3h76gqrp6l;
  assign qp_qdf85kgmrdv0g  = m01nkyoco0x75jz9u;
  assign dulmf_uxmfqqtg2l  = 2'b11;
  assign dyakcoiio7g_syixx88j = (bnuk7i1r040vc == 2'b11);
  assign t0y69cfh1u7o0doo239h = (bnuk7i1r040vc == 2'b01);
  assign mfpiw_tv_z1eky7kc85o_ = jhfh0wvubm4_3h_0llx;
  assign ypi9wk4jnw81_n4nch6    = 1'b0  
                             | gi4_hly49c98avr
                             ;



  
  
  
  
  
  assign yq4iwd6ozbphw48uqdu = lr2o95dm_bbktf7tl9hpwh6;
  assign uc521p6zdkn7p02dbc22 = j8_netqgm7ehavktx6w1_;
  assign whh06cku29tn0bl88w7c = lr2o95dm_bbktf7tl9hpwh6 & s7l5s1wmqz91n6j1gc;
  wire fu0fi0bd7j0nbd30s = lr2o95dm_bbktf7tl9hpwh6 & s7l5s1wmqz91n6j1gc & ewtcvmi5tj2tjjcu;
  

  
  
  
  
  
  
  wire vt1kqrcdzdoo1a1h28v_;
  wire oddmmblr4q85ue4qqlh7 = gppkfp8cx1th0k6k4aoct3vdgmpav | fu0fi0bd7j0nbd30s;
  wire v_r_ekvjgf5f25ztv58gp = dym9qcd2znn | hhmod6mrlp;
  wire ptzq_rxuk6qbkgutd9xt8bm4 = oddmmblr4q85ue4qqlh7 & ~v_r_ekvjgf5f25ztv58gp;
  wire b3agdhne85zo2qobzl63c = oddmmblr4q85ue4qqlh7 | v_r_ekvjgf5f25ztv58gp;
  ux607_gnrl_dfflr #(1) jsno3sy7yo3wm9liwas8yl8 (b3agdhne85zo2qobzl63c, ptzq_rxuk6qbkgutd9xt8bm4, vt1kqrcdzdoo1a1h28v_, gf33atgy, ru_wi);
  assign w90yio82brq3k1uvzp57esy = vt1kqrcdzdoo1a1h28v_;


  wire trdufzx9h1f4miot;
  wire d3gv5fe87lj2n05x_xzane9 = mrxv14k2syk5_0eo_prc3491vu2;
  wire bhtr1bniwer509qtd94vb = dym9qcd2znn | hhmod6mrlp;
  wire u4jlvs82lbjq9cspmuyk = d3gv5fe87lj2n05x_xzane9 & ~bhtr1bniwer509qtd94vb;
  wire vsgcsdjn0s54c2vwpmty = d3gv5fe87lj2n05x_xzane9 | bhtr1bniwer509qtd94vb;
  ux607_gnrl_dfflr #(1) vy9aptf3pt5rsdh83bk2nmk (vsgcsdjn0s54c2vwpmty, u4jlvs82lbjq9cspmuyk, trdufzx9h1f4miot, gf33atgy, ru_wi);
  assign kbv_rf0mvydplzwef_3qe = trdufzx9h1f4miot;


endmodule















































module xnkv2ixv6wqo (
  input                                           ru_wi,
  input                                           gf33atgy,

  input                                           g3ljqli3ukatw2132ssx,
  
  input                                           qhne8m65goz1y091ss8, 
  input [27-1:0]                    z83wiqsi0hgv, 
  input                                           mqi6hv3p07axtj, 
  input [1:0]                                     r6p4z7df65i25fz, 
  output                                          zgpvz622wmbpuyplhsxe2y, 
  output                                          h7x7oqrhyprsd9fpyf7ukcq, 
  output                                          q4u0u5t961_a5u67h7zrv, 
  output [55-1:0]              qn5go609a7uekpxe4, 
  output                                          uxqm4y8nwwoy7a4manunpmrxz2a, 
  output                                          tjdyq2su0gawzvcig32cszgu749r, 
  
  
  input                                           qjkug4xiqzawij13384vr4, 
  input                                           pb3pms28fol8dfr0gr8dkit, 
  input                                           cj92o34fmt9lj4qchqzk6arhow, 
  input [16-1:0]                    qr21q8rwg0cu, 
  input [27-1:0]                    g1400sa7kyme0jubnk7du, 
  output                                          l875nvn0_y6wu72ui7ogut, 
  
  
  input                                           j9xmer7ue4wnuw7ba9gy, 
  input [27-1:0]                    kqjz41lwlrrv, 
  input [1:0]                                     ha7j195sl8e_t5, 
  output                                          t0xxoojg_0iodq0py, 
  output                                          mm9g9a4egd29oz9vvgscmya, 
  output                                          qouo17x2sfmp8hi9d3pto43t1, 
  output [51-1:0]              l5xpteag34o1wqsgx, 
  output                                          g2vry3iwllflk3zzplwitn3eq7gc, 
  output                                          ilj8lhiujxv57r4qqghj0_nntz, 
  
  
  input                                           z1l_kkshyf_56cwmaq2dm, 
  input [16-1:0]                    w7u50np_chxy7wq5n9et_q, 
  input [20-1:0]                      l2dse4sd3runnrb1rcbydauc,  
  input                                           kr1rhzlb5gr_wty1pe392s5oqet, 
  input [1:0]                                     ox2ptuhum_e2aodz8wine6h, 
  input                                           g_qmxgznvfin609fmm97kuc2dm02, 
  input                                           i9oln6xm1pi9dzsd61s1kg4dmo7j, 
  
  input                                           yf_5vs18cke5xg660my, 
  input                                           sneofd4rq3b0m9eu91r8,
  input [8*1-1:0]               d6vb8lyc7vlnm0o3arpqw68r, 
  input [8*1-1:0]               pxmnhz1pxp2i2mmdb6540, 
  input [8*1-1:0]               pfeolrpx0uzt9jq1ndjruu_, 
  input [8*2-1:0]               xa286l0j7185h2h8cym8, 
  input [8*1-1:0]               vs6zhd0u5jdq_fconvsekj, 
  input [8*32-1:0]      n9tjosvoxai4p0sj6mb, 
  

  
  output                                          i0acx70llka5qu09r5jd, 
  output                                          e44u8ctdv_z5u19to, 
  output                                          h7k_k0xxi7vktla, 
  output                                          v_vouzmjecsvtjxt, 
  output [66-1:0]               ef9y8yyld9onuy00de7o, 
  output [66-1:0]               ammhazyeeglt3ewt4p, 
  output [6-1:0]              xvwzwg7_3ek2tx, 
  input  [66-1:0]               y8sg6kbsyavoh4usiqn, 
  input  [66-1:0]               gnqkycbjc0k9k4_edoube, 
  
  
  
  output                                          xib8tki1lzl05e71ry, 
  input                                           hdle8ta5fimb1inf1z, 
  output [32-1:0]                      trtxm7l0l_kp36i9y,
  output [1:0]                                    p0akg_4worvsnfq_q36vp,
  output                                          mqdc73rtez0bzh2_1,
  output                                          oj6rvjf7ujgb34264,
  output                                          vjfz03uzu8p_0jhhvvev,
  output                                          vl5p5iump0rpm1hbr,
  input                                           p1qeemcgwrrzzt73bl,
  output                                          ertspxpg0txqgp9i6fx53,
  input                                           z3xt8rx_qs6z0goo1,
  input [64-1:0]                          ln7r12q36ofpcd6m6u,

  output                                          trtkzwpsx6l

);

  wire                                            kbi8qdl8tmgm5j0uu1p1xu0;
  wire                                            on37whxvtxni09my52drx;
  wire                                            ntychvakx3t8mzzgh8_ev;
  wire [27-1:0]                     k11nc9vg2x3_cg_semdn;
  wire [27-1:0]                     y0__7wpxqx83r42pl;

  wire                                            w9_jhj6c4a6df_4pxyyb;
  wire [55-1:0]                oh3gt3hus6shq_f5p7d;
  wire                                            zs5xuhg0c8f60zy_nv1v987v74;
  
  wire                                            ezhgcskig85uffd7xor0c;
  wire [51-1:0]                tbassexmaytz0vwwh79gt;
  wire                                            ibq_47zipoy6cbbw2uwa2jy_1o;

  wire                                            nvupfco9fb64lzc1ej;
  wire                                            hi_bckth818lxu0y4nnr6xzf;

  wire                                            xhehq_1td3fs;
  wire                                            m0rgjbiqu6nadc33k5;

  wire                                            m01i4z2a2meu;
  wire                                            mou2g2qz02878jxn;
  wire                                            yyz7lhabpe7x17h10y;
  wire [16-1:0]                     j3d84gxpt2b4pd8;
  wire                                            ew6x7412r46;

  wire                                            ata0drtuuh;
  wire                                            k9ocj6wlczbbe2;
  wire                                            se_0n3327r;
  wire                                            rxosbn3wj_1o6y20fv;
  wire                                            w90yio82brq3k1uvzp57esy;
  wire                                            kbv_rf0mvydplzwef_3qe;


  wire [20-1:0]                       kpl3digtonftoyh;
  wire [1:0]                                      ermcr77dq4jhq99jq;
  wire                                            mnac5hr2jmri8kx5xj;
  wire                                            o44hlt5z77imds2;
  wire                                            he47fcvawyr15g;
  wire                                            oclzmsyeij5bw;
  wire                                            vv_afyrrunvcjbtl2_;
  wire                                            n9qmjt3s04yv75d;
  wire                                            cf1ozmszcxohbmdmqv;

  
  wire [27-1:0]                     uhegwov_bgw;
  wire                                            b0l_kaqp;
  wire                                            tlygxd1cs0w;
  wire                                            i3o6jvv3t7i;
  wire                                            xwd9yye9seo2l;

  wire                                            hhmod6mrlp = 1'b0; 

  wire [32-1:0]                        fwt3o39z4wp7kgxvw1t;
  wire                                            mvs_fsi6kfei3;
  wire                                            pctmewhh2f_cwcf5s69;
  wire                                            ulxix1i53xn713u9xj7;
  wire                                            b5beplnhdi2bmdath3b7;
  

  wire                                            wgzv30ij6tqvr1ykebebnmf;

  wire [32-1:0]                        aehmj46c34ed6a0pb0;
  wire                                            zev6d96kah47qb;
  wire                                            cra0dkwdvx0ihnd_xh6rgjlj_9;
  wire                                            ilq7084h434m7cfiznn;
  wire                                            lblyw80ur;
  
  wire                                            uffg2hvo7n434unl4s45oodbr;
  wire                                            im060noyiuihen00u8qh;
  wire                                            p9_d39xvr2hasr1_h1b7;
  wire                                            gyalmuzig9xbui_og;
  wire                                            lxkixcjuqcytzy;
  wire                                            ynkkniwzqhh9y0le;
  wire [32-1:0]                        gkxwt91rch3ir_gn4353q;
  wire                                            qof8e1wj8wm0vj_;

  wire                                            a12zdb8h90f5;

  wire                                            zhvjiiwk09so1foo5i_o9x;
  wire                                            pxtixm9y0620ihre7hd2pu5l;
  wire [32-1:0  ]                      q08dlg0s0csrtgosqa;
  wire [1:0]                                      u5wdh8xtwsdew0fpf5sj8y;
  wire                                            lh4tjxmbn7t8pk6toyz7c;
  wire                                            r0ly0j_gqyee2z0tun10r;
  wire                                            qsh14wsvd8onhwmjnf;
  wire [64-1:0]                           cboj5whx27x6ubhsumzjzqq;

  wire                                            r4_c53bcpygr5c;
  wire                                            d4ab_e8ynn1a53_52a3;

  wire [1:0]                                      s6u3f028i2i9ac9e94l;
  wire [1:0]                                      crlyza4dmh_xv3objkjm;

  n9qdnl9_3k0n2m1yo4pxt j_nvjhyum5d7o_gn_mlk0(
    .ru_wi                  (ru_wi),
    .gf33atgy                    (gf33atgy),

    .g3ljqli3ukatw2132ssx     (g3ljqli3ukatw2132ssx),
    .fkuqlh34r              (z1l_kkshyf_56cwmaq2dm),
    .hnc10arn_rd              (w7u50np_chxy7wq5n9et_q),
    .rm1dxjejhq7dh3q5m           (kr1rhzlb5gr_wty1pe392s5oqet),
    .st2zalpx0uf            (ox2ptuhum_e2aodz8wine6h),
    .ni01kj42oob2x            (g_qmxgznvfin609fmm97kuc2dm02),
    .ah8kjlmvnaxzbi            (i9oln6xm1pi9dzsd61s1kg4dmo7j),
    .toox2fc0snvsr_n           (crlyza4dmh_xv3objkjm),

    .f_yktlpn8eslyt9akam        (i0acx70llka5qu09r5jd),
    .lf2bvnvn_k5yqtn5od        (e44u8ctdv_z5u19to),
    .vy13vm0dqfvofi_2dp09        (h7k_k0xxi7vktla),
    .klkyy__rhf1ui9omvg        (v_vouzmjecsvtjxt),
    .wqhbmg7dvocz1j9wy9     (ef9y8yyld9onuy00de7o),
    .tp8gw47qpcwgagtuvei     (ammhazyeeglt3ewt4p),
    .jw_o9pbzjnqwneo0t          (xvwzwg7_3ek2tx),
    .qbksws8auoc48qp3sb      (y8sg6kbsyavoh4usiqn),
    .xyeddoohku7q6ja9pvnp      (gnqkycbjc0k9k4_edoube),

    .kbi8qdl8tmgm5j0uu1p1xu0     (kbi8qdl8tmgm5j0uu1p1xu0),
    .on37whxvtxni09my52drx      (on37whxvtxni09my52drx),
    .ntychvakx3t8mzzgh8_ev     (ntychvakx3t8mzzgh8_ev),
    .k11nc9vg2x3_cg_semdn        (k11nc9vg2x3_cg_semdn),
    .y0__7wpxqx83r42pl        (y0__7wpxqx83r42pl),

    .w9_jhj6c4a6df_4pxyyb       (w9_jhj6c4a6df_4pxyyb),
    .oh3gt3hus6shq_f5p7d       (oh3gt3hus6shq_f5p7d),
    .zs5xuhg0c8f60zy_nv1v987v74 (zs5xuhg0c8f60zy_nv1v987v74),
    
    .ezhgcskig85uffd7xor0c       (ezhgcskig85uffd7xor0c),
    .tbassexmaytz0vwwh79gt       (tbassexmaytz0vwwh79gt),
    .ibq_47zipoy6cbbw2uwa2jy_1o (ibq_47zipoy6cbbw2uwa2jy_1o),

    .nvupfco9fb64lzc1ej      (nvupfco9fb64lzc1ej),
    .hi_bckth818lxu0y4nnr6xzf    (hi_bckth818lxu0y4nnr6xzf),
    
    .xhehq_1td3fs           (xhehq_1td3fs),
    .m0rgjbiqu6nadc33k5        (m0rgjbiqu6nadc33k5),
    

    .m01i4z2a2meu           (m01i4z2a2meu),
    .mou2g2qz02878jxn        (mou2g2qz02878jxn),
    .yyz7lhabpe7x17h10y      (yyz7lhabpe7x17h10y),
    .j3d84gxpt2b4pd8            (j3d84gxpt2b4pd8),
    .ew6x7412r46            (ew6x7412r46),

    .b3ymasxx4cnt            (ata0drtuuh),
    .j48quvipiuwft           (k9ocj6wlczbbe2),
    .pffig1fl4xtnw          (se_0n3327r),
    .rxosbn3wj_1o6y20fv          (rxosbn3wj_1o6y20fv),
    .w90yio82brq3k1uvzp57esy   (w90yio82brq3k1uvzp57esy),
    .kbv_rf0mvydplzwef_3qe     (kbv_rf0mvydplzwef_3qe),

    .kpl3digtonftoyh            (kpl3digtonftoyh),
    .ermcr77dq4jhq99jq      (ermcr77dq4jhq99jq),
    .mnac5hr2jmri8kx5xj          (mnac5hr2jmri8kx5xj),
    .o44hlt5z77imds2          (o44hlt5z77imds2),
    .he47fcvawyr15g          (he47fcvawyr15g),
    .oclzmsyeij5bw          (oclzmsyeij5bw),
    .vv_afyrrunvcjbtl2_          (vv_afyrrunvcjbtl2_),
    .n9qmjt3s04yv75d          (n9qmjt3s04yv75d),
    .cf1ozmszcxohbmdmqv          (cf1ozmszcxohbmdmqv),

    .uhegwov_bgw                 (uhegwov_bgw),
    .b0l_kaqp                (b0l_kaqp),
    .tlygxd1cs0w               (tlygxd1cs0w),
    .i3o6jvv3t7i              (i3o6jvv3t7i),
    .xwd9yye9seo2l             (xwd9yye9seo2l),
    
    .d4ab_e8ynn1a53_52a3      (d4ab_e8ynn1a53_52a3)


  );


  sgcljp8bjyetj1gfifd kbpt281lapcyhbj4uyv1m0n(
    .ru_wi                  (ru_wi),
    .gf33atgy                    (gf33atgy),


    .b0l_kaqp                (b0l_kaqp),
    .tlygxd1cs0w               (tlygxd1cs0w),
    .i3o6jvv3t7i              (i3o6jvv3t7i),
    .xwd9yye9seo2l             (xwd9yye9seo2l),
    .uhegwov_bgw                 (uhegwov_bgw),
    .hhmod6mrlp              (hhmod6mrlp),

    .ata0drtuuh               (ata0drtuuh),
    .k9ocj6wlczbbe2              (k9ocj6wlczbbe2),
    .se_0n3327r             (se_0n3327r),
    .rxosbn3wj_1o6y20fv          (rxosbn3wj_1o6y20fv),
    .w90yio82brq3k1uvzp57esy   (w90yio82brq3k1uvzp57esy),
    .kbv_rf0mvydplzwef_3qe     (kbv_rf0mvydplzwef_3qe),
    .kpl3digtonftoyh            (kpl3digtonftoyh),
    .ermcr77dq4jhq99jq      (ermcr77dq4jhq99jq),
    .mnac5hr2jmri8kx5xj          (mnac5hr2jmri8kx5xj),
    .o44hlt5z77imds2          (o44hlt5z77imds2),
    .he47fcvawyr15g          (he47fcvawyr15g),
    .oclzmsyeij5bw          (oclzmsyeij5bw),
    .vv_afyrrunvcjbtl2_          (vv_afyrrunvcjbtl2_),
    .n9qmjt3s04yv75d          (n9qmjt3s04yv75d),
    .cf1ozmszcxohbmdmqv          (cf1ozmszcxohbmdmqv),


    .fwt3o39z4wp7kgxvw1t         (fwt3o39z4wp7kgxvw1t),
    .mvs_fsi6kfei3           (mvs_fsi6kfei3),
    .pctmewhh2f_cwcf5s69       (pctmewhh2f_cwcf5s69),
    .ulxix1i53xn713u9xj7         (ulxix1i53xn713u9xj7),
    .b5beplnhdi2bmdath3b7        (b5beplnhdi2bmdath3b7),
    
    .fratob3hz3uz8_es            (lblyw80ur),
    .cpltrra0abys2mc67       (a12zdb8h90f5),
    
    .wgzv30ij6tqvr1ykebebnmf (wgzv30ij6tqvr1ykebebnmf),

    .ax9vq1cjvpo685qhrq8y      (zhvjiiwk09so1foo5i_o9x),
    .e7xoepkekhele1jha9      (pxtixm9y0620ihre7hd2pu5l),
    .qp_qdf85kgmrdv0g       (q08dlg0s0csrtgosqa),
    .dulmf_uxmfqqtg2l       (u5wdh8xtwsdew0fpf5sj8y),
    .ypi9wk4jnw81_n4nch6         (mqdc73rtez0bzh2_1),
    .dyakcoiio7g_syixx88j      (oj6rvjf7ujgb34264),
    .t0y69cfh1u7o0doo239h      (vjfz03uzu8p_0jhhvvev),
    .mfpiw_tv_z1eky7kc85o_      (vl5p5iump0rpm1hbr),
    .s7l5s1wmqz91n6j1gc      (lh4tjxmbn7t8pk6toyz7c),
    .yq4iwd6ozbphw48uqdu      (r0ly0j_gqyee2z0tun10r),
    .ewtcvmi5tj2tjjcu        (qsh14wsvd8onhwmjnf),
    .j8_netqgm7ehavktx6w1_       (cboj5whx27x6ubhsumzjzqq),

    .b2ulqcjb               (l2dse4sd3runnrb1rcbydauc),
    .rm1dxjejhq7dh3q5m           (kr1rhzlb5gr_wty1pe392s5oqet),
    .st2zalpx0uf            (ox2ptuhum_e2aodz8wine6h),
    .ni01kj42oob2x            (g_qmxgznvfin609fmm97kuc2dm02),
    .ah8kjlmvnaxzbi            (i9oln6xm1pi9dzsd61s1kg4dmo7j),
    .ih7iqx5fe57              (s6u3f028i2i9ac9e94l),
    .r4_c53bcpygr5c         (r4_c53bcpygr5c)

  );

   assign xib8tki1lzl05e71ry   = zhvjiiwk09so1foo5i_o9x;
   assign pxtixm9y0620ihre7hd2pu5l = hdle8ta5fimb1inf1z;
   assign trtxm7l0l_kp36i9y    = q08dlg0s0csrtgosqa;
   assign p0akg_4worvsnfq_q36vp    = u5wdh8xtwsdew0fpf5sj8y;
   assign lh4tjxmbn7t8pk6toyz7c = p1qeemcgwrrzzt73bl;
   assign ertspxpg0txqgp9i6fx53   = r0ly0j_gqyee2z0tun10r;
   assign qsh14wsvd8onhwmjnf   = z3xt8rx_qs6z0goo1;
   assign cboj5whx27x6ubhsumzjzqq  = ln7r12q36ofpcd6m6u;

 wire [32-1:0] j8gryhjp7trqw17xi0 = aehmj46c34ed6a0pb0;
  wc2lipjaiimwuy7fx9zp32mr znyaw1u_6z94cmoqfg6bq6y(
    .e98zc_xde8d                 (j8gryhjp7trqw17xi0),
    .lms849k                   (lblyw80ur),
    .dhzk00cwbk               (zev6d96kah47qb)
  );


 wire [32-1:0] ff7r40h7yzdrkij9j = gkxwt91rch3ir_gn4353q;
  d7stl61zflp21cls1tg g_gi1g9jygnc2ow8nwskl4d(
    .sxvvsxtbhyvt             (yf_5vs18cke5xg660my),
    .pcr4upio7_tx37              (n9tjosvoxai4p0sj6mb),
    .uzklqlncpqqm1rav           (d6vb8lyc7vlnm0o3arpqw68r),
    .ortueunvnkx_l5m_j           (pxmnhz1pxp2i2mmdb6540),
    .hwuhtb7ucto_utk56           (pfeolrpx0uzt9jq1ndjruu_),
    .i1env2kmns7qvvuuc           (xa286l0j7185h2h8cym8),
    .g3s3vpafvy3i           (vs6zhd0u5jdq_fconvsekj),

    
    .rm1dxjejhq7dh3q5m           (1'b0),
    .xatytj_r0fv14q           (1'b0),
    .u2k4dyp52s_m                (1'b0),
    .bktu0z1mk56                (p9_d39xvr2hasr1_h1b7),
    .oily7                    (1'b1),
    .ly3dor8                    (1'b0),
    .p1m                    (1'b0),
    .e98zc_xde8d                 (ff7r40h7yzdrkij9j),

    .foj6m18                  (qof8e1wj8wm0vj_)
  );


  
  
  wire vqdwf6w8nvntlzotmu41o;
  wire jiv3l9v2dpzhh0hme8edwu = qhne8m65goz1y091ss8;
  wire at1hi4jzjhwc8t7hqw8i0ow98t = (qhne8m65goz1y091ss8 != vqdwf6w8nvntlzotmu41o);
  ux607_gnrl_dfflr #(1) pobs_k5_54hrdwjnp6vx2e716uye2 (at1hi4jzjhwc8t7hqw8i0ow98t, jiv3l9v2dpzhh0hme8edwu, vqdwf6w8nvntlzotmu41o, gf33atgy, ru_wi);

  wire m65gi_yrqy2n2gq1lnt;
  wire k5y2_x7ozp0odhr_ = mqi6hv3p07axtj;
  wire j721gkykckv8t7cu = (m65gi_yrqy2n2gq1lnt != mqi6hv3p07axtj) & qhne8m65goz1y091ss8;
  ux607_gnrl_dfflr #(1) g65imjpgsx8z0hlzijna (j721gkykckv8t7cu, k5y2_x7ozp0odhr_, m65gi_yrqy2n2gq1lnt, gf33atgy, ru_wi);

  wire kbz6obn9xlyv25r8r2famz;
  ux607_gnrl_dffr #(1) i7sb3ihi4hdbze2pa_xo08n21fs (qjkug4xiqzawij13384vr4, kbz6obn9xlyv25r8r2famz, gf33atgy, ru_wi);

  wire tt1b119l__9dfouqco51ej5 = (qhne8m65goz1y091ss8 & (~vqdwf6w8nvntlzotmu41o | zgpvz622wmbpuyplhsxe2y)) | (qjkug4xiqzawij13384vr4 & ~kbz6obn9xlyv25r8r2famz); 

  wire [27-1:0] pkvucbkmjxaxt;
  wire [27-1:0] wevavulyowll8wq = qjkug4xiqzawij13384vr4 ? g1400sa7kyme0jubnk7du : z83wiqsi0hgv;
  wire cyvpjddes0c4jnu = tt1b119l__9dfouqco51ej5; 
  ux607_gnrl_dfflr #(27) ovl1530s74h7dw_o7rxxp (cyvpjddes0c4jnu, wevavulyowll8wq, pkvucbkmjxaxt, gf33atgy, ru_wi);


  
  wire saqaunfb1hccihzq7tm3ppyd;
  wire ie_arn5f3iehr0lw3eki0v5w = j9xmer7ue4wnuw7ba9gy;
  wire p1s14jq1v4_vn29nu03ta9f = (j9xmer7ue4wnuw7ba9gy != saqaunfb1hccihzq7tm3ppyd);
  ux607_gnrl_dfflr #(1) bouuhp5heey61x7zue693p84_ay8m (p1s14jq1v4_vn29nu03ta9f, ie_arn5f3iehr0lw3eki0v5w, saqaunfb1hccihzq7tm3ppyd, gf33atgy, ru_wi);

  wire shrx523ghhwyg4oi80uhpx9z = j9xmer7ue4wnuw7ba9gy & (~saqaunfb1hccihzq7tm3ppyd | t0xxoojg_0iodq0py); 

  wire [27-1:0] e20yfuej9280mxmn;
  wire [27-1:0] eutswaterpfbkszhj7f = kqjz41lwlrrv;
  wire owyvta3gedzdwkkdy5j = shrx523ghhwyg4oi80uhpx9z;
  ux607_gnrl_dfflr #(27) u0s6v06q_oxf5h5_0 (owyvta3gedzdwkkdy5j, eutswaterpfbkszhj7f, e20yfuej9280mxmn, gf33atgy, ru_wi);
  
  assign s6u3f028i2i9ac9e94l    = xhehq_1td3fs    ? r6p4z7df65i25fz : ha7j195sl8e_t5;
  assign crlyza4dmh_xv3objkjm = m0rgjbiqu6nadc33k5 ? r6p4z7df65i25fz : ha7j195sl8e_t5;
  
  assign a12zdb8h90f5        = xhehq_1td3fs    ? sneofd4rq3b0m9eu91r8 : 1'b0; 
  
  
  
  
  
  
  

  
  assign kbi8qdl8tmgm5j0uu1p1xu0 = qhne8m65goz1y091ss8;
  assign on37whxvtxni09my52drx  = mqi6hv3p07axtj;
  assign ntychvakx3t8mzzgh8_ev = j9xmer7ue4wnuw7ba9gy;
  assign k11nc9vg2x3_cg_semdn    = pkvucbkmjxaxt;
  assign y0__7wpxqx83r42pl    = e20yfuej9280mxmn;

  assign m01i4z2a2meu       = qjkug4xiqzawij13384vr4;
  assign mou2g2qz02878jxn    = pb3pms28fol8dfr0gr8dkit;
  assign yyz7lhabpe7x17h10y  = cj92o34fmt9lj4qchqzk6arhow;
  assign j3d84gxpt2b4pd8        = qr21q8rwg0cu;

  assign ilq7084h434m7cfiznn =  zev6d96kah47qb & cra0dkwdvx0ihnd_xh6rgjlj_9;
  assign wgzv30ij6tqvr1ykebebnmf = ilq7084h434m7cfiznn | qof8e1wj8wm0vj_;



  
  
  
  
  

  assign aehmj46c34ed6a0pb0 = fwt3o39z4wp7kgxvw1t;
  assign cra0dkwdvx0ihnd_xh6rgjlj_9 = pctmewhh2f_cwcf5s69;

 
  assign uffg2hvo7n434unl4s45oodbr = (ox2ptuhum_e2aodz8wine6h == 2'b11);
  assign im060noyiuihen00u8qh      = (s6u3f028i2i9ac9e94l == 2'b11);
  assign p9_d39xvr2hasr1_h1b7      = a12zdb8h90f5;
  assign gyalmuzig9xbui_og = ulxix1i53xn713u9xj7;
  assign lxkixcjuqcytzy = b5beplnhdi2bmdath3b7;
  assign ynkkniwzqhh9y0le = pctmewhh2f_cwcf5s69;
  assign gkxwt91rch3ir_gn4353q = aehmj46c34ed6a0pb0;



  
  
  
  
  
  
  assign zgpvz622wmbpuyplhsxe2y          = w9_jhj6c4a6df_4pxyyb;
  assign h7x7oqrhyprsd9fpyf7ukcq         = nvupfco9fb64lzc1ej;
  assign q4u0u5t961_a5u67h7zrv       = hi_bckth818lxu0y4nnr6xzf;
  assign qn5go609a7uekpxe4          = oh3gt3hus6shq_f5p7d;
  assign uxqm4y8nwwoy7a4manunpmrxz2a    = zs5xuhg0c8f60zy_nv1v987v74;
  assign tjdyq2su0gawzvcig32cszgu749r    = zs5xuhg0c8f60zy_nv1v987v74;
  assign l875nvn0_y6wu72ui7ogut        = ew6x7412r46;

  assign t0xxoojg_0iodq0py          = ezhgcskig85uffd7xor0c;
  assign mm9g9a4egd29oz9vvgscmya         = nvupfco9fb64lzc1ej;
  assign qouo17x2sfmp8hi9d3pto43t1       = hi_bckth818lxu0y4nnr6xzf;
  assign l5xpteag34o1wqsgx          = tbassexmaytz0vwwh79gt;
  assign g2vry3iwllflk3zzplwitn3eq7gc    = ibq_47zipoy6cbbw2uwa2jy_1o;
  assign ilj8lhiujxv57r4qqghj0_nntz    = ibq_47zipoy6cbbw2uwa2jy_1o;


  wire mwilep4hzy69z0r                  = r4_c53bcpygr5c | d4ab_e8ynn1a53_52a3;
  wire ei_cr4ztwk5vk; 
  ux607_gnrl_dffr #(1)  q61z_8s3_p6v930_n (mwilep4hzy69z0r, ei_cr4ztwk5vk, gf33atgy, ru_wi);
  assign trtkzwpsx6l                     = mwilep4hzy69z0r | ei_cr4ztwk5vk; 

endmodule





























module gd24zygbbl9zyo7b5kh11q(
  input   gf33atgy,
  input   ru_wi,
  input   vjpwi,
  output  nuyn4ii2ammwp0,
  output  eqgtpngp18n_lvdz,
  input   vekdxlkh3krc8nq2,
  input   pn5bg45cenp8r81fqkq8
);

  reg  k_y41r7s_yex4;

  wire lmw44bcdnncus7 = vjpwi & vekdxlkh3krc8nq2;
  assign eqgtpngp18n_lvdz = vjpwi & (~k_y41r7s_yex4);

  always @(posedge gf33atgy or negedge ru_wi) begin
    if (~ru_wi) begin
      k_y41r7s_yex4 <= 1'h0;
    end else begin
      if (pn5bg45cenp8r81fqkq8) begin
        k_y41r7s_yex4 <= 1'h0;
      end else begin
        if (lmw44bcdnncus7) begin
          k_y41r7s_yex4 <= 1'h1;
        end
      end
    end
  end

  assign nuyn4ii2ammwp0 = k_y41r7s_yex4; 

endmodule



















module kf2la1880s333ws # (
    parameter tzf9ikb5_qqg1y_e = 3,
    parameter cat22hy7y76lujwa2 = 8,
    parameter gymxwkxs0wahkw_0yn7y0u = 3,
                                    
                                    
                                    
                                    
                                    
                                    
    parameter sewtft9yusm1lav = 0  
)(
  input   dk2xhkj77a,
  input   gf33atgy,
  input   ru_wi,

  input                      th06du2c8e2_b7k,
  output                     irjoi8wvo25u209f_5,
  input  [26-1:0]            zvk11dhgg2s67mkq, 
  input                      zxe59xihintdqfy9d, 
  input  [32-1:0]            u4r4b_6kp09q767q,
  
  output                     klkflmsyyf5w7ar,
  input                      wy36iirxspfw56864,
  output [32-1:0]            h7f6k_ims_9p3,

  output                     aaxhz6kul1ot1yaavzv,
  input  [cat22hy7y76lujwa2-1:0]  da_yai4b0c6,
  input  x_cq40qmp6a,
  output ysjo7jpbga9zbsp,
  output qszs2_0t9_mzkmv3
);




localparam hfcds5urpxlqveoo4e = (((cat22hy7y76lujwa2-1)/32) + 1);

 wire h5maomnmovgqtb7    = th06du2c8e2_b7k & irjoi8wvo25u209f_5;
 wire fz_isl8q3blzlbl2zzf = h5maomnmovgqtb7 & (~zxe59xihintdqfy9d); 
 



 wire [cat22hy7y76lujwa2-1:0]  a82oi6zpkqk83n2oipe7;
 wire [cat22hy7y76lujwa2-1:0]  qoi4fkr36973x72kew7;
 wire [cat22hy7y76lujwa2-1:0]  x62v1om841jew61n144hf;
 wire [cat22hy7y76lujwa2-1:0]  p3agy5z87wpvbnlbhd2pd;

 assign aaxhz6kul1ot1yaavzv = (|qoi4fkr36973x72kew7) | th06du2c8e2_b7k | klkflmsyyf5w7ar;

 wire [cat22hy7y76lujwa2-1:0]  f9n2ww4tvkzba2;
 wire [cat22hy7y76lujwa2-1:0]  p8uxid5kkyo7df5k;


 wire k2ncd2i1iim;
 wire [gymxwkxs0wahkw_0yn7y0u-1:0] uv44wf1j65v2 ;
 wire [gymxwkxs0wahkw_0yn7y0u-1:0] uf7de7zpp08vpoty6 ;
 
 wire c6fzou5v7;
 wire [gymxwkxs0wahkw_0yn7y0u-1:0] bnee_q3n ;
 wire [gymxwkxs0wahkw_0yn7y0u-1:0] s0mhddnef29v_gz ;
 

 wire [cat22hy7y76lujwa2-1:0]  ycrua2947m8x_55;
 wire [cat22hy7y76lujwa2-1:0]  j238od4yrv064ch24;
 wire [cat22hy7y76lujwa2-1:0]  s4uzyyk17lonk9k;
 wire [cat22hy7y76lujwa2-1:0]  yt01u8f0y42y;
 wire [hfcds5urpxlqveoo4e*32-1:0] zht4b3od6bzai2;  

 
 wire [hfcds5urpxlqveoo4e-1:0] fantfusosj7k6mrx;
 wire vl6_9ba2i5fx_xhmtfj;
 wire pkefsp2mb5due9eg0;
 

 
 wire oq7f2ib0dpl9z_mae8kc;
 wire bgzc9eqams6teg5;
 wire [tzf9ikb5_qqg1y_e-1:0] sihkmzttdo2b46; 
 wire [tzf9ikb5_qqg1y_e-1:0] z4ngztakowuu_  ; 
 wire gzr345bh_m8fi3bytd;
 wire idzmafdadoa77;
 wire [tzf9ikb5_qqg1y_e-1:0] way393gdsud2z_4dt; 
 wire [tzf9ikb5_qqg1y_e-1:0] wsqdephh3t2_  ; 

 wire [cat22hy7y76lujwa2-1:0]  w6c2akdrlid9avjvlb;
 wire [cat22hy7y76lujwa2-1:0]  ukjgoxolihuosd;
 wire [tzf9ikb5_qqg1y_e-1:0] gzoacqf2vtdijy5 [cat22hy7y76lujwa2-1:0];
 wire [tzf9ikb5_qqg1y_e-1:0] jyddq3a8ly9p [cat22hy7y76lujwa2-1:0];  
 wire [tzf9ikb5_qqg1y_e-1:0] ojtjwtgewqnaz9w1 [cat22hy7y76lujwa2-1:0];  

 wire mnt6z_bia7o8jv25yt8cf2  [512-1:0] ; 
 wire c47kbapo3fucxthlu5uzd  [256-1:0] ; 
 wire x1cdf7ca0olalffgri6auam  [128-1:0] ; 
 wire jeks0uk13f18yrd295nxpbo  [64-1:0]  ; 
 wire drt3ivzqqm_zyfc5ms4blmk  [32-1:0]  ; 
 wire l9s0fv2odn20c3n085b8  [16-1:0]  ; 
 wire vl9cwqm4dvxgfvmhfxjb  [8-1:0]   ; 
 wire djdaznlzdvhirrro3bg5mvs  [4-1:0]   ; 
 wire h5dh32hx4hsm9pjp8k7z  [2-1:0]   ; 
 wire vpsdxay6t9ljxoyw              ; 

 wire [tzf9ikb5_qqg1y_e-1:0] taob615tstphkxxs [1024-1:0] ; 
 wire [tzf9ikb5_qqg1y_e-1:0] cjzyc77dhoop82t  [512-1:0]  ; 
 wire [tzf9ikb5_qqg1y_e-1:0] y5a1pxovhgosn88n7c  [256-1:0]  ; 
 wire [tzf9ikb5_qqg1y_e-1:0] dnl33ng1rj2vi6ja0s8k  [128-1:0]  ; 
 wire [tzf9ikb5_qqg1y_e-1:0] bvs105isqq0g96g8jx0w[128-1:0]  ; 
 wire [tzf9ikb5_qqg1y_e-1:0] s1hhz3yk0pzhjwixzfqx  [64-1:0]   ; 
 wire [tzf9ikb5_qqg1y_e-1:0] ngkgea6_5gf9bvty  [32-1:0]   ; 
 wire [tzf9ikb5_qqg1y_e-1:0] ygvbbw84u2q0jtj9w50  [16-1:0]   ; 
 wire [tzf9ikb5_qqg1y_e-1:0] yp17di68g8f71mkmlk  [8-1:0]    ; 
 wire [tzf9ikb5_qqg1y_e-1:0] rju3my9lv8y3cbnfo  [4-1:0]    ; 
 wire [tzf9ikb5_qqg1y_e-1:0] te1e5seip8x1q777t  [2-1:0]    ; 
 wire [tzf9ikb5_qqg1y_e-1:0] nwtyfej2utyqgylmb               ; 
 wire [tzf9ikb5_qqg1y_e-1:0] a_dpaxoovd9h29hvz6zc             ; 
                                                                         
 wire [gymxwkxs0wahkw_0yn7y0u-1:0] c41xupq5w7388f27ukm [1024-1:0] ; 
 wire [gymxwkxs0wahkw_0yn7y0u-1:0] d7sy37oab43wukk  [512-1:0]  ; 
 wire [gymxwkxs0wahkw_0yn7y0u-1:0] fnh2cmjnh1_hp96  [256-1:0]  ; 
 wire [gymxwkxs0wahkw_0yn7y0u-1:0] qx0fz6gcnv73y_0zp  [128-1:0]  ; 
 wire [gymxwkxs0wahkw_0yn7y0u-1:0] ryv52yptw9dd5mfovnd[128-1:0]  ; 
 wire [gymxwkxs0wahkw_0yn7y0u-1:0] jxa3a8yqpc1jhrki  [64-1:0]   ; 
 wire [gymxwkxs0wahkw_0yn7y0u-1:0] sn2z9v_g4vkwm1bjb  [32-1:0]   ; 
 wire [gymxwkxs0wahkw_0yn7y0u-1:0] ihyj00khkjbc53z  [16-1:0]   ; 
 wire [gymxwkxs0wahkw_0yn7y0u-1:0] skag4ov5g18bfa3i  [8-1:0]    ; 
 wire [gymxwkxs0wahkw_0yn7y0u-1:0] h7ti6hf70p_ygpnajl  [4-1:0]    ; 
 wire [gymxwkxs0wahkw_0yn7y0u-1:0] mhk558i74bszw0z8  [2-1:0]    ; 
 wire [gymxwkxs0wahkw_0yn7y0u-1:0] hzxz7_d7he6               ; 
 wire [gymxwkxs0wahkw_0yn7y0u-1:0] v_51t44hy95z4p2q             ; 

 wire i_422iukgabh4_dkcm [1024-1:0] ; 
 wire ccnqw_x78a8ay54  [512-1:0]  ; 
 wire f13p8x8ox9qsm6y1  [256-1:0]  ; 
 wire fiu0qb12a90ooc  [128-1:0]  ; 
 wire h4bf06qwiscpvvhd6it[128-1:0]  ; 
 wire idq0i_2dyhcoc  [64-1:0]   ; 
 wire nqx5hep9lxcyrql  [32-1:0]   ; 
 wire emy2mk07ej8qf9gk6e  [16-1:0]   ; 
 wire fwnr2gdp6_pibp  [8-1:0]    ; 
 wire wju5k5n9lhgub7qki  [4-1:0]    ; 
 wire tvp2h1cn5o__x  [2-1:0]    ; 
 wire qaglq05v3wynay2               ; 
 wire fouwrienzarllyb2fj             ; 

 
 wire nojmco2vlex76odckhff8  [512-1:0] ; 
 wire v0v4_plwgcip0eli19cj4h  [256-1:0] ; 
 wire b7wpmpcjii__wknsiyk  [128-1:0] ; 
 wire ngnhy7oxdfylctzylt7  [64-1:0]  ; 
 wire ah07i0clghk1utzvu16  [32-1:0]  ; 
 wire rywdk18g2nr2sc0b8ted  [16-1:0]  ; 
 wire ze6ri1l8jxyy7vw76nj34io  [8-1:0]   ; 
 wire wocc028fu283icuysd5g  [4-1:0]   ; 
 wire wqlvfvo8odxv10r2sv  [2-1:0]   ; 
 wire edfyaofcnrbis37co              ; 

 wire [tzf9ikb5_qqg1y_e-1:0] d79e9q763xm3qc2w [1024-1:0] ; 
 wire [tzf9ikb5_qqg1y_e-1:0] sjcqdgwcznwwqgrpc  [512-1:0]  ; 
 wire [tzf9ikb5_qqg1y_e-1:0] lkqnhmlmzjz1bkmcw  [256-1:0]  ; 
 wire [tzf9ikb5_qqg1y_e-1:0] rnhybhgneoipqsg9  [128-1:0]  ; 
 wire [tzf9ikb5_qqg1y_e-1:0] aq1acidhrbz5buewmkqnbi[128-1:0]  ; 
 wire [tzf9ikb5_qqg1y_e-1:0] gera2jf_uijkoww5_y  [64-1:0]   ; 
 wire [tzf9ikb5_qqg1y_e-1:0] ydi_qu5xqtkc83mfteyr  [32-1:0]   ; 
 wire [tzf9ikb5_qqg1y_e-1:0] ca8pwmy0m3o74x6g04ns  [16-1:0]   ; 
 wire [tzf9ikb5_qqg1y_e-1:0] zpqijbukenuthcnz  [8-1:0]    ; 
 wire [tzf9ikb5_qqg1y_e-1:0] jofphxs6hhru826m  [4-1:0]    ; 
 wire [tzf9ikb5_qqg1y_e-1:0] q0aeo4xujtc3994  [2-1:0]    ; 
 wire [tzf9ikb5_qqg1y_e-1:0] a96b5jn_1zoh4r4dl               ; 
 wire [tzf9ikb5_qqg1y_e-1:0] phh1y4aj3l80kp6nzh             ; 
                                                                         
 wire [gymxwkxs0wahkw_0yn7y0u-1:0] hpp0o9m70w_yyawskm4 [1024-1:0] ; 
 wire [gymxwkxs0wahkw_0yn7y0u-1:0] o63o5r4a81d02q  [512-1:0]  ; 
 wire [gymxwkxs0wahkw_0yn7y0u-1:0] pkd63dc3q4g7uq  [256-1:0]  ; 
 wire [gymxwkxs0wahkw_0yn7y0u-1:0] afvbwh_mufmgrqitkv  [128-1:0]  ; 
 wire [gymxwkxs0wahkw_0yn7y0u-1:0] s1ld8kn7xezto9wljz[128-1:0]  ; 
 wire [gymxwkxs0wahkw_0yn7y0u-1:0] kioexjpglrhp8t  [64-1:0]   ; 
 wire [gymxwkxs0wahkw_0yn7y0u-1:0] zbhpz_qu0faflzfu  [32-1:0]   ; 
 wire [gymxwkxs0wahkw_0yn7y0u-1:0] l0_uj2d8l_j_zr  [16-1:0]   ; 
 wire [gymxwkxs0wahkw_0yn7y0u-1:0] e0nof8mn01h_d  [8-1:0]    ; 
 wire [gymxwkxs0wahkw_0yn7y0u-1:0] m_x8lyyazk62n2ukc  [4-1:0]    ; 
 wire [gymxwkxs0wahkw_0yn7y0u-1:0] cohsp6_l2cjuue0  [2-1:0]    ; 
 wire [gymxwkxs0wahkw_0yn7y0u-1:0] wus473noq42               ; 
 wire [gymxwkxs0wahkw_0yn7y0u-1:0] licry2hg31jq4jakm9             ; 

 wire y_kb1j0en14pj5vd [1024-1:0] ; 
 wire nij7ab8cnxi38  [512-1:0]  ; 
 wire kj4e8svtm6gqdr  [256-1:0]  ; 
 wire jof5rwhigzpntt_a  [128-1:0]  ; 
 wire qdmzjcafcd5bb5nd[128-1:0]  ; 
 wire jlbts1peb_9sr  [64-1:0]   ; 
 wire mwn76z37n1w_0q  [32-1:0]   ; 
 wire rjuh1rgifxl4f1epk  [16-1:0]   ; 
 wire vudsnti_nryt5  [8-1:0]    ; 
 wire gdenr1jqhz1pjs8ih  [4-1:0]    ; 
 wire incpiir4oag9ckdn_  [2-1:0]    ; 
 wire l2esmim0kdiv3df               ; 
 wire r6ky4y12q0pg1             ; 

 wire          ih9z547j1im23m4t [hfcds5urpxlqveoo4e-1:0];
 wire          ifhzvsn6_t5yeg0     [hfcds5urpxlqveoo4e-1:0];
 wire [32-1:0] vstsr81jy_a9ecyd     [hfcds5urpxlqveoo4e-1:0];
 wire [32-1:0] rsfbyutx87j       [hfcds5urpxlqveoo4e-1:0];
 wire [32-1:0] db8zucrxnds60se0    [hfcds5urpxlqveoo4e-1:0];
 wire          f0j5gjqjz49gutt84th [hfcds5urpxlqveoo4e-1:0];
 wire          gxcuwj3vrh47     [hfcds5urpxlqveoo4e-1:0];
 wire [32-1:0] tt7q5u7zduz0_6rp     [hfcds5urpxlqveoo4e-1:0];
 wire [32-1:0] ewg_wzpr6f       [hfcds5urpxlqveoo4e-1:0];
 wire [32-1:0] q8mi7ol7is1aa    [hfcds5urpxlqveoo4e-1:0];

 genvar i;
 integer nzd5e;

 generate 

     if(sewtft9yusm1lav == 1) begin: ey9a0xfbof0e8e4n
          ux607_gnrl_dffr #(1) pwpf50qmh_rwhiai9(k2ncd2i1iim , qszs2_0t9_mzkmv3, gf33atgy, ru_wi);
          ux607_gnrl_dffr #(gymxwkxs0wahkw_0yn7y0u) xo8vak3exlixf5lcob0(uv44wf1j65v2 , uf7de7zpp08vpoty6, gf33atgy, ru_wi);
          
     end
     else begin: hm8humg_aww9kg31817h
          assign qszs2_0t9_mzkmv3 = k2ncd2i1iim ;
          assign uf7de7zpp08vpoty6 = uv44wf1j65v2;
          
     end
     if(sewtft9yusm1lav == 1) begin: dgw03buuof8h48_r
          ux607_gnrl_dffr #(1) zctkie7qya_g8wvh4h(c6fzou5v7 , ysjo7jpbga9zbsp, gf33atgy, ru_wi);
          ux607_gnrl_dffr #(gymxwkxs0wahkw_0yn7y0u) j2hsfax1kcte2e8c8(bnee_q3n , s0mhddnef29v_gz, gf33atgy, ru_wi);
          
     end
     else begin: de7gm7n9xkcxpq0gml
          assign ysjo7jpbga9zbsp = c6fzou5v7 ;
          assign s0mhddnef29v_gz = bnee_q3n;
          
     end

     assign p3agy5z87wpvbnlbhd2pd[0] = 1'b0;
     assign a82oi6zpkqk83n2oipe7[0] = 1'b0;
     assign qoi4fkr36973x72kew7   [0] = 1'b0;
     assign x62v1om841jew61n144hf[0] = 1'b0;

     assign ycrua2947m8x_55[0] = 1'b0;
     assign j238od4yrv064ch24[0] = 1'b0;
     assign s4uzyyk17lonk9k[0] = 1'b0;
     assign yt01u8f0y42y[0] = 1'b0;
     assign zht4b3od6bzai2  [0] = 1'b0;

     assign ukjgoxolihuosd[0] = 1'b0;
     assign gzoacqf2vtdijy5[0] = {tzf9ikb5_qqg1y_e{1'b0}};
     assign jyddq3a8ly9p[0]   = {tzf9ikb5_qqg1y_e{1'b0}};
 
     assign ojtjwtgewqnaz9w1[0] = {tzf9ikb5_qqg1y_e{1'b0}};

   for(i=1; i<cat22hy7y76lujwa2;i=i+1) begin: f7ve5vb6bqmg5m
       
       
       
     gd24zygbbl9zyo7b5kh11q kjcm5uvixk_7iie (
       
       .gf33atgy      (dk2xhkj77a),
       .ru_wi    (ru_wi),
       .vjpwi    (da_yai4b0c6[i]),
       .nuyn4ii2ammwp0    (qoi4fkr36973x72kew7[i]),
       .eqgtpngp18n_lvdz   (a82oi6zpkqk83n2oipe7[i]),
       .vekdxlkh3krc8nq2   (x62v1om841jew61n144hf[i]),
       .pn5bg45cenp8r81fqkq8(p8uxid5kkyo7df5k[i])
     );

     assign p3agy5z87wpvbnlbhd2pd[i] = a82oi6zpkqk83n2oipe7[i] & x62v1om841jew61n144hf[i];

       
       
       
     
     assign x62v1om841jew61n144hf[i] = (~zht4b3od6bzai2[i]);

        
     assign ycrua2947m8x_55[i] = p3agy5z87wpvbnlbhd2pd[i];
        
        
        
     assign j238od4yrv064ch24[i] = f9n2ww4tvkzba2[i];
     assign s4uzyyk17lonk9k[i] = (ycrua2947m8x_55[i] | j238od4yrv064ch24[i]);
     assign yt01u8f0y42y[i] = (ycrua2947m8x_55[i] | (~j238od4yrv064ch24[i]));

        
     ux607_gnrl_dfflr #(1) k_egyjray93xrto(s4uzyyk17lonk9k[i] , yt01u8f0y42y[i], zht4b3od6bzai2[i], dk2xhkj77a, ru_wi);

       
       
       
       
     assign ukjgoxolihuosd[i] = fz_isl8q3blzlbl2zzf & w6c2akdrlid9avjvlb[i];
     assign gzoacqf2vtdijy5[i] = u4r4b_6kp09q767q[tzf9ikb5_qqg1y_e-1:0];
     ux607_gnrl_dfflr #(tzf9ikb5_qqg1y_e) ihqdw6k_czai7m8z(ukjgoxolihuosd[i] , gzoacqf2vtdijy5[i], jyddq3a8ly9p[i], gf33atgy, ru_wi);
 
       
       
       
     assign ojtjwtgewqnaz9w1[i] = jyddq3a8ly9p[i] & {tzf9ikb5_qqg1y_e{zht4b3od6bzai2[i]}};
   end

   for(i=cat22hy7y76lujwa2; i<(hfcds5urpxlqveoo4e*32);i=i+1) begin: ttcwnr94f3i3
       assign zht4b3od6bzai2[i] = 1'b0;
   end

       
       
       
   for(i=0; i<(hfcds5urpxlqveoo4e);i=i+1) begin: mfh_v76dj45ak
     
     assign ifhzvsn6_t5yeg0[i] = ih9z547j1im23m4t[i] & fz_isl8q3blzlbl2zzf;
     ux607_gnrl_dfflr #(32) syzgda_k0w3s4a60_8(ifhzvsn6_t5yeg0[i], vstsr81jy_a9ecyd[i], rsfbyutx87j[i], gf33atgy, ru_wi);

     if(i == 0)begin: nf1xhk08j1ho
         if(hfcds5urpxlqveoo4e == 1) begin:uerysy5xvf6xfxcqm
            assign vstsr81jy_a9ecyd[i] = {u4r4b_6kp09q767q[cat22hy7y76lujwa2-1:1], 1'b0};
         end
         else begin:c0_gojxwcrsqub4npvu35y
            assign vstsr81jy_a9ecyd[i] = {u4r4b_6kp09q767q[31:1], 1'b0};
         end
     end
     else if((hfcds5urpxlqveoo4e-1) == i) begin:ht7xenld3si8
         if((cat22hy7y76lujwa2%32) == 0) begin:wuzomz93g60fm8tmxy_o
           assign vstsr81jy_a9ecyd[i] = u4r4b_6kp09q767q[31:0];
         end
         else begin:a5qc4uk__rbnll4wxw3grf
           assign vstsr81jy_a9ecyd[i] = u4r4b_6kp09q767q[(cat22hy7y76lujwa2%32)-1:0];
         end
     end
     else begin:vusq6iha_lu8x87
       assign vstsr81jy_a9ecyd[i] = u4r4b_6kp09q767q[31:0];
     end

   end
   for(i=0; i<(hfcds5urpxlqveoo4e);i=i+1) begin: ppn318q29njr62g
     
     assign gxcuwj3vrh47[i] = f0j5gjqjz49gutt84th[i] & fz_isl8q3blzlbl2zzf;
     ux607_gnrl_dfflr #(32) nosoa107bbdsfn(gxcuwj3vrh47[i], tt7q5u7zduz0_6rp[i], ewg_wzpr6f[i], gf33atgy, ru_wi);

     if(i == 0)begin: nf1xhk08j1ho
         if(hfcds5urpxlqveoo4e == 1) begin:uerysy5xvf6xfxcqm
            assign tt7q5u7zduz0_6rp[i] = {u4r4b_6kp09q767q[cat22hy7y76lujwa2-1:1], 1'b0};
         end
         else begin:c0_gojxwcrsqub4npvu35y
            assign tt7q5u7zduz0_6rp[i] = {u4r4b_6kp09q767q[31:1], 1'b0};
         end
     end
     else if((hfcds5urpxlqveoo4e-1) == i) begin:ht7xenld3si8
         if((cat22hy7y76lujwa2%32) == 0) begin:wuzomz93g60fm8tmxy_o
           assign tt7q5u7zduz0_6rp[i] = u4r4b_6kp09q767q[31:0];
         end
         else begin:a5qc4uk__rbnll4wxw3grf
           assign tt7q5u7zduz0_6rp[i] = u4r4b_6kp09q767q[(cat22hy7y76lujwa2%32)-1:0];
         end
     end
     else begin:vusq6iha_lu8x87
       assign tt7q5u7zduz0_6rp[i] = u4r4b_6kp09q767q[31:0];
     end

   end

   
       
       
       
       
   wire xs1z6dglk0h1if0w;
   wire klrmtxecl22oi;
   wire chg36rpc_i821dypx5;
   wire j7egvh62h85nvye0lg;

   wire an53efkcwwxbak7tjca = fz_isl8q3blzlbl2zzf & oq7f2ib0dpl9z_mae8kc;
   wire dgm12u9xzfps2on7uz3 = fz_isl8q3blzlbl2zzf & gzr345bh_m8fi3bytd;

   assign bgzc9eqams6teg5 = an53efkcwwxbak7tjca ; 
                         
                         
                         
                         
   assign idzmafdadoa77 = dgm12u9xzfps2on7uz3 ; 

   

   assign sihkmzttdo2b46 = u4r4b_6kp09q767q[tzf9ikb5_qqg1y_e-1:0];
   
                    
                    
                    
   assign way393gdsud2z_4dt = u4r4b_6kp09q767q[tzf9ikb5_qqg1y_e-1:0];

   ux607_gnrl_dfflr #(tzf9ikb5_qqg1y_e) ho3_ofb4vqzyrzd(bgzc9eqams6teg5 , sihkmzttdo2b46, z4ngztakowuu_, gf33atgy, ru_wi);
   ux607_gnrl_dfflr #(tzf9ikb5_qqg1y_e) snjgmc1z8loxvjgx(idzmafdadoa77 , way393gdsud2z_4dt, wsqdephh3t2_, gf33atgy, ru_wi);

   
   
   
   
   
   
   

   
   
   
   
   
   
   
   
   
   
   



     
     
     
     
     
         
             
             
             
             
             
         assign taob615tstphkxxs[0] = {tzf9ikb5_qqg1y_e{1'b0}};  
         assign c41xupq5w7388f27ukm  [0] = {gymxwkxs0wahkw_0yn7y0u{1'b0}};
         assign i_422iukgabh4_dkcm  [0] = 1'b0;
         assign db8zucrxnds60se0[0][0]  = 1'b0;
         assign d79e9q763xm3qc2w[0] = {tzf9ikb5_qqg1y_e{1'b0}};  
         assign hpp0o9m70w_yyawskm4  [0] = {gymxwkxs0wahkw_0yn7y0u{1'b0}};
         assign y_kb1j0en14pj5vd  [0] = 1'b0;
         assign q8mi7ol7is1aa[0][0]  = 1'b0;
     for(i=1; i<cat22hy7y76lujwa2;i=i+1) begin: gwtmuqg71vqzj20
            
         assign db8zucrxnds60se0[i/32][i%32] = (rsfbyutx87j[i/32][i%32] 
                                         | ((~x_cq40qmp6a) & ewg_wzpr6f[i/32][i%32])
                                         )
                                         ;
        assign q8mi7ol7is1aa[i/32][i%32] = (x_cq40qmp6a & ewg_wzpr6f[i/32][i%32]);
            
         assign taob615tstphkxxs[i] = ojtjwtgewqnaz9w1[i] & {tzf9ikb5_qqg1y_e{db8zucrxnds60se0[i/32][i%32]}};
         assign c41xupq5w7388f27ukm  [i] = i[gymxwkxs0wahkw_0yn7y0u-1:0];
         assign i_422iukgabh4_dkcm  [i] = zht4b3od6bzai2[i] & db8zucrxnds60se0[i/32][i%32];
         assign d79e9q763xm3qc2w[i] = ojtjwtgewqnaz9w1[i] & {tzf9ikb5_qqg1y_e{q8mi7ol7is1aa[i/32][i%32]}};
         assign hpp0o9m70w_yyawskm4  [i] = i[gymxwkxs0wahkw_0yn7y0u-1:0];
         assign y_kb1j0en14pj5vd  [i] = zht4b3od6bzai2[i] & q8mi7ol7is1aa[i/32][i%32];

     end

     for(i=cat22hy7y76lujwa2; i<32*hfcds5urpxlqveoo4e; i=i+1) begin: dbmtbmmhjkv66td4jstzd8i_xcpouil
         assign db8zucrxnds60se0[i/32][i%32] = 1'b0;
         assign q8mi7ol7is1aa[i/32][i%32] = 1'b0;
     end
     for(i=cat22hy7y76lujwa2; i<1024;i=i+1) begin: o1o7cansg6fjuqpt2k1qov97bg
         assign taob615tstphkxxs[i] = {tzf9ikb5_qqg1y_e{1'b0}};  
         assign c41xupq5w7388f27ukm  [i] = {gymxwkxs0wahkw_0yn7y0u{1'b0}};
         assign i_422iukgabh4_dkcm  [i] = 1'b0;
         assign d79e9q763xm3qc2w[i] = {tzf9ikb5_qqg1y_e{1'b0}};  
         assign hpp0o9m70w_yyawskm4  [i] = {gymxwkxs0wahkw_0yn7y0u{1'b0}};
         assign y_kb1j0en14pj5vd  [i] = 1'b0;
     end


         
     for(i=0; i<512;i=i+1) begin: urf7puwurdc7nugl5b
         assign mnt6z_bia7o8jv25yt8cf2[i] = (taob615tstphkxxs[2*i] < taob615tstphkxxs[(2*i)+1]); 
         assign cjzyc77dhoop82t[i] = mnt6z_bia7o8jv25yt8cf2[i] ? taob615tstphkxxs[(2*i)+1] : taob615tstphkxxs[2*i];
         assign d7sy37oab43wukk  [i] = mnt6z_bia7o8jv25yt8cf2[i] ? c41xupq5w7388f27ukm  [(2*i)+1] : c41xupq5w7388f27ukm  [2*i];
         assign ccnqw_x78a8ay54  [i] = mnt6z_bia7o8jv25yt8cf2[i] ? i_422iukgabh4_dkcm  [(2*i)+1] : i_422iukgabh4_dkcm  [2*i];
         assign nojmco2vlex76odckhff8[i] = (d79e9q763xm3qc2w[2*i] < d79e9q763xm3qc2w[(2*i)+1]); 
         assign sjcqdgwcznwwqgrpc[i] = nojmco2vlex76odckhff8[i] ? d79e9q763xm3qc2w[(2*i)+1] : d79e9q763xm3qc2w[2*i];
         assign o63o5r4a81d02q  [i] = nojmco2vlex76odckhff8[i] ? hpp0o9m70w_yyawskm4  [(2*i)+1] : hpp0o9m70w_yyawskm4  [2*i];
         assign nij7ab8cnxi38  [i] = nojmco2vlex76odckhff8[i] ? y_kb1j0en14pj5vd  [(2*i)+1] : y_kb1j0en14pj5vd  [2*i];
     end
         
     for(i=0; i<256;i=i+1) begin: wc3v_g425z367q1mue1
         assign c47kbapo3fucxthlu5uzd[i] = (cjzyc77dhoop82t[2*i] < cjzyc77dhoop82t[(2*i)+1]); 
         assign y5a1pxovhgosn88n7c[i] = c47kbapo3fucxthlu5uzd[i] ? cjzyc77dhoop82t[(2*i)+1] : cjzyc77dhoop82t[2*i];
         assign fnh2cmjnh1_hp96  [i] = c47kbapo3fucxthlu5uzd[i] ? d7sy37oab43wukk  [(2*i)+1] : d7sy37oab43wukk  [2*i];
         assign f13p8x8ox9qsm6y1  [i] = c47kbapo3fucxthlu5uzd[i] ? ccnqw_x78a8ay54  [(2*i)+1] : ccnqw_x78a8ay54  [2*i];
         assign v0v4_plwgcip0eli19cj4h[i] = (sjcqdgwcznwwqgrpc[2*i] < sjcqdgwcznwwqgrpc[(2*i)+1]); 
         assign lkqnhmlmzjz1bkmcw[i] = v0v4_plwgcip0eli19cj4h[i] ? sjcqdgwcznwwqgrpc[(2*i)+1] : sjcqdgwcznwwqgrpc[2*i];
         assign pkd63dc3q4g7uq  [i] = v0v4_plwgcip0eli19cj4h[i] ? o63o5r4a81d02q  [(2*i)+1] : o63o5r4a81d02q  [2*i];
         assign kj4e8svtm6gqdr  [i] = v0v4_plwgcip0eli19cj4h[i] ? nij7ab8cnxi38  [(2*i)+1] : nij7ab8cnxi38  [2*i];
     end
         
     for(i=0; i<128;i=i+1) begin: mqjkd_lrrz3fh3cwm7668y
         assign x1cdf7ca0olalffgri6auam[i] = (y5a1pxovhgosn88n7c[2*i] < y5a1pxovhgosn88n7c[(2*i)+1]); 
         assign dnl33ng1rj2vi6ja0s8k[i] = x1cdf7ca0olalffgri6auam[i] ? y5a1pxovhgosn88n7c[(2*i)+1] : y5a1pxovhgosn88n7c[2*i];
         assign qx0fz6gcnv73y_0zp  [i] = x1cdf7ca0olalffgri6auam[i] ? fnh2cmjnh1_hp96  [(2*i)+1] : fnh2cmjnh1_hp96  [2*i];
         assign fiu0qb12a90ooc  [i] = x1cdf7ca0olalffgri6auam[i] ? f13p8x8ox9qsm6y1  [(2*i)+1] : f13p8x8ox9qsm6y1  [2*i];
         assign b7wpmpcjii__wknsiyk[i] = (lkqnhmlmzjz1bkmcw[2*i] < lkqnhmlmzjz1bkmcw[(2*i)+1]); 
         assign rnhybhgneoipqsg9[i] = b7wpmpcjii__wknsiyk[i] ? lkqnhmlmzjz1bkmcw[(2*i)+1] : lkqnhmlmzjz1bkmcw[2*i];
         assign afvbwh_mufmgrqitkv  [i] = b7wpmpcjii__wknsiyk[i] ? pkd63dc3q4g7uq  [(2*i)+1] : pkd63dc3q4g7uq  [2*i];
         assign jof5rwhigzpntt_a  [i] = b7wpmpcjii__wknsiyk[i] ? kj4e8svtm6gqdr  [(2*i)+1] : kj4e8svtm6gqdr  [2*i];
     end
    for(i=0; i<128;i=i+1) begin: ex6h4y03yg5mumwu0x
    ux607_gnrl_dffr #(tzf9ikb5_qqg1y_e) ouv56pdmpcufxyaagm1360rgpsn24(dnl33ng1rj2vi6ja0s8k[i],bvs105isqq0g96g8jx0w[i],gf33atgy,ru_wi);  
    ux607_gnrl_dffr #(1) ntqkw3lxejo6bmu3g5j1o(fiu0qb12a90ooc[i],h4bf06qwiscpvvhd6it[i],gf33atgy,ru_wi);  
    ux607_gnrl_dffr #(gymxwkxs0wahkw_0yn7y0u) rx8xd53e7pv7993sdudq(qx0fz6gcnv73y_0zp[i],ryv52yptw9dd5mfovnd[i],gf33atgy,ru_wi);  
    ux607_gnrl_dffr #(tzf9ikb5_qqg1y_e) mkc2540wi55eb81c4q8pc_jwmfw(rnhybhgneoipqsg9[i],aq1acidhrbz5buewmkqnbi[i],gf33atgy,ru_wi);  
    ux607_gnrl_dffr #(1) tcqelo0oxpe89vh8n43nsp(jof5rwhigzpntt_a[i],qdmzjcafcd5bb5nd[i],gf33atgy,ru_wi);  
    ux607_gnrl_dffr #(gymxwkxs0wahkw_0yn7y0u) pwctfdyvq5_i35c4ak2vo(afvbwh_mufmgrqitkv[i],s1ld8kn7xezto9wljz[i],gf33atgy,ru_wi);  
    end

         
     for(i=0; i<64;i=i+1) begin: skn1r4f7vtna16hnlfx
         assign jeks0uk13f18yrd295nxpbo[i] = (bvs105isqq0g96g8jx0w[2*i] < bvs105isqq0g96g8jx0w[(2*i)+1]); 
         assign s1hhz3yk0pzhjwixzfqx[i] = jeks0uk13f18yrd295nxpbo[i] ? bvs105isqq0g96g8jx0w[(2*i)+1] : bvs105isqq0g96g8jx0w[2*i];
         assign jxa3a8yqpc1jhrki  [i] = jeks0uk13f18yrd295nxpbo[i] ? ryv52yptw9dd5mfovnd  [(2*i)+1] : ryv52yptw9dd5mfovnd  [2*i];
         assign idq0i_2dyhcoc  [i] = jeks0uk13f18yrd295nxpbo[i] ? h4bf06qwiscpvvhd6it  [(2*i)+1] : h4bf06qwiscpvvhd6it  [2*i];
         assign ngnhy7oxdfylctzylt7[i] = (aq1acidhrbz5buewmkqnbi[2*i] < aq1acidhrbz5buewmkqnbi[(2*i)+1]); 
         assign gera2jf_uijkoww5_y[i] = ngnhy7oxdfylctzylt7[i] ? aq1acidhrbz5buewmkqnbi[(2*i)+1] : aq1acidhrbz5buewmkqnbi[2*i];
         assign kioexjpglrhp8t  [i] = ngnhy7oxdfylctzylt7[i] ? s1ld8kn7xezto9wljz  [(2*i)+1] : s1ld8kn7xezto9wljz  [2*i];
         assign jlbts1peb_9sr  [i] = ngnhy7oxdfylctzylt7[i] ? qdmzjcafcd5bb5nd  [(2*i)+1] : qdmzjcafcd5bb5nd  [2*i];
     end
         
     for(i=0; i<32;i=i+1) begin: xcws65db8uymiaoyop6
         assign drt3ivzqqm_zyfc5ms4blmk[i] = (s1hhz3yk0pzhjwixzfqx[2*i] < s1hhz3yk0pzhjwixzfqx[(2*i)+1]); 
         assign ngkgea6_5gf9bvty[i] = drt3ivzqqm_zyfc5ms4blmk[i] ? s1hhz3yk0pzhjwixzfqx[(2*i)+1] : s1hhz3yk0pzhjwixzfqx[2*i];
         assign sn2z9v_g4vkwm1bjb  [i] = drt3ivzqqm_zyfc5ms4blmk[i] ? jxa3a8yqpc1jhrki  [(2*i)+1] : jxa3a8yqpc1jhrki  [2*i];
         assign nqx5hep9lxcyrql  [i] = drt3ivzqqm_zyfc5ms4blmk[i] ? idq0i_2dyhcoc  [(2*i)+1] : idq0i_2dyhcoc  [2*i];
         assign ah07i0clghk1utzvu16[i] = (gera2jf_uijkoww5_y[2*i] < gera2jf_uijkoww5_y[(2*i)+1]); 
         assign ydi_qu5xqtkc83mfteyr[i] = ah07i0clghk1utzvu16[i] ? gera2jf_uijkoww5_y[(2*i)+1] : gera2jf_uijkoww5_y[2*i];
         assign zbhpz_qu0faflzfu  [i] = ah07i0clghk1utzvu16[i] ? kioexjpglrhp8t  [(2*i)+1] : kioexjpglrhp8t  [2*i];
         assign mwn76z37n1w_0q  [i] = ah07i0clghk1utzvu16[i] ? jlbts1peb_9sr  [(2*i)+1] : jlbts1peb_9sr  [2*i];
     end
         
     for(i=0; i<16;i=i+1) begin: tg8js04ob2c6l_h3uoe9
         assign l9s0fv2odn20c3n085b8[i] = (ngkgea6_5gf9bvty[2*i] < ngkgea6_5gf9bvty[(2*i)+1]); 
         assign ygvbbw84u2q0jtj9w50[i] = l9s0fv2odn20c3n085b8[i] ? ngkgea6_5gf9bvty[(2*i)+1] : ngkgea6_5gf9bvty[2*i];
         assign ihyj00khkjbc53z  [i] = l9s0fv2odn20c3n085b8[i] ? sn2z9v_g4vkwm1bjb  [(2*i)+1] : sn2z9v_g4vkwm1bjb  [2*i];
         assign emy2mk07ej8qf9gk6e  [i] = l9s0fv2odn20c3n085b8[i] ? nqx5hep9lxcyrql  [(2*i)+1] : nqx5hep9lxcyrql  [2*i];
         assign rywdk18g2nr2sc0b8ted[i] = (ydi_qu5xqtkc83mfteyr[2*i] < ydi_qu5xqtkc83mfteyr[(2*i)+1]); 
         assign ca8pwmy0m3o74x6g04ns[i] = rywdk18g2nr2sc0b8ted[i] ? ydi_qu5xqtkc83mfteyr[(2*i)+1] : ydi_qu5xqtkc83mfteyr[2*i];
         assign l0_uj2d8l_j_zr  [i] = rywdk18g2nr2sc0b8ted[i] ? zbhpz_qu0faflzfu  [(2*i)+1] : zbhpz_qu0faflzfu  [2*i];
         assign rjuh1rgifxl4f1epk  [i] = rywdk18g2nr2sc0b8ted[i] ? mwn76z37n1w_0q  [(2*i)+1] : mwn76z37n1w_0q  [2*i];
     end
         
     for(i=0; i<8;i=i+1) begin: re0wlw7suywy3dyogou
         assign vl9cwqm4dvxgfvmhfxjb[i] = (ygvbbw84u2q0jtj9w50[2*i] < ygvbbw84u2q0jtj9w50[(2*i)+1]); 
         assign yp17di68g8f71mkmlk[i] = vl9cwqm4dvxgfvmhfxjb[i] ? ygvbbw84u2q0jtj9w50[(2*i)+1] : ygvbbw84u2q0jtj9w50[2*i];
         assign skag4ov5g18bfa3i  [i] = vl9cwqm4dvxgfvmhfxjb[i] ? ihyj00khkjbc53z  [(2*i)+1] : ihyj00khkjbc53z  [2*i];
         assign fwnr2gdp6_pibp  [i] = vl9cwqm4dvxgfvmhfxjb[i] ? emy2mk07ej8qf9gk6e  [(2*i)+1] : emy2mk07ej8qf9gk6e  [2*i];
         assign ze6ri1l8jxyy7vw76nj34io[i] = (ca8pwmy0m3o74x6g04ns[2*i] < ca8pwmy0m3o74x6g04ns[(2*i)+1]); 
         assign zpqijbukenuthcnz[i] = ze6ri1l8jxyy7vw76nj34io[i] ? ca8pwmy0m3o74x6g04ns[(2*i)+1] : ca8pwmy0m3o74x6g04ns[2*i];
         assign e0nof8mn01h_d  [i] = ze6ri1l8jxyy7vw76nj34io[i] ? l0_uj2d8l_j_zr  [(2*i)+1] : l0_uj2d8l_j_zr  [2*i];
         assign vudsnti_nryt5  [i] = ze6ri1l8jxyy7vw76nj34io[i] ? rjuh1rgifxl4f1epk  [(2*i)+1] : rjuh1rgifxl4f1epk  [2*i];
     end
         
     for(i=0; i<4;i=i+1) begin: psptlzby4f1z2uux_h
         assign djdaznlzdvhirrro3bg5mvs[i] = (yp17di68g8f71mkmlk[2*i] < yp17di68g8f71mkmlk[(2*i)+1]); 
         assign rju3my9lv8y3cbnfo[i] = djdaznlzdvhirrro3bg5mvs[i] ? yp17di68g8f71mkmlk[(2*i)+1] : yp17di68g8f71mkmlk[2*i];
         assign h7ti6hf70p_ygpnajl  [i] = djdaznlzdvhirrro3bg5mvs[i] ? skag4ov5g18bfa3i  [(2*i)+1] : skag4ov5g18bfa3i  [2*i];
         assign wju5k5n9lhgub7qki  [i] = djdaznlzdvhirrro3bg5mvs[i] ? fwnr2gdp6_pibp  [(2*i)+1] : fwnr2gdp6_pibp  [2*i];
         assign wocc028fu283icuysd5g[i] = (zpqijbukenuthcnz[2*i] < zpqijbukenuthcnz[(2*i)+1]); 
         assign jofphxs6hhru826m[i] = wocc028fu283icuysd5g[i] ? zpqijbukenuthcnz[(2*i)+1] : zpqijbukenuthcnz[2*i];
         assign m_x8lyyazk62n2ukc  [i] = wocc028fu283icuysd5g[i] ? e0nof8mn01h_d  [(2*i)+1] : e0nof8mn01h_d  [2*i];
         assign gdenr1jqhz1pjs8ih  [i] = wocc028fu283icuysd5g[i] ? vudsnti_nryt5  [(2*i)+1] : vudsnti_nryt5  [2*i];
     end
         
     for(i=0; i<2;i=i+1) begin: ui067tw1gk66engyjixnwg
         assign h5dh32hx4hsm9pjp8k7z[i] = (rju3my9lv8y3cbnfo[2*i] < rju3my9lv8y3cbnfo[(2*i)+1]); 
         assign te1e5seip8x1q777t[i] = h5dh32hx4hsm9pjp8k7z[i] ? rju3my9lv8y3cbnfo[(2*i)+1] : rju3my9lv8y3cbnfo[2*i];
         assign mhk558i74bszw0z8  [i] = h5dh32hx4hsm9pjp8k7z[i] ? h7ti6hf70p_ygpnajl  [(2*i)+1] : h7ti6hf70p_ygpnajl  [2*i];
         assign tvp2h1cn5o__x  [i] = h5dh32hx4hsm9pjp8k7z[i] ? wju5k5n9lhgub7qki  [(2*i)+1] : wju5k5n9lhgub7qki  [2*i];
         assign wqlvfvo8odxv10r2sv[i] = (jofphxs6hhru826m[2*i] < jofphxs6hhru826m[(2*i)+1]); 
         assign q0aeo4xujtc3994[i] = wqlvfvo8odxv10r2sv[i] ? jofphxs6hhru826m[(2*i)+1] : jofphxs6hhru826m[2*i];
         assign cohsp6_l2cjuue0  [i] = wqlvfvo8odxv10r2sv[i] ? m_x8lyyazk62n2ukc  [(2*i)+1] : m_x8lyyazk62n2ukc  [2*i];
         assign incpiir4oag9ckdn_  [i] = wqlvfvo8odxv10r2sv[i] ? gdenr1jqhz1pjs8ih  [(2*i)+1] : gdenr1jqhz1pjs8ih  [2*i];
     end
 endgenerate

     assign vpsdxay6t9ljxoyw = (te1e5seip8x1q777t[0] < te1e5seip8x1q777t[1]); 
     assign nwtyfej2utyqgylmb    = vpsdxay6t9ljxoyw ? te1e5seip8x1q777t[1] : te1e5seip8x1q777t[0];
     assign hzxz7_d7he6      = vpsdxay6t9ljxoyw ? mhk558i74bszw0z8  [1] : mhk558i74bszw0z8  [0];
     assign qaglq05v3wynay2      = vpsdxay6t9ljxoyw ? tvp2h1cn5o__x  [1] : tvp2h1cn5o__x  [0];
     assign edfyaofcnrbis37co = (q0aeo4xujtc3994[0] < q0aeo4xujtc3994[1]); 
     assign a96b5jn_1zoh4r4dl    = edfyaofcnrbis37co ? q0aeo4xujtc3994[1] : q0aeo4xujtc3994[0];
     assign wus473noq42      = edfyaofcnrbis37co ? cohsp6_l2cjuue0  [1] : cohsp6_l2cjuue0  [0];
     assign l2esmim0kdiv3df      = edfyaofcnrbis37co ? incpiir4oag9ckdn_  [1] : incpiir4oag9ckdn_  [0];

    ux607_gnrl_dffr #(tzf9ikb5_qqg1y_e) v4fc2fwwoxcoc3ivcjqqmp(nwtyfej2utyqgylmb,a_dpaxoovd9h29hvz6zc,gf33atgy,ru_wi);  
    ux607_gnrl_dffr #(1) ochpue39eg2lk909rb(qaglq05v3wynay2,fouwrienzarllyb2fj,gf33atgy,ru_wi);  
    ux607_gnrl_dffr #(gymxwkxs0wahkw_0yn7y0u) sdekzmnso6xnza99p(hzxz7_d7he6,v_51t44hy95z4p2q,gf33atgy,ru_wi);  
    ux607_gnrl_dffr #(tzf9ikb5_qqg1y_e) g8dljgvx_mfdn4djxwaaftj(a96b5jn_1zoh4r4dl,phh1y4aj3l80kp6nzh,gf33atgy,ru_wi);  
    ux607_gnrl_dffr #(1) rnlb3xz8cbv3fjlulyr5w(l2esmim0kdiv3df,r6ky4y12q0pg1,gf33atgy,ru_wi);  
    ux607_gnrl_dffr #(gymxwkxs0wahkw_0yn7y0u) upp3ltryzslaetn12q(wus473noq42,licry2hg31jq4jakm9,gf33atgy,ru_wi);  

     assign k2ncd2i1iim           = fouwrienzarllyb2fj & (a_dpaxoovd9h29hvz6zc > z4ngztakowuu_);
     assign uv44wf1j65v2          = v_51t44hy95z4p2q;
     assign c6fzou5v7           = r6ky4y12q0pg1 & (phh1y4aj3l80kp6nzh > wsqdephh3t2_);
     assign bnee_q3n          = licry2hg31jq4jakm9;

   
   
   
   


 
   
    
 generate 
   
         
   
         
         
         
         
    wire [31:0] n061advnk8sndlqu[cat22hy7y76lujwa2-1:0];
    wire [31:0] ur9lzpso4q6_74[hfcds5urpxlqveoo4e-1:0];
    wire [31:0] tdmds3o0p_7r5m[hfcds5urpxlqveoo4e-1:0];
    wire [31:0] lagc5e6e2o465[hfcds5urpxlqveoo4e-1:0];

   for(i=0; i<cat22hy7y76lujwa2;i=i+1) begin: jf0c_8hslf7q1
     assign n061advnk8sndlqu[i] = i*4;
     assign w6c2akdrlid9avjvlb[i] = (zvk11dhgg2s67mkq == $unsigned(n061advnk8sndlqu[i][25:0])); 
   end
   
         
         
         
   for(i=0; i<(hfcds5urpxlqveoo4e);i=i+1) begin: x9ha87h5vniaj
     assign ur9lzpso4q6_74[i] = i*4;
     assign fantfusosj7k6mrx[i] = (zvk11dhgg2s67mkq == ($unsigned(ur9lzpso4q6_74[i][25:0]) + 26'h1000)); 
   end

   
         
         
         
         
     for(i=0; i<(hfcds5urpxlqveoo4e);i=i+1) begin: gt5es1b8emcdp9
       assign tdmds3o0p_7r5m[i] = i*4;
       assign ih9z547j1im23m4t[i] = (zvk11dhgg2s67mkq == ($unsigned(tdmds3o0p_7r5m[i][25:0]) + 26'h2000)); 
     end
   for(i=0; i<(hfcds5urpxlqveoo4e);i=i+1) begin: lg122ts0otkotnsb
       assign lagc5e6e2o465[i] = i*4;
       assign f0j5gjqjz49gutt84th[i] = (zvk11dhgg2s67mkq == ($unsigned(lagc5e6e2o465[i][25:0]) + 26'h2080)); 
   end
   
         
         
         
       assign oq7f2ib0dpl9z_mae8kc = (zvk11dhgg2s67mkq ==  (26'h200000)); 
       assign vl6_9ba2i5fx_xhmtfj = (zvk11dhgg2s67mkq ==  (26'h200004)); 
       assign gzr345bh_m8fi3bytd = (zvk11dhgg2s67mkq ==  (26'h201000)); 
       assign pkefsp2mb5due9eg0 = (zvk11dhgg2s67mkq ==  (26'h201004)); 
       
        
 endgenerate

   
   
   
   
   reg [32-1:0] rgm5uxc7w5_q4yy;
   reg [32-1:0] jqch2dr_p9q8tvl37f;
   reg [32-1:0] l7tz2iqt9co8irq3srw;

   always @* begin:r6ynkpony176lm09iw
       rgm5uxc7w5_q4yy = 32'b0;

       for(nzd5e=0; nzd5e<cat22hy7y76lujwa2;nzd5e=nzd5e+1) begin: jf0c_8hslf7q1
         rgm5uxc7w5_q4yy = rgm5uxc7w5_q4yy | ({32{w6c2akdrlid9avjvlb[nzd5e]}} & jyddq3a8ly9p[nzd5e] );
       end
   end

   always @* begin:s5gdq0fuicnklmb052dg6
       jqch2dr_p9q8tvl37f = 32'b0;

       for(nzd5e=0; nzd5e<(hfcds5urpxlqveoo4e);nzd5e=nzd5e+1) begin: x9ha87h5vniaj
         jqch2dr_p9q8tvl37f = jqch2dr_p9q8tvl37f | ({32{fantfusosj7k6mrx[nzd5e]}} &  
                             {
                                zht4b3od6bzai2[nzd5e*32+31], zht4b3od6bzai2[nzd5e*32+30], zht4b3od6bzai2[nzd5e*32+29], zht4b3od6bzai2[nzd5e*32+28], 
                                zht4b3od6bzai2[nzd5e*32+27], zht4b3od6bzai2[nzd5e*32+26], zht4b3od6bzai2[nzd5e*32+25], zht4b3od6bzai2[nzd5e*32+24], 
                                zht4b3od6bzai2[nzd5e*32+23], zht4b3od6bzai2[nzd5e*32+22], zht4b3od6bzai2[nzd5e*32+21], zht4b3od6bzai2[nzd5e*32+20], 
                                zht4b3od6bzai2[nzd5e*32+19], zht4b3od6bzai2[nzd5e*32+18], zht4b3od6bzai2[nzd5e*32+17], zht4b3od6bzai2[nzd5e*32+16], 
                                zht4b3od6bzai2[nzd5e*32+15], zht4b3od6bzai2[nzd5e*32+14], zht4b3od6bzai2[nzd5e*32+13], zht4b3od6bzai2[nzd5e*32+12], 
                                zht4b3od6bzai2[nzd5e*32+11], zht4b3od6bzai2[nzd5e*32+10], zht4b3od6bzai2[nzd5e*32+09], zht4b3od6bzai2[nzd5e*32+08], 
                                zht4b3od6bzai2[nzd5e*32+07], zht4b3od6bzai2[nzd5e*32+06], zht4b3od6bzai2[nzd5e*32+05], zht4b3od6bzai2[nzd5e*32+04], 
                                zht4b3od6bzai2[nzd5e*32+03], zht4b3od6bzai2[nzd5e*32+02], zht4b3od6bzai2[nzd5e*32+01], zht4b3od6bzai2[nzd5e*32+00]  
                             });
       end
   end

   always @* begin:fsuyegekquivx0tyoz85
       l7tz2iqt9co8irq3srw = 32'b0;

       
       l7tz2iqt9co8irq3srw = l7tz2iqt9co8irq3srw | ({32{oq7f2ib0dpl9z_mae8kc}} & {{32-tzf9ikb5_qqg1y_e  {1'b0}},z4ngztakowuu_}); 
       l7tz2iqt9co8irq3srw = l7tz2iqt9co8irq3srw | ({32{vl6_9ba2i5fx_xhmtfj}} & {{32-gymxwkxs0wahkw_0yn7y0u{1'b0}},uf7de7zpp08vpoty6});
       l7tz2iqt9co8irq3srw = l7tz2iqt9co8irq3srw | ({32{gzr345bh_m8fi3bytd}} & {{32-tzf9ikb5_qqg1y_e  {1'b0}},wsqdephh3t2_}); 
       l7tz2iqt9co8irq3srw = l7tz2iqt9co8irq3srw | ({32{pkefsp2mb5due9eg0}} & {{32-gymxwkxs0wahkw_0yn7y0u{1'b0}},s0mhddnef29v_gz});
       
       for(nzd5e=0; nzd5e<(hfcds5urpxlqveoo4e);nzd5e=nzd5e+1) begin: w8a8p2f05i0cwgloj1
           l7tz2iqt9co8irq3srw = l7tz2iqt9co8irq3srw | ({32{ih9z547j1im23m4t[nzd5e]}} & rsfbyutx87j[nzd5e]);
       end
       for(nzd5e=0; nzd5e<(hfcds5urpxlqveoo4e);nzd5e=nzd5e+1) begin: o256pauxvbijm
           l7tz2iqt9co8irq3srw = l7tz2iqt9co8irq3srw | ({32{f0j5gjqjz49gutt84th[nzd5e]}} & ewg_wzpr6f[nzd5e]);
       end
       
   end

   wire [32-1:0] vf_r9hn9ty7axn = rgm5uxc7w5_q4yy | jqch2dr_p9q8tvl37f | l7tz2iqt9co8irq3srw;


   localparam knhydck6no_65 = 35; 

   wire vpkceiwyiwes_;
   wire k833g5eg4xayl5j66o;
   wire t1pz5o51yu5vuy;
   wire [knhydck6no_65-1:0] iwxu78sftoab_xrp;
   wire [knhydck6no_65-1:0] em0tq6kd5rq9f = {
                                            vf_r9hn9ty7axn,
                                            zxe59xihintdqfy9d,
                                            pkefsp2mb5due9eg0,
                                            vl6_9ba2i5fx_xhmtfj
                                          };

   assign {
           h7f6k_ims_9p3,
           t1pz5o51yu5vuy,
           vpkceiwyiwes_,
           k833g5eg4xayl5j66o
                                    } = iwxu78sftoab_xrp;

        ux607_gnrl_pipe_stage # (
          .CUT_READY(0),
          .DP(1),
          .DW(knhydck6no_65)
        ) cqc6bg2e20t9lh9m3z0ggh (
          .i_vld  (th06du2c8e2_b7k),
          .i_rdy  (irjoi8wvo25u209f_5),
          .i_dat  (em0tq6kd5rq9f),
          .o_vld  (klkflmsyyf5w7ar),
          .o_rdy  (wy36iirxspfw56864),  
          .o_dat  (iwxu78sftoab_xrp),   
        
          .clk  (gf33atgy),
          .rst_n(ru_wi)
        );

   wire   jetszpnn_3n3x0k4d = klkflmsyyf5w7ar & wy36iirxspfw56864;
   wire   wk6gqnfmstzo2w9ixs5 = jetszpnn_3n3x0k4d & t1pz5o51yu5vuy;

   assign xs1z6dglk0h1if0w = k833g5eg4xayl5j66o & wk6gqnfmstzo2w9ixs5;
   assign klrmtxecl22oi = vl6_9ba2i5fx_xhmtfj & fz_isl8q3blzlbl2zzf;
   assign chg36rpc_i821dypx5 = vpkceiwyiwes_ & wk6gqnfmstzo2w9ixs5;
   assign j7egvh62h85nvye0lg = pkefsp2mb5due9eg0 & fz_isl8q3blzlbl2zzf;

   generate 
   
   for(i=0; i<cat22hy7y76lujwa2;i=i+1) begin: wly_cw09ctboc29tlj163

                                       
     assign f9n2ww4tvkzba2[i] = (h7f6k_ims_9p3 == $unsigned(i)) & ((db8zucrxnds60se0[i/32][i%32] & xs1z6dglk0h1if0w) | (q8mi7ol7is1aa[i/32][i%32] & chg36rpc_i821dypx5));
                                       
     assign p8uxid5kkyo7df5k[i] = (u4r4b_6kp09q767q == $unsigned(i)) & ((db8zucrxnds60se0[i/32][i%32] & klrmtxecl22oi) | (q8mi7ol7is1aa[i/32][i%32] & j7egvh62h85nvye0lg));


   end
   endgenerate


endmodule



















module qc2dx_wo71_o92_z4(
  input   dk2xhkj77a ,
  input   gf33atgy,
  input   ru_wi,

  output        b13zu8ysd3u,

  input                      v9ov1b3vn5k4ctkb,
  output                     ub9pjiu4juf6nuqoq2w6,
  input  [32-1:0]            aw0a19a967dn7n0x25w, 
  input                      ogvavqa7ta836s, 
  input  [32-1:0]            sc169gxpr38lpe8,
  input  [ 4-1:0]            hg1g2yh6yktfe_btdst7,
                              
                              
  input                      ty6a2k41y0e9ir8_yzg,
  input                      cwkq4r6_upg_2884r,
  
  output                     dy9ll1o6t6ytby71hf4,
  input                      ow4hbh48f0mt6le4o,
  output [32-1:0]            dek0xt7q6guk2vf6,
  output                     uzwj715coelxmfqs,

  input [32:1] da_yai4b0c6,
  input   x_cq40qmp6a,
  output  ysjo7jpbga9zbsp,
  output  qszs2_0t9_mzkmv3
);

  wire                     klkflmsyyf5w7ar;
  wire                     wy36iirxspfw56864;
  wire [32-1:0]            h7f6k_ims_9p3;

  ux607_gnrl_fifo # (
        .CUT_READY (1),
        .MSKO      (0),
        .DP  (1),
        .DW  (32)
  ) dr57pnc5s_2fzk6x (
        .i_vld(klkflmsyyf5w7ar),
        .i_rdy(wy36iirxspfw56864),
        .i_dat(h7f6k_ims_9p3),
        .o_vld(dy9ll1o6t6ytby71hf4),
        .o_rdy(ow4hbh48f0mt6le4o),  
        .o_dat(dek0xt7q6guk2vf6),  
      
        .clk  (gf33atgy),
        .rst_n(ru_wi)
  );
  wire rmxmly8p_7ju2zn5xm9vbtbukb4h = klkflmsyyf5w7ar & wy36iirxspfw56864;
  wire g1ayxtymznjy9agkm1a8ivxy3ipe = dy9ll1o6t6ytby71hf4 & ow4hbh48f0mt6le4o;

localparam tzf9ikb5_qqg1y_e = 3;
localparam cat22hy7y76lujwa2 = 32+1;
localparam gymxwkxs0wahkw_0yn7y0u = (cat22hy7y76lujwa2<=2)?1:(cat22hy7y76lujwa2<=4)?2:(cat22hy7y76lujwa2<=8)?3:(cat22hy7y76lujwa2<=16)?4:(cat22hy7y76lujwa2<=32)?5:(cat22hy7y76lujwa2<=64)?6:(cat22hy7y76lujwa2<=128)?7:(cat22hy7y76lujwa2<=256)?8:(cat22hy7y76lujwa2<=512)?9:(cat22hy7y76lujwa2<=1024)?10:(cat22hy7y76lujwa2<=2048)?11:(cat22hy7y76lujwa2<=4096)?12:-1;

wire [32:0] fleckfvg71haq0xl8 = {
                  da_yai4b0c6,
                  1'b0 };

wire aaxhz6kul1ot1yaavzv;

kf2la1880s333ws #(
    .tzf9ikb5_qqg1y_e   (tzf9ikb5_qqg1y_e),
    .cat22hy7y76lujwa2      (cat22hy7y76lujwa2),
    .gymxwkxs0wahkw_0yn7y0u (gymxwkxs0wahkw_0yn7y0u),
    .sewtft9yusm1lav   (0) 
) ieqeish335xi51b7(
    .dk2xhkj77a        (dk2xhkj77a        ),      
    .gf33atgy            (gf33atgy),      
    .ru_wi          (ru_wi          ),

    .th06du2c8e2_b7k  (v9ov1b3vn5k4ctkb),
    .irjoi8wvo25u209f_5  (ub9pjiu4juf6nuqoq2w6),
    .zvk11dhgg2s67mkq   (aw0a19a967dn7n0x25w[26-1:0] ),
    .zxe59xihintdqfy9d   (ogvavqa7ta836s ),
    .u4r4b_6kp09q767q  (sc169gxpr38lpe8),
                    
    .klkflmsyyf5w7ar  (klkflmsyyf5w7ar),
    .wy36iirxspfw56864  (wy36iirxspfw56864),
    .h7f6k_ims_9p3  (h7f6k_ims_9p3),

    .aaxhz6kul1ot1yaavzv (aaxhz6kul1ot1yaavzv),

    .da_yai4b0c6 (fleckfvg71haq0xl8),
    .x_cq40qmp6a (x_cq40qmp6a),
    .ysjo7jpbga9zbsp (ysjo7jpbga9zbsp), 
    .qszs2_0t9_mzkmv3 (qszs2_0t9_mzkmv3) 
);

  assign uzwj715coelxmfqs = 1'b0;
  assign b13zu8ysd3u = aaxhz6kul1ot1yaavzv 
                     | g1ayxtymznjy9agkm1a8ivxy3ipe
                     | rmxmly8p_7ju2zn5xm9vbtbukb4h
                     ;


endmodule



















module w3ji4naj4ajyji(
  input           jewtb_k,
  input  [32-2-1:0] wj5ongbu6, 
  output [32-1:0] e0w_why77quoq  
  );


  wire [32-1:0] dws_i84z4ie9lw = {wj5ongbu6, 2'b11}; 

  wire [32-1:0] hsepvqpwkkjmfe32f_zdwd5; 
  wire [32-1:0] zap0dyhammhw6a88_2mm15a = {hsepvqpwkkjmfe32f_zdwd5[32-1-1:0],1'b0}; 

  wire [32-1:0] gyuikqhht8b3aaabz;  

  genvar i;
  generate
    for (i=0; i<32; i=i+1) begin: e4z7n36x1bqp88hk8njp
        if(i==0) begin:xvpcp9wjmb99kn
            assign hsepvqpwkkjmfe32f_zdwd5[0] = 1'b0;
            assign gyuikqhht8b3aaabz[0]   = 1'b0;
        end
        else begin:mltk61kc_oi7ew4w
            assign hsepvqpwkkjmfe32f_zdwd5[i] = (~dws_i84z4ie9lw[i]) & dws_i84z4ie9lw[i-1]; 
            assign gyuikqhht8b3aaabz[i]   = |zap0dyhammhw6a88_2mm15a[i:0];
        end
    end
  endgenerate

  assign e0w_why77quoq = jewtb_k ? {(~({32-2{1'b0}})),2'b00} : gyuikqhht8b3aaabz; 

endmodule



















module d7stl61zflp21cls1tg(

  input sxvvsxtbhyvt,

  input [8*32-1:0] pcr4upio7_tx37, 
  input [8*1-1:0] uzklqlncpqqm1rav,
  input [8*1-1:0] ortueunvnkx_l5m_j,
  input [8*1-1:0] hwuhtb7ucto_utk56,
  input [8*2-1:0] i1env2kmns7qvvuuc,
  input [8*1-1:0] g3s3vpafvy3i,


  input  rm1dxjejhq7dh3q5m,
  input  xatytj_r0fv14q,
  input  u2k4dyp52s_m,
  input  bktu0z1mk56,
  input  oily7,
  input  ly3dor8,
  input  p1m,
  input  [32-1:0] e98zc_xde8d ,
  output foj6m18   
  );


  genvar i;

  wire [32-1:0] wj5ongbu6       [8-1:0]; 
  wire [32-1:0] e0w_why77quoq  [8-1:0];
  wire                  l5dwr36cp4xs      [8-1:0];
  wire                  ievzogco14      [8-1:0];
  wire                  n78fb03bj00v      [8-1:0];
  wire [2-1:0]          zn3av2_qfxg      [8-1:0];
  wire                  alkw6cq4ei      [8-1:0];

  wire  [8-1:0] de9vb1p7mqzggq3c0v4b3  ;
  wire  [8-1:0] cg31jos3lwbosp1uo  ;


  wire  [8-1:0] rbkhedejfse33j8  ;
  wire  [8-1:0] p7icye18y8l6l  ;
  wire  [8-1:0] hlhcnhvw4wjmcl8k_oq;

  wire  [8-1:0] hztrxxh8s9k988m7i ;
  wire  [8-1:0] ab01vsjb5jhs3    ;
  wire  [8-1:0] v4l5fg97ku084rrubqysv;

  generate 
    for (i=0; i<8; i=i+1) begin: kdmkvmzy0w
      assign wj5ongbu6 [i] = pcr4upio7_tx37   [(i*32+32-1) : i*32];
      assign l5dwr36cp4xs[i] = uzklqlncpqqm1rav[(i*1+1-1) : i*1];
      assign ievzogco14[i] = ortueunvnkx_l5m_j[(i*1+1-1) : i*1];
      assign n78fb03bj00v[i] = hwuhtb7ucto_utk56[(i*1+1-1) : i*1];
      assign zn3av2_qfxg[i] = i1env2kmns7qvvuuc[(i*2+2-1) : i*2];
      assign alkw6cq4ei[i] = g3s3vpafvy3i[(i*1+1-1) : i*1];
    end
  endgenerate





  wire fwmbk3wv_1qt = (bktu0z1mk56 ? sxvvsxtbhyvt : 1'b1) & rm1dxjejhq7dh3q5m;

  
  wire jmr5or9glw48yt6 = ( (oily7 | ly3dor8) & fwmbk3wv_1qt) ? xatytj_r0fv14q : (u2k4dyp52s_m | bktu0z1mk56);
  wire z30_md1zf_cg0 = (~jmr5or9glw48yt6);

  generate 
    for (i=0; i<8; i=i+1) begin: g0rwttdjgy4g
      assign rbkhedejfse33j8[i] = (zn3av2_qfxg[i] == 2'b00);
      
      
      assign p7icye18y8l6l[i] = 1'b0;  
      assign hlhcnhvw4wjmcl8k_oq[i] = (zn3av2_qfxg[i] == 2'b11);

      

      w3ji4naj4ajyji p1tra6jm653sl_3cnidz(.jewtb_k(p7icye18y8l6l[i]), .wj5ongbu6(wj5ongbu6[i][32-2-1:0]), .e0w_why77quoq(e0w_why77quoq[i][32-1:0])  );
      
      
      
      
      
      
      
      
      
      
      assign hztrxxh8s9k988m7i[i] = ( (e98zc_xde8d & e0w_why77quoq[i]) == ({wj5ongbu6[i][32-2-1:0],2'b0} & e0w_why77quoq[i][32-1:0]) ); 

      
      assign ab01vsjb5jhs3[i] = ((hlhcnhvw4wjmcl8k_oq[i] | p7icye18y8l6l[i]) & hztrxxh8s9k988m7i[i]);

      if(i == 0) begin: xvpcp9wjmb99kn
          assign v4l5fg97ku084rrubqysv[i] = ab01vsjb5jhs3[i];
      end
      else begin: efbb_rw4_pjzu4jx64w
          assign v4l5fg97ku084rrubqysv[i] = ab01vsjb5jhs3[i] & (~(|ab01vsjb5jhs3[i-1:0]));
      end

      assign de9vb1p7mqzggq3c0v4b3[i] = (oily7 ? l5dwr36cp4xs[i] : 1'b1) & (ly3dor8 ? ievzogco14[i] : 1'b1) & (p1m ? n78fb03bj00v[i] : 1'b1);

      assign cg31jos3lwbosp1uo[i] = 
                                        
                                    jmr5or9glw48yt6 ? ( (~alkw6cq4ei[i]) |  de9vb1p7mqzggq3c0v4b3[i])
                                        
                                                 : de9vb1p7mqzggq3c0v4b3[i];
 
    end
  endgenerate

  wire sgdlgdu7mr13um_lh = ~(|ab01vsjb5jhs3);

  wire ejgn5tadlr039fb = |(cg31jos3lwbosp1uo & v4l5fg97ku084rrubqysv);












































  wire qn11430de9 = (jmr5or9glw48yt6 ? sgdlgdu7mr13um_lh : 1'b0) | ejgn5tadlr039fb;

  assign foj6m18 = ~qn11430de9;

endmodule




















module y123rdlyxl0o(
  input rb050tnl,
  input a94vd35etec4,
  input el7_p8jit09,
  input [12-1:0] e1go3iu,
  input izhvh9xxvwe2,
  input  [64-1:0] vf5xcr67bqhzlo43_,
  output [64-1:0] l9erxxpnphqd26vg9,
  output u2dvoyt5e7o_03z9z5,

  output [8*32-1:0] pcr4upio7_tx37, 
  output [8*1-1:0] uzklqlncpqqm1rav,
  output [8*1-1:0] ortueunvnkx_l5m_j,
  output [8*1-1:0] hwuhtb7ucto_utk56,
  output [8*2-1:0] i1env2kmns7qvvuuc,
  output [8*1-1:0] g3s3vpafvy3i,

  input  gf33atgy,
  input  ru_wi

  );

  localparam	l_llawuowq1w9__k97nb3	= 16 ;

  wire [32-1:0] mwfdpj5fmqn8yboei  [0:l_llawuowq1w9__k97nb3-1]; 
  wire [32-1:0] wj5ongbu6  [0:l_llawuowq1w9__k97nb3-1]; 
  wire [32-1:0] htr5woms2zu1w8wv  [0:l_llawuowq1w9__k97nb3-1]; 
  wire [l_llawuowq1w9__k97nb3-1:0] vxsp5_xnwx7uki; 

  wire                  l5dwr36cp4xs [0:l_llawuowq1w9__k97nb3-1];
  wire                  ievzogco14 [0:l_llawuowq1w9__k97nb3-1];
  wire                  n78fb03bj00v [0:l_llawuowq1w9__k97nb3-1];
  wire [2-1:0]          zn3av2_qfxg [0:l_llawuowq1w9__k97nb3-1];
  wire                  alkw6cq4ei [0:l_llawuowq1w9__k97nb3-1];

  wire                  lvbsm8d9etdwan [0:l_llawuowq1w9__k97nb3-1];

  wire [64-1:0] dtr5k0nv2e4  [0:l_llawuowq1w9__k97nb3/8-1]; 

  wire [8-1:0] k8fiqgty83a   [0:l_llawuowq1w9__k97nb3-1]; 
  wire [8-1:0] ak8fp_     [0:l_llawuowq1w9__k97nb3-1]; 
  wire [8-1:0] xya8xzutptj1i3e [0:l_llawuowq1w9__k97nb3-1]; 
  wire         kplu05bi8rtxdt [0:l_llawuowq1w9__k97nb3-1];

  genvar i;

  generate 
    for (i=0; i<8; i=i+1) begin: kdmkvmzy0w
      assign pcr4upio7_tx37    [(i*32+32-1) : i*32] = wj5ongbu6 [i];
      assign uzklqlncpqqm1rav [(i*1+1-1) : i*1]                   = l5dwr36cp4xs[i];
      assign ortueunvnkx_l5m_j [(i*1+1-1) : i*1]                   = ievzogco14[i];
      assign hwuhtb7ucto_utk56 [(i*1+1-1) : i*1]                   = n78fb03bj00v[i];
      assign i1env2kmns7qvvuuc [(i*2+2-1) : i*2]                   = zn3av2_qfxg[i];
      assign g3s3vpafvy3i [(i*1+1-1) : i*1]                   = alkw6cq4ei[i];
    end
  endgenerate






















  wire[l_llawuowq1w9__k97nb3/8-1:0] f9mi9f4wgttfuvh;
  wire[l_llawuowq1w9__k97nb3/8-1:0] cqdf4hy8g8073s;
  wire[l_llawuowq1w9__k97nb3/8-1:0] x17x8iuk2nd7egtz;
  wire[l_llawuowq1w9__k97nb3/8-1:0] rgxbp_8e2wjpdachmxi4;

  wire[l_llawuowq1w9__k97nb3-1:0] wiyfv0zoxthq9d;
  wire[l_llawuowq1w9__k97nb3-1:0] nitbp_u4hkep2;
  wire[l_llawuowq1w9__k97nb3-1:0] ferpmry2dcmhe;
  wire[l_llawuowq1w9__k97nb3-1:0] gkiybei3mif_ggx;


  generate 
    for (i=0; i<l_llawuowq1w9__k97nb3/8; i=i+1) begin: m7ywpx2_8dut9x
      assign f9mi9f4wgttfuvh[i] = (e1go3iu == (12'h3A0 + {i[10:0],1'b0}));
      if (i<8/8) begin: n12eccxq1a7ypm0iiuxaa
        assign cqdf4hy8g8073s[i]  = el7_p8jit09 & f9mi9f4wgttfuvh[i];
        assign x17x8iuk2nd7egtz[i]  = a94vd35etec4 & f9mi9f4wgttfuvh[i];
        assign rgxbp_8e2wjpdachmxi4[i]  = (x17x8iuk2nd7egtz[i]  & izhvh9xxvwe2);
        assign dtr5k0nv2e4[i] = {ak8fp_[8*i+7], ak8fp_[8*i+6], ak8fp_[8*i+5], ak8fp_[8*i+4],
                                ak8fp_[8*i+3], ak8fp_[8*i+2], ak8fp_[8*i+1], ak8fp_[8*i]};
      end
      else begin: pbeg7ab23hn6qimxtpl1ntz5 
        assign cqdf4hy8g8073s[i]  = 1'b0;
        assign x17x8iuk2nd7egtz[i]  = 1'b0;
        assign rgxbp_8e2wjpdachmxi4[i]  = 1'b0;
        assign dtr5k0nv2e4[i] = {64{1'b0}};
      end
    end

    for (i=0; i<l_llawuowq1w9__k97nb3; i=i+1) begin: mm4tvvv_vb4ajq4pd1
      assign wiyfv0zoxthq9d[i] = (e1go3iu == (12'h3B0 + i[11:0]));
      if (i<8) begin: lovnmithyqtuuml45yatbn
        assign nitbp_u4hkep2[i]  = el7_p8jit09 & wiyfv0zoxthq9d[i];
        assign ferpmry2dcmhe[i]  = a94vd35etec4 & wiyfv0zoxthq9d[i];
        assign gkiybei3mif_ggx[i]  = (ferpmry2dcmhe[i] & izhvh9xxvwe2);
      end
      else begin: kvq0ra43amle4lp_xcnnbnn98y_ 
        assign nitbp_u4hkep2[i]  = 1'b0;
        assign ferpmry2dcmhe[i]  = 1'b0;
        assign gkiybei3mif_ggx[i]  = 1'b0;
      end
      if(i < (l_llawuowq1w9__k97nb3-1)) begin: bzo9jrg3dckmpbbk1lc9
        assign vxsp5_xnwx7uki[i] = gkiybei3mif_ggx[i] & (~( alkw6cq4ei[i] | lvbsm8d9etdwan[i+1] ));
      end
      if(i == (l_llawuowq1w9__k97nb3-1)) begin: q0tsqspg5zvf3j
        assign vxsp5_xnwx7uki[i] = gkiybei3mif_ggx[i] & (~( alkw6cq4ei[i] | 1'b0 ));
      end









      assign kplu05bi8rtxdt[i] = rgxbp_8e2wjpdachmxi4[i/8] & (~alkw6cq4ei[i]);



      assign lvbsm8d9etdwan[i] = 1'b0;


      assign xya8xzutptj1i3e[i][2:0] = vf5xcr67bqhzlo43_[((i%8)*8+2):((i%8)*8)];
      assign xya8xzutptj1i3e[i][4:3] = (vf5xcr67bqhzlo43_[((i%8)*8+4)] ^ vf5xcr67bqhzlo43_[((i%8)*8+3)]) ? 2'b00 : vf5xcr67bqhzlo43_[((i%8)*8+4):((i%8)*8+3)]; 
      assign xya8xzutptj1i3e[i][6:5] = 2'b0;
      assign xya8xzutptj1i3e[i][7]   = vf5xcr67bqhzlo43_[(i%8)*8+7];

      ux607_gnrl_dfflr #(8) eomoqdmimdwwtm (kplu05bi8rtxdt[i], xya8xzutptj1i3e[i], k8fiqgty83a[i], gf33atgy, ru_wi);

      assign ak8fp_[i][2:0] = k8fiqgty83a[i][2:0];

      assign ak8fp_[i][4:3] = k8fiqgty83a[i][4:3];
      assign ak8fp_[i][6:5] = 2'b0;
      assign ak8fp_[i][7]   = k8fiqgty83a[i][7]  ;

      assign l5dwr36cp4xs[i] = ak8fp_[i][0];
      assign ievzogco14[i] = ak8fp_[i][1];
      assign n78fb03bj00v[i] = ak8fp_[i][2];
      assign zn3av2_qfxg[i] = ak8fp_[i][4:3];
      assign alkw6cq4ei[i] = ak8fp_[i][7];

      assign htr5woms2zu1w8wv[i] = {2'b0,vf5xcr67bqhzlo43_[32-2-1:0]};



      assign wj5ongbu6[i][10-2:0]  = {10-1{1'b1}};
      ux607_gnrl_dfflr #(32+1-10) knk59gfmpt3wr2bb (vxsp5_xnwx7uki[i], htr5woms2zu1w8wv[i][32-1:10-1], wj5ongbu6[i][32-1:10-1], gf33atgy, ru_wi);

      assign mwfdpj5fmqn8yboei[i] = zn3av2_qfxg[i][1] ? wj5ongbu6[i] : {wj5ongbu6[i][32-1:10], {10{1'b0}}};


    end
  endgenerate








  reg [64-1:0] dd9uliud2umvee0juc7yk;
  reg u0c5hinsd9vyuxr5qv5;

  integer j;

  always @ (*) begin : j2pngj0ie
      dd9uliud2umvee0juc7yk = 64'b0;
      u0c5hinsd9vyuxr5qv5 = 1'b0;
      for(j = 0; j < l_llawuowq1w9__k97nb3/8; j = j+1) begin
        dd9uliud2umvee0juc7yk = dd9uliud2umvee0juc7yk | ({64{cqdf4hy8g8073s[j]}} & dtr5k0nv2e4[j]);
        u0c5hinsd9vyuxr5qv5 = u0c5hinsd9vyuxr5qv5 | f9mi9f4wgttfuvh[j]; 
      end

      for(j = 0; j < l_llawuowq1w9__k97nb3; j = j+1) begin


        dd9uliud2umvee0juc7yk = dd9uliud2umvee0juc7yk | ({64{nitbp_u4hkep2[j]}} & mwfdpj5fmqn8yboei[j]);
        u0c5hinsd9vyuxr5qv5 = u0c5hinsd9vyuxr5qv5 | wiyfv0zoxthq9d[j]; 
      end
  end

  assign l9erxxpnphqd26vg9 = dd9uliud2umvee0juc7yk;
  assign u2dvoyt5e7o_03z9z5 = u0c5hinsd9vyuxr5qv5;

endmodule


























































module svx57a7v0ddpyua9ju (
  input  dk2xhkj77a,    
  input  gf33atgy,        
  input  ru_wi,      
  input  gc4b3kdcan6do88ta_,  




  input  kxmsn0p4ualeps,

  input  b7ch4h6nrw1vm0,
  output rcernpf1zf4,

  input  y12wg4mlovhn13,
  output ais_l7yddpa00,

  input  b13zu8ysd3u,
  output itcmps0ezqld,



  input  j4xe_w_yjq2,
  input  aui65oshqn8b5_iz6,
  input  jmoafuo8zb_i1t,
  input  sa5of37yr6xn0s3e,
  input  j2t29hqv0s6c7,

  output o_dsdljul,
  output juyzxopct4k03sl,
  output qyqw_37_fxv8z,
  output hyw0m71z3q3rpt1,
  output fx_h7chccf02z,

  input  bf61lpqg8z,
  output dnl01g_,

  input  wz_if_2q_23jhl2,
  output n1wslu68m9v,
  output jxdeeywnwq,

  input  dyl5g2vgrvy4mb3,
  output viuu21jzrv,

  input  trtkzwpsx6l,
  output h87jx93oz7,

  input  h8xul8_er09on,
  input  emc_bywzarijbo,
  input  umnrzb6pv8dzc,
  input  nv5a7f_68p9ebw,
  input  e592323mqvany,
  input  bebngvg8sove,
  input  qz0hhqemjh,
  output ub65ja5c,
  input  vlb2az38tbnj4,
  output s_lnrw,

  output o5q5hev,
  output c8fchlpwl,
  output fid1178x5nxb,
  output erv7j3wmd3gb_dp,

  output oi60pknul, 


  output ip80u6bjne,
  output imsbh3sgxkg4,

  output klwwlfrft 
);





      
      
      
  wire yiaqce6msyt71     = kxmsn0p4ualeps | (j4xe_w_yjq2    );
  wire bgby5xqs44dvk8gqh4 = kxmsn0p4ualeps | (aui65oshqn8b5_iz6);
  wire ph3l3mocrkww4d5 = kxmsn0p4ualeps | (jmoafuo8zb_i1t);
  wire r__phg4kums7367e = kxmsn0p4ualeps | (sa5of37yr6xn0s3e);
  wire ona4gl0zwi62nzv  = kxmsn0p4ualeps | (j2t29hqv0s6c7);

  wire lhz6myl0n1vxl7 = kxmsn0p4ualeps | (h8xul8_er09on);




  wire czb4bez_5q = kxmsn0p4ualeps | (emc_bywzarijbo);
  wire hasv9p6e_t = kxmsn0p4ualeps | (umnrzb6pv8dzc);
  wire u2lp1121c2sn = kxmsn0p4ualeps | (nv5a7f_68p9ebw);
  wire lksehj4lfza2j = kxmsn0p4ualeps | (e592323mqvany);
  wire o0zbexb7mcpy10ga = kxmsn0p4ualeps | (bebngvg8sove);




  
  ux607_clkgate x4zyef7q1j752jf01(
    .clk_in   (dk2xhkj77a    ),
    .clkgate_bypass(gc4b3kdcan6do88ta_  ),
    .clock_en (y12wg4mlovhn13),
    .clk_out  (ais_l7yddpa00)
  );

  
  ux607_clkgate b40xk0vcg866n7xw(
    .clk_in   (dk2xhkj77a    ),
    .clkgate_bypass(gc4b3kdcan6do88ta_  ),
    .clock_en (b13zu8ysd3u),
    .clk_out  (itcmps0ezqld)
  );

  
  ux607_clkgate kr7d3bdmk3pmbms_(
    .clk_in   (dk2xhkj77a    ),
    .clkgate_bypass(gc4b3kdcan6do88ta_  ),
    .clock_en (b7ch4h6nrw1vm0),
    .clk_out  (rcernpf1zf4)
  );



  ux607_clkgate fwlfd3ea3mg14(
    .clk_in   (gf33atgy        ),
    .clkgate_bypass(gc4b3kdcan6do88ta_  ),
    .clock_en (yiaqce6msyt71),
    .clk_out  (o_dsdljul)
  );

  ux607_clkgate n3p_dw37_q9g7n6j0upzq(
    .clk_in   (gf33atgy        ),
    .clkgate_bypass(gc4b3kdcan6do88ta_  ),
    .clock_en (bgby5xqs44dvk8gqh4),
    .clk_out  (juyzxopct4k03sl)
  );
  ux607_clkgate l34crj101608xp2ms(
    .clk_in   (gf33atgy        ),
    .clkgate_bypass(gc4b3kdcan6do88ta_  ),
    .clock_en (ph3l3mocrkww4d5),
    .clk_out  (qyqw_37_fxv8z)
  );
  ux607_clkgate hr8y4877xfk0adn5e3eg(
    .clk_in   (gf33atgy        ),
    .clkgate_bypass(gc4b3kdcan6do88ta_  ),
    .clock_en (r__phg4kums7367e),
    .clk_out  (hyw0m71z3q3rpt1)
  );
  ux607_clkgate pz57svu1g81ykcfkp(
    .clk_in   (gf33atgy        ),
    .clkgate_bypass(gc4b3kdcan6do88ta_  ),
    .clock_en (ona4gl0zwi62nzv),
    .clk_out  (fx_h7chccf02z)
  );

  ux607_clkgate jrmzv9jq9bl5x(
    .clk_in   (gf33atgy        ),
    .clkgate_bypass(gc4b3kdcan6do88ta_  ),
    .clock_en (lhz6myl0n1vxl7),
    .clk_out  (o5q5hev)
  );

  ux607_clkgate kk_0xexqyxrrz1d(
    .clk_in   (gf33atgy        ),
    .clkgate_bypass(gc4b3kdcan6do88ta_  ),
    .clock_en (czb4bez_5q),
    .clk_out  (c8fchlpwl)
  );

  ux607_clkgate hvktokln0ezqb7c4cg(
    .clk_in   (gf33atgy        ),
    .clkgate_bypass(gc4b3kdcan6do88ta_  ),
    .clock_en (lksehj4lfza2j),
    .clk_out  (erv7j3wmd3gb_dp)
  );

  ux607_clkgate rq4gc83k_325c(
    .clk_in   (dk2xhkj77a        ),
    .clkgate_bypass(gc4b3kdcan6do88ta_  ),
    .clock_en (hasv9p6e_t),
    .clk_out  (fid1178x5nxb)
  );

  ux607_clkgate z12xs3_s_cbvvmy(
    .clk_in   (dk2xhkj77a        ),
    .clkgate_bypass(gc4b3kdcan6do88ta_  ),
    .clock_en (u2lp1121c2sn),
    .clk_out  (klwwlfrft)
  );

  ux607_clkgate ez9g00i3n88489or1f(
    .clk_in   (dk2xhkj77a        ),
    .clkgate_bypass(gc4b3kdcan6do88ta_  ),
    .clock_en (o0zbexb7mcpy10ga),
    .clk_out  (oi60pknul)
  );






  wire fls32p3vxwfiw = kxmsn0p4ualeps | wz_if_2q_23jhl2;
  assign jxdeeywnwq = ~fls32p3vxwfiw;

  ux607_clkgate mdb6ky1jikvicdpid8768(
    .clk_in   (gf33atgy        ),
    .clkgate_bypass(gc4b3kdcan6do88ta_  ),
    .clock_en (fls32p3vxwfiw),
    .clk_out  (n1wslu68m9v)
  );




  wire maa1zk26ruj16jkl_i = kxmsn0p4ualeps | dyl5g2vgrvy4mb3;
  wire dur4xgsa4i3 = ~maa1zk26ruj16jkl_i;

  ux607_clkgate okrcwiyckpri2eb84(
    .clk_in   (dk2xhkj77a        ),
    .clkgate_bypass(gc4b3kdcan6do88ta_  ),
    .clock_en (maa1zk26ruj16jkl_i),
    .clk_out  (viuu21jzrv)
  );

      
      
      
  wire aw2kqfi3l_ = kxmsn0p4ualeps | trtkzwpsx6l;

  ux607_clkgate zypp3q6_e18kf(
    .clk_in   (gf33atgy        ),
    .clkgate_bypass(gc4b3kdcan6do88ta_  ),
    .clock_en (aw2kqfi3l_),
    .clk_out  (h87jx93oz7)
  );




  wire jee2mgu95ygdk2 = kxmsn0p4ualeps | bf61lpqg8z;

  ux607_clkgate yhw8x2fnylfosm(
    .clk_in   (gf33atgy        ),
    .clkgate_bypass(gc4b3kdcan6do88ta_  ),
    .clock_en (jee2mgu95ygdk2),
    .clk_out  (dnl01g_)
  );

      
      
      
      
  wire grpf922iqr = kxmsn0p4ualeps | qz0hhqemjh;
  assign ub65ja5c = ~grpf922iqr;

  ux607_clkgate lleyqa9ezwywn(
    .clk_in   (dk2xhkj77a        ),
    .clkgate_bypass(gc4b3kdcan6do88ta_  ),
    .clock_en (grpf922iqr),
    .clk_out  (ip80u6bjne)
  );

      
      
      
      
  wire kzvoot3amvkbyop = kxmsn0p4ualeps | vlb2az38tbnj4;
  assign s_lnrw = ~kzvoot3amvkbyop;

  ux607_clkgate w7iux9eezpvls4sub(
    .clk_in   (dk2xhkj77a        ),
    .clkgate_bypass(gc4b3kdcan6do88ta_  ),
    .clock_en (kzvoot3amvkbyop),
    .clk_out  (imsbh3sgxkg4)
  );

endmodule



















module ux607_clkgate (
  input   clk_in,
  input   clkgate_bypass,
  input   clock_en,
  output  clk_out
);








reg enb;

always@(*)
  if (!clk_in)
    enb <= (clock_en | clkgate_bypass);

    assign clk_out = enb & clk_in;





endmodule 





















module ux607_reset_sync (
  input  clk,        
  input  rst_n_a,    
  input  reset_bypass,  
  output rst_n_sync 
);


localparam RST_SYNC_LEVEL = 2;

reg [RST_SYNC_LEVEL-1:0] rst_sync_r; 


always @(posedge clk or negedge rst_n_a)
begin:gen_rst_sync_PROC
  if(rst_n_a == 1'b0)
    begin
      rst_sync_r[RST_SYNC_LEVEL-1:0] <= {RST_SYNC_LEVEL{1'b0}};
    end
  else
    begin
      rst_sync_r[RST_SYNC_LEVEL-1:0] <= {rst_sync_r[RST_SYNC_LEVEL-2:0],1'b1};
    end
end

 assign rst_n_sync = reset_bypass ? rst_n_a : rst_sync_r[2-1];



endmodule




















module u9lwna1kfmt_pjd_ (

  output w41ourymsjpvm8q1e,
  input  dk2xhkj77a,    
  input  kdnujwd70g0p,
  input  k9yxnxeuf0w1,
  input  yez0ldac23i95,  








  output rb077g2alw88,


  output frilyw4z 

);


wire  i4fpck7;


wire  lx_s8lo9nrd5tedr = yez0ldac23i95 ? 1'b1 : 
                       (
                         k9yxnxeuf0w1
                       );

assign i4fpck7 = (kdnujwd70g0p & lx_s8lo9nrd5tedr);

wire pb9ckxfoinjwff;















ux607_reset_sync u_ux607_reset_sync(
  .clk      (dk2xhkj77a),
  .rst_n_a  (i4fpck7),
  .reset_bypass(yez0ldac23i95),
  .rst_n_sync(pb9ckxfoinjwff)   
);























 assign rb077g2alw88 = pb9ckxfoinjwff;


 assign frilyw4z = pb9ckxfoinjwff;

 
 
 
 
  wire c4ughu0qm5sfai;
  ux607_gnrl_dffrs #(1) dbvgqgz185u8yqz4kvb4g (1'b0, c4ughu0qm5sfai, dk2xhkj77a, rb077g2alw88);
  assign w41ourymsjpvm8q1e = c4ughu0qm5sfai;



endmodule








module u7uyomlq26a_3s81cs ( 
input  j0ln_h, 
input  p2fq1i8, 
input  pg17e0, 
output qqk5yk, 
output khfri3vm7, 
output x7bl2zxqiftsf, 
output kgg1udim46o  
);








wire   j4d0jtvzt; 
wire   ik97c06rajp2j9f3;

ux607_gnrl_dffr #(1) j9a0f3g59tmi_vntp4i_ (pg17e0, ik97c06rajp2j9f3, p2fq1i8, j0ln_h);









ux607_gnrl_dffr #(1) sp9mdoi19v9mo0_ (ik97c06rajp2j9f3, qqk5yk, p2fq1i8, j0ln_h);









ux607_gnrl_dffr #(1) hf9369s7lfrdc258m8q (qqk5yk, j4d0jtvzt, p2fq1i8, j0ln_h);









assign khfri3vm7 = qqk5yk && !j4d0jtvzt;
assign x7bl2zxqiftsf = !(qqk5yk || !j4d0jtvzt);
assign kgg1udim46o = qqk5yk ^ j4d0jtvzt;

endmodule
