 /*                                                                      
  *  Copyright (c) 2018-2020 Nuclei System Technology, Inc.              
  *  All rights reserved.                                                
  */                                                                     
                                                                         


















`include "ux607_defines.v" 

module ux607_sim_ram 
#(parameter DP = 512,
  parameter FORCE_X2ZERO = 0,
  parameter DW = 32,
  parameter MW = 4,
  parameter AW = 32 
)
(
  input             clk, 
  input  [DW-1  :0] din, 
  input  [AW-1  :0] addr,
  input             cs,
  input  [MW-1:0]   wem,
  output [DW-1:0]   dout
);

    reg [MW*8-1:0] mem_r [0:DP-1];
    reg [AW-1:0] addr_r;
    wire [MW-1:0] wen;
    wire ren;

    assign ren = cs;
    assign wen = ({MW{cs}} & wem);


    wire [MW*8-1:0] i_din; 
    generate
      if(DW == (MW*8)) begin:dw_eq_mw8
          assign i_din = din; 
      end
      else begin: dw_ne_mw8
          assign i_din = {{MW*8-DW{1'b0}},din}; 
      end
    endgenerate

    genvar i;

    always @(posedge clk)
    begin
        if (ren) begin
            addr_r <= addr;
        end
    end

    generate
      for (i = 0; i < MW; i = i+1) begin :mem
          always @(posedge clk) begin
            if (wen[i]) begin
               mem_r[addr][8*i+7:8*i] <= i_din[8*i+7:8*i];
            end
          end
      end
    endgenerate

  wire [MW*8-1:0] dout_pre;
  assign dout_pre = mem_r[addr_r];

  generate
   if(FORCE_X2ZERO == 1) begin: force_x_to_zero
      for (i = 0; i < DW; i = i+1) begin:force_x_gen 
          `ifndef SYNTHESIS
         assign dout[i] = (dout_pre[i] === 1'bx) ? 1'b0 : dout_pre[i];
          `else
         assign dout[i] = dout_pre[i];
          `endif
      end
   end
   else begin:no_force_x_to_zero
     assign dout = dout_pre[DW-1:0];
   end
  endgenerate

 
endmodule

module ux607_sim_ram_bit_en
#(parameter DP = 512,
  parameter FORCE_X2ZERO = 0,
  parameter DW = 32,
  parameter AW = 32 
)
(
  input             clk, 
  input  [DW-1  :0] din, 
  input  [AW-1  :0] addr,
  input             cs,
  input             wem,
  output [DW-1:0]   dout
);

    reg [DW-1:0] mem_r [0:DP-1];
    reg [AW-1:0] addr_r;
    wire wen;
    wire ren;

    assign ren = cs;
    assign wen = cs & wem;


    always @(posedge clk)
    begin
        if (ren) begin
            addr_r <= addr;
        end
    end

  always @(posedge clk) begin
    if (wen) begin
       mem_r[addr] <= din;
    end
  end

  wire [DW-1:0] dout_pre;
  assign dout_pre = mem_r[addr_r];

  genvar i;
  generate
   if(FORCE_X2ZERO == 1) begin: force_x_to_zero
      for (i = 0; i < DW; i = i+1) begin:force_x_gen 
          `ifndef SYNTHESIS
         assign dout[i] = (dout_pre[i] === 1'bx) ? 1'b0 : dout_pre[i];
          `else
         assign dout[i] = dout_pre[i];
          `endif
      end
   end
   else begin:no_force_x_to_zero
     assign dout = dout_pre[DW-1:0];
   end
  endgenerate

 
endmodule
